//Key = 1100000111010010100100000111101010100001110011101011001111110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354;

XOR2_X1 U748 ( .A(G107), .B(n1040), .Z(G9) );
NOR3_X1 U749 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
XNOR2_X1 U750 ( .A(KEYINPUT30), .B(n1044), .ZN(n1041) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1047), .A2(G953), .A3(G952), .ZN(n1046) );
NOR4_X1 U753 ( .A1(n1048), .A2(n1049), .A3(n1047), .A4(n1050), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
AND4_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1051) );
AND2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
AND4_X1 U757 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1047) );
NOR4_X1 U758 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
XNOR2_X1 U759 ( .A(G478), .B(n1067), .ZN(n1066) );
XOR2_X1 U760 ( .A(n1068), .B(n1069), .Z(n1063) );
NOR3_X1 U761 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1061) );
INV_X1 U762 ( .A(n1073), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
NAND2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1060) );
XOR2_X1 U765 ( .A(KEYINPUT46), .B(n1078), .Z(n1059) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1078) );
NAND3_X1 U767 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1048) );
NAND2_X1 U768 ( .A1(n1056), .A2(n1082), .ZN(n1081) );
NAND2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U770 ( .A1(n1058), .A2(n1085), .A3(n1086), .ZN(n1084) );
NAND2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NAND2_X1 U772 ( .A1(n1053), .A2(n1089), .ZN(n1088) );
XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n1090), .ZN(n1089) );
NAND2_X1 U774 ( .A1(n1055), .A2(n1091), .ZN(n1087) );
NAND2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND3_X1 U776 ( .A1(n1094), .A2(n1072), .A3(KEYINPUT8), .ZN(n1093) );
NAND2_X1 U777 ( .A1(n1055), .A2(n1095), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND3_X1 U779 ( .A1(n1094), .A2(n1072), .A3(n1098), .ZN(n1097) );
NOR3_X1 U780 ( .A1(n1065), .A2(KEYINPUT8), .A3(n1058), .ZN(n1098) );
NAND2_X1 U781 ( .A1(n1053), .A2(n1099), .ZN(n1096) );
NAND3_X1 U782 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1103), .ZN(n1102) );
NAND2_X1 U784 ( .A1(n1058), .A2(n1104), .ZN(n1100) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND3_X1 U786 ( .A1(G214), .A2(n1107), .A3(n1108), .ZN(n1106) );
NAND2_X1 U787 ( .A1(n1057), .A2(n1052), .ZN(n1105) );
INV_X1 U788 ( .A(KEYINPUT52), .ZN(n1052) );
NAND3_X1 U789 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1079) );
AND3_X1 U790 ( .A1(n1056), .A2(n1058), .A3(n1112), .ZN(n1111) );
INV_X1 U791 ( .A(n1113), .ZN(n1056) );
XNOR2_X1 U792 ( .A(n1086), .B(KEYINPUT44), .ZN(n1110) );
XNOR2_X1 U793 ( .A(n1053), .B(KEYINPUT48), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U797 ( .A1(n1120), .A2(n1080), .ZN(n1119) );
AND2_X1 U798 ( .A1(G227), .A2(G900), .ZN(n1120) );
AND3_X1 U799 ( .A1(n1118), .A2(n1121), .A3(G953), .ZN(n1116) );
NOR2_X1 U800 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1122) );
XOR2_X1 U802 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U803 ( .A1(KEYINPUT26), .A2(n1128), .ZN(n1127) );
NAND2_X1 U804 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
OR2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U806 ( .A(n1133), .B(KEYINPUT2), .Z(n1129) );
NAND2_X1 U807 ( .A1(n1132), .A2(n1131), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1134), .A2(G953), .ZN(n1114) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(G69) );
NOR2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U811 ( .A1(G224), .A2(n1080), .ZN(n1137) );
NOR3_X1 U812 ( .A1(KEYINPUT53), .A2(n1139), .A3(n1140), .ZN(n1135) );
NOR3_X1 U813 ( .A1(n1141), .A2(n1138), .A3(n1142), .ZN(n1140) );
AND3_X1 U814 ( .A1(n1141), .A2(n1080), .A3(n1142), .ZN(n1139) );
XOR2_X1 U815 ( .A(n1143), .B(KEYINPUT38), .Z(n1142) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U818 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U819 ( .A1(n1075), .A2(n1150), .ZN(n1149) );
NAND2_X1 U820 ( .A1(KEYINPUT16), .A2(n1151), .ZN(n1148) );
XOR2_X1 U821 ( .A(KEYINPUT61), .B(n1152), .Z(n1151) );
NOR2_X1 U822 ( .A1(n1146), .A2(n1153), .ZN(G63) );
XNOR2_X1 U823 ( .A(n1154), .B(n1155), .ZN(n1153) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1150), .ZN(n1155) );
NOR3_X1 U825 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(G60) );
AND3_X1 U826 ( .A1(KEYINPUT63), .A2(G953), .A3(G952), .ZN(n1159) );
NOR2_X1 U827 ( .A1(KEYINPUT63), .A2(n1160), .ZN(n1158) );
INV_X1 U828 ( .A(n1146), .ZN(n1160) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U830 ( .A(KEYINPUT51), .B(n1163), .Z(n1162) );
NOR2_X1 U831 ( .A1(n1164), .A2(n1150), .ZN(n1163) );
XNOR2_X1 U832 ( .A(G104), .B(n1165), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1146), .A2(n1166), .ZN(G57) );
XOR2_X1 U834 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U835 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U836 ( .A1(n1171), .A2(n1150), .ZN(n1170) );
NAND2_X1 U837 ( .A1(KEYINPUT41), .A2(n1172), .ZN(n1169) );
XOR2_X1 U838 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U840 ( .A(n1177), .B(KEYINPUT33), .ZN(n1173) );
NOR2_X1 U841 ( .A1(n1146), .A2(n1178), .ZN(G54) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U843 ( .A1(n1077), .A2(n1150), .ZN(n1180) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
XOR2_X1 U845 ( .A(n1183), .B(KEYINPUT40), .Z(n1182) );
NAND2_X1 U846 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U847 ( .A(KEYINPUT4), .B(n1186), .Z(n1184) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1186), .ZN(n1181) );
XNOR2_X1 U849 ( .A(n1187), .B(n1188), .ZN(n1186) );
NAND2_X1 U850 ( .A1(G227), .A2(n1080), .ZN(n1187) );
NOR2_X1 U851 ( .A1(n1146), .A2(n1189), .ZN(G51) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U853 ( .A1(n1192), .A2(n1150), .ZN(n1190) );
NAND2_X1 U854 ( .A1(G902), .A2(n1049), .ZN(n1150) );
NAND3_X1 U855 ( .A1(n1144), .A2(n1193), .A3(n1134), .ZN(n1049) );
AND4_X1 U856 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1134) );
NOR4_X1 U857 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1203), .ZN(n1196) );
NOR3_X1 U859 ( .A1(n1090), .A2(n1204), .A3(n1101), .ZN(n1203) );
NOR3_X1 U860 ( .A1(n1205), .A2(n1206), .A3(n1065), .ZN(n1202) );
NAND3_X1 U861 ( .A1(n1207), .A2(n1208), .A3(n1055), .ZN(n1205) );
NAND2_X1 U862 ( .A1(KEYINPUT62), .A2(n1204), .ZN(n1208) );
NAND2_X1 U863 ( .A1(n1209), .A2(n1210), .ZN(n1207) );
INV_X1 U864 ( .A(KEYINPUT62), .ZN(n1210) );
XOR2_X1 U865 ( .A(KEYINPUT37), .B(n1145), .Z(n1193) );
AND3_X1 U866 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1145) );
OR2_X1 U867 ( .A1(n1214), .A2(n1044), .ZN(n1213) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1216), .ZN(n1211) );
NAND2_X1 U869 ( .A1(n1090), .A2(n1043), .ZN(n1216) );
AND4_X1 U870 ( .A1(n1217), .A2(n1165), .A3(n1218), .A4(n1219), .ZN(n1144) );
NAND3_X1 U871 ( .A1(n1057), .A2(n1220), .A3(n1221), .ZN(n1218) );
XNOR2_X1 U872 ( .A(KEYINPUT13), .B(n1043), .ZN(n1220) );
NAND3_X1 U873 ( .A1(n1221), .A2(n1057), .A3(n1222), .ZN(n1165) );
INV_X1 U874 ( .A(n1042), .ZN(n1221) );
NAND3_X1 U875 ( .A1(n1223), .A2(n1224), .A3(n1058), .ZN(n1042) );
NAND3_X1 U876 ( .A1(n1223), .A2(n1103), .A3(n1225), .ZN(n1217) );
NOR2_X1 U877 ( .A1(n1080), .A2(G952), .ZN(n1146) );
XOR2_X1 U878 ( .A(G146), .B(n1200), .Z(G48) );
AND2_X1 U879 ( .A1(n1222), .A2(n1226), .ZN(n1200) );
XNOR2_X1 U880 ( .A(G143), .B(n1194), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1057), .ZN(n1194) );
XNOR2_X1 U882 ( .A(G140), .B(n1195), .ZN(G42) );
NAND4_X1 U883 ( .A1(n1222), .A2(n1086), .A3(n1229), .A4(n1103), .ZN(n1195) );
XOR2_X1 U884 ( .A(G137), .B(n1230), .Z(G39) );
NOR2_X1 U885 ( .A1(n1231), .A2(n1065), .ZN(n1230) );
XOR2_X1 U886 ( .A(n1232), .B(KEYINPUT42), .Z(n1231) );
NAND3_X1 U887 ( .A1(n1229), .A2(n1233), .A3(n1055), .ZN(n1232) );
XOR2_X1 U888 ( .A(G134), .B(n1199), .Z(G36) );
NOR3_X1 U889 ( .A1(n1204), .A2(n1043), .A3(n1101), .ZN(n1199) );
XNOR2_X1 U890 ( .A(G131), .B(n1234), .ZN(G33) );
NAND4_X1 U891 ( .A1(n1222), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1234) );
OR2_X1 U892 ( .A1(n1229), .A2(KEYINPUT3), .ZN(n1237) );
INV_X1 U893 ( .A(n1204), .ZN(n1229) );
NAND2_X1 U894 ( .A1(KEYINPUT3), .A2(n1209), .ZN(n1236) );
NAND2_X1 U895 ( .A1(n1092), .A2(n1238), .ZN(n1209) );
INV_X1 U896 ( .A(n1223), .ZN(n1092) );
INV_X1 U897 ( .A(n1101), .ZN(n1235) );
NAND2_X1 U898 ( .A1(n1228), .A2(n1086), .ZN(n1101) );
INV_X1 U899 ( .A(n1065), .ZN(n1086) );
NAND2_X1 U900 ( .A1(n1108), .A2(n1239), .ZN(n1065) );
NAND2_X1 U901 ( .A1(G214), .A2(n1107), .ZN(n1239) );
NAND2_X1 U902 ( .A1(n1240), .A2(n1241), .ZN(G30) );
NAND2_X1 U903 ( .A1(n1198), .A2(n1242), .ZN(n1241) );
XOR2_X1 U904 ( .A(KEYINPUT14), .B(n1243), .Z(n1240) );
NOR2_X1 U905 ( .A1(n1198), .A2(n1242), .ZN(n1243) );
AND2_X1 U906 ( .A1(n1226), .A2(n1112), .ZN(n1198) );
NOR3_X1 U907 ( .A1(n1206), .A2(n1044), .A3(n1204), .ZN(n1226) );
NAND2_X1 U908 ( .A1(n1223), .A2(n1238), .ZN(n1204) );
INV_X1 U909 ( .A(n1057), .ZN(n1044) );
XNOR2_X1 U910 ( .A(G101), .B(n1219), .ZN(G3) );
NAND3_X1 U911 ( .A1(n1228), .A2(n1223), .A3(n1225), .ZN(n1219) );
XOR2_X1 U912 ( .A(G125), .B(n1201), .Z(G27) );
AND3_X1 U913 ( .A1(n1053), .A2(n1222), .A3(n1244), .ZN(n1201) );
AND3_X1 U914 ( .A1(n1057), .A2(n1238), .A3(n1103), .ZN(n1244) );
NAND2_X1 U915 ( .A1(n1113), .A2(n1245), .ZN(n1238) );
NAND3_X1 U916 ( .A1(G902), .A2(n1246), .A3(n1123), .ZN(n1245) );
NOR2_X1 U917 ( .A1(n1080), .A2(G900), .ZN(n1123) );
XNOR2_X1 U918 ( .A(G122), .B(n1247), .ZN(G24) );
NAND2_X1 U919 ( .A1(n1248), .A2(n1057), .ZN(n1247) );
XOR2_X1 U920 ( .A(n1214), .B(KEYINPUT34), .Z(n1248) );
NAND4_X1 U921 ( .A1(n1227), .A2(n1053), .A3(n1058), .A4(n1224), .ZN(n1214) );
AND2_X1 U922 ( .A1(n1249), .A2(n1250), .ZN(n1227) );
XNOR2_X1 U923 ( .A(n1251), .B(KEYINPUT59), .ZN(n1249) );
XNOR2_X1 U924 ( .A(G119), .B(n1212), .ZN(G21) );
NAND3_X1 U925 ( .A1(n1053), .A2(n1233), .A3(n1225), .ZN(n1212) );
INV_X1 U926 ( .A(n1206), .ZN(n1233) );
NAND2_X1 U927 ( .A1(n1252), .A2(n1064), .ZN(n1206) );
XNOR2_X1 U928 ( .A(KEYINPUT1), .B(n1253), .ZN(n1252) );
XOR2_X1 U929 ( .A(G116), .B(n1254), .Z(G18) );
NOR3_X1 U930 ( .A1(n1255), .A2(KEYINPUT36), .A3(n1043), .ZN(n1254) );
INV_X1 U931 ( .A(n1112), .ZN(n1043) );
NOR2_X1 U932 ( .A1(n1256), .A2(n1250), .ZN(n1112) );
XOR2_X1 U933 ( .A(n1257), .B(n1258), .Z(G15) );
XNOR2_X1 U934 ( .A(G113), .B(KEYINPUT27), .ZN(n1258) );
NAND2_X1 U935 ( .A1(KEYINPUT58), .A2(n1259), .ZN(n1257) );
NAND2_X1 U936 ( .A1(n1215), .A2(n1222), .ZN(n1259) );
INV_X1 U937 ( .A(n1090), .ZN(n1222) );
NAND2_X1 U938 ( .A1(n1250), .A2(n1256), .ZN(n1090) );
INV_X1 U939 ( .A(n1255), .ZN(n1215) );
NAND4_X1 U940 ( .A1(n1053), .A2(n1228), .A3(n1057), .A4(n1224), .ZN(n1255) );
NOR2_X1 U941 ( .A1(n1253), .A2(n1260), .ZN(n1228) );
NOR2_X1 U942 ( .A1(n1261), .A2(n1072), .ZN(n1053) );
XNOR2_X1 U943 ( .A(G110), .B(n1262), .ZN(G12) );
NAND3_X1 U944 ( .A1(n1225), .A2(n1103), .A3(n1263), .ZN(n1262) );
XNOR2_X1 U945 ( .A(n1223), .B(KEYINPUT0), .ZN(n1263) );
NOR2_X1 U946 ( .A1(n1094), .A2(n1072), .ZN(n1223) );
AND2_X1 U947 ( .A1(G221), .A2(n1264), .ZN(n1072) );
INV_X1 U948 ( .A(n1261), .ZN(n1094) );
XOR2_X1 U949 ( .A(n1076), .B(n1265), .Z(n1261) );
NOR2_X1 U950 ( .A1(KEYINPUT47), .A2(n1077), .ZN(n1265) );
INV_X1 U951 ( .A(G469), .ZN(n1077) );
AND2_X1 U952 ( .A1(n1266), .A2(n1267), .ZN(n1076) );
XNOR2_X1 U953 ( .A(n1188), .B(n1268), .ZN(n1266) );
XNOR2_X1 U954 ( .A(n1269), .B(n1270), .ZN(n1268) );
NOR2_X1 U955 ( .A1(KEYINPUT49), .A2(n1185), .ZN(n1270) );
XNOR2_X1 U956 ( .A(n1271), .B(n1272), .ZN(n1185) );
XNOR2_X1 U957 ( .A(n1273), .B(n1274), .ZN(n1272) );
XNOR2_X1 U958 ( .A(KEYINPUT28), .B(n1275), .ZN(n1274) );
INV_X1 U959 ( .A(G104), .ZN(n1275) );
XOR2_X1 U960 ( .A(n1276), .B(n1128), .Z(n1271) );
XNOR2_X1 U961 ( .A(n1277), .B(n1278), .ZN(n1128) );
NAND2_X1 U962 ( .A1(KEYINPUT55), .A2(n1279), .ZN(n1277) );
XNOR2_X1 U963 ( .A(G146), .B(n1280), .ZN(n1279) );
XOR2_X1 U964 ( .A(n1175), .B(n1281), .Z(n1276) );
NOR2_X1 U965 ( .A1(G107), .A2(KEYINPUT18), .ZN(n1281) );
NOR2_X1 U966 ( .A1(KEYINPUT21), .A2(n1121), .ZN(n1269) );
INV_X1 U967 ( .A(G227), .ZN(n1121) );
XNOR2_X1 U968 ( .A(G110), .B(n1282), .ZN(n1188) );
NAND2_X1 U969 ( .A1(n1283), .A2(n1284), .ZN(n1103) );
NAND2_X1 U970 ( .A1(n1058), .A2(n1285), .ZN(n1284) );
INV_X1 U971 ( .A(KEYINPUT1), .ZN(n1285) );
NOR2_X1 U972 ( .A1(n1253), .A2(n1064), .ZN(n1058) );
NAND3_X1 U973 ( .A1(n1260), .A2(n1253), .A3(KEYINPUT1), .ZN(n1283) );
NAND3_X1 U974 ( .A1(n1286), .A2(n1287), .A3(n1073), .ZN(n1253) );
NAND2_X1 U975 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U976 ( .A1(KEYINPUT24), .A2(n1075), .ZN(n1287) );
OR3_X1 U977 ( .A1(n1074), .A2(KEYINPUT24), .A3(n1075), .ZN(n1286) );
NAND2_X1 U978 ( .A1(G217), .A2(n1264), .ZN(n1075) );
NAND2_X1 U979 ( .A1(n1288), .A2(n1267), .ZN(n1264) );
AND2_X1 U980 ( .A1(n1152), .A2(n1267), .ZN(n1074) );
XNOR2_X1 U981 ( .A(n1289), .B(n1290), .ZN(n1152) );
XOR2_X1 U982 ( .A(G137), .B(n1291), .Z(n1290) );
NOR2_X1 U983 ( .A1(KEYINPUT23), .A2(n1292), .ZN(n1291) );
XOR2_X1 U984 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U985 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U986 ( .A(G125), .B(G119), .Z(n1296) );
XOR2_X1 U987 ( .A(KEYINPUT7), .B(G146), .Z(n1295) );
XOR2_X1 U988 ( .A(n1297), .B(n1278), .Z(n1293) );
XNOR2_X1 U989 ( .A(n1298), .B(n1299), .ZN(n1297) );
NAND2_X1 U990 ( .A1(KEYINPUT19), .A2(n1282), .ZN(n1298) );
NAND2_X1 U991 ( .A1(G221), .A2(n1300), .ZN(n1289) );
INV_X1 U992 ( .A(n1064), .ZN(n1260) );
XOR2_X1 U993 ( .A(n1301), .B(n1171), .Z(n1064) );
INV_X1 U994 ( .A(G472), .ZN(n1171) );
NAND2_X1 U995 ( .A1(n1302), .A2(n1267), .ZN(n1301) );
XOR2_X1 U996 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U997 ( .A(n1176), .B(n1167), .ZN(n1304) );
XNOR2_X1 U998 ( .A(n1305), .B(n1273), .ZN(n1167) );
INV_X1 U999 ( .A(G101), .ZN(n1273) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U1001 ( .A(n1307), .B(n1308), .ZN(n1176) );
XOR2_X1 U1002 ( .A(KEYINPUT29), .B(G119), .Z(n1308) );
XOR2_X1 U1003 ( .A(n1309), .B(G113), .Z(n1307) );
NAND2_X1 U1004 ( .A1(KEYINPUT57), .A2(G116), .ZN(n1309) );
XNOR2_X1 U1005 ( .A(n1177), .B(n1310), .ZN(n1303) );
XNOR2_X1 U1006 ( .A(n1311), .B(KEYINPUT25), .ZN(n1310) );
NAND2_X1 U1007 ( .A1(KEYINPUT56), .A2(n1175), .ZN(n1311) );
XNOR2_X1 U1008 ( .A(n1131), .B(n1312), .ZN(n1175) );
XNOR2_X1 U1009 ( .A(KEYINPUT17), .B(n1132), .ZN(n1312) );
XNOR2_X1 U1010 ( .A(G131), .B(KEYINPUT32), .ZN(n1132) );
XOR2_X1 U1011 ( .A(G134), .B(G137), .Z(n1131) );
AND3_X1 U1012 ( .A1(n1057), .A2(n1224), .A3(n1055), .ZN(n1225) );
NOR2_X1 U1013 ( .A1(n1250), .A2(n1251), .ZN(n1055) );
INV_X1 U1014 ( .A(n1256), .ZN(n1251) );
NAND2_X1 U1015 ( .A1(n1313), .A2(n1314), .ZN(n1256) );
NAND2_X1 U1016 ( .A1(n1315), .A2(n1156), .ZN(n1314) );
INV_X1 U1017 ( .A(G478), .ZN(n1156) );
XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(n1067), .ZN(n1315) );
NAND2_X1 U1019 ( .A1(n1316), .A2(G478), .ZN(n1313) );
XOR2_X1 U1020 ( .A(n1067), .B(KEYINPUT9), .Z(n1316) );
NAND2_X1 U1021 ( .A1(n1317), .A2(n1267), .ZN(n1067) );
XNOR2_X1 U1022 ( .A(KEYINPUT12), .B(n1318), .ZN(n1317) );
INV_X1 U1023 ( .A(n1154), .ZN(n1318) );
XNOR2_X1 U1024 ( .A(n1319), .B(n1320), .ZN(n1154) );
XOR2_X1 U1025 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1026 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1027 ( .A1(KEYINPUT43), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1028 ( .A(KEYINPUT5), .B(G134), .Z(n1325) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1300), .ZN(n1323) );
AND2_X1 U1030 ( .A1(G234), .A2(n1080), .ZN(n1300) );
XOR2_X1 U1031 ( .A(n1326), .B(n1327), .Z(n1319) );
NOR2_X1 U1032 ( .A1(KEYINPUT60), .A2(G107), .ZN(n1327) );
XNOR2_X1 U1033 ( .A(G122), .B(G116), .ZN(n1326) );
XNOR2_X1 U1034 ( .A(n1328), .B(n1069), .ZN(n1250) );
XNOR2_X1 U1035 ( .A(n1164), .B(KEYINPUT11), .ZN(n1069) );
INV_X1 U1036 ( .A(G475), .ZN(n1164) );
NAND2_X1 U1037 ( .A1(KEYINPUT54), .A2(n1068), .ZN(n1328) );
NAND2_X1 U1038 ( .A1(n1161), .A2(n1267), .ZN(n1068) );
XNOR2_X1 U1039 ( .A(n1329), .B(n1330), .ZN(n1161) );
XOR2_X1 U1040 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1041 ( .A(n1333), .B(n1124), .Z(n1332) );
XNOR2_X1 U1042 ( .A(G125), .B(n1282), .ZN(n1124) );
INV_X1 U1043 ( .A(G140), .ZN(n1282) );
XOR2_X1 U1044 ( .A(n1334), .B(n1335), .Z(n1331) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1306), .ZN(n1335) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1306) );
NAND2_X1 U1047 ( .A1(KEYINPUT39), .A2(G146), .ZN(n1334) );
XOR2_X1 U1048 ( .A(n1336), .B(n1337), .Z(n1329) );
XOR2_X1 U1049 ( .A(KEYINPUT20), .B(G131), .Z(n1337) );
XNOR2_X1 U1050 ( .A(G104), .B(n1338), .ZN(n1336) );
NOR2_X1 U1051 ( .A1(KEYINPUT31), .A2(n1280), .ZN(n1338) );
INV_X1 U1052 ( .A(G143), .ZN(n1280) );
NAND2_X1 U1053 ( .A1(n1113), .A2(n1339), .ZN(n1224) );
NAND3_X1 U1054 ( .A1(n1138), .A2(n1246), .A3(G902), .ZN(n1339) );
NOR2_X1 U1055 ( .A1(G898), .A2(n1080), .ZN(n1138) );
NAND3_X1 U1056 ( .A1(n1246), .A2(n1080), .A3(G952), .ZN(n1113) );
NAND2_X1 U1057 ( .A1(G237), .A2(n1288), .ZN(n1246) );
XOR2_X1 U1058 ( .A(G234), .B(KEYINPUT10), .Z(n1288) );
NOR2_X1 U1059 ( .A1(n1108), .A2(n1340), .ZN(n1057) );
AND2_X1 U1060 ( .A1(G214), .A2(n1107), .ZN(n1340) );
XNOR2_X1 U1061 ( .A(n1341), .B(n1192), .ZN(n1108) );
NAND2_X1 U1062 ( .A1(G210), .A2(n1107), .ZN(n1192) );
NAND2_X1 U1063 ( .A1(n1342), .A2(n1343), .ZN(n1107) );
INV_X1 U1064 ( .A(G237), .ZN(n1343) );
XNOR2_X1 U1065 ( .A(KEYINPUT45), .B(n1267), .ZN(n1342) );
INV_X1 U1066 ( .A(G902), .ZN(n1267) );
OR2_X1 U1067 ( .A1(n1191), .A2(G902), .ZN(n1341) );
XNOR2_X1 U1068 ( .A(n1344), .B(n1345), .ZN(n1191) );
XOR2_X1 U1069 ( .A(G125), .B(n1346), .Z(n1345) );
AND2_X1 U1070 ( .A1(n1080), .A2(G224), .ZN(n1346) );
INV_X1 U1071 ( .A(G953), .ZN(n1080) );
XNOR2_X1 U1072 ( .A(n1143), .B(n1347), .ZN(n1344) );
INV_X1 U1073 ( .A(n1177), .ZN(n1347) );
XNOR2_X1 U1074 ( .A(n1321), .B(G146), .ZN(n1177) );
XNOR2_X1 U1075 ( .A(G143), .B(n1278), .ZN(n1321) );
XNOR2_X1 U1076 ( .A(n1242), .B(KEYINPUT6), .ZN(n1278) );
INV_X1 U1077 ( .A(G128), .ZN(n1242) );
XOR2_X1 U1078 ( .A(n1348), .B(n1349), .Z(n1143) );
XNOR2_X1 U1079 ( .A(n1333), .B(n1350), .ZN(n1349) );
XNOR2_X1 U1080 ( .A(n1351), .B(n1352), .ZN(n1350) );
NOR2_X1 U1081 ( .A1(G119), .A2(KEYINPUT35), .ZN(n1352) );
NOR2_X1 U1082 ( .A1(KEYINPUT15), .A2(n1353), .ZN(n1351) );
XNOR2_X1 U1083 ( .A(G104), .B(G107), .ZN(n1353) );
XOR2_X1 U1084 ( .A(G113), .B(G122), .Z(n1333) );
XNOR2_X1 U1085 ( .A(G101), .B(n1354), .ZN(n1348) );
XNOR2_X1 U1086 ( .A(G116), .B(n1299), .ZN(n1354) );
INV_X1 U1087 ( .A(G110), .ZN(n1299) );
endmodule


