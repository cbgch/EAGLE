//Key = 0001001101111010011111101000001101001001001000011001101010000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XOR2_X1 U721 ( .A(n1009), .B(n1010), .Z(G9) );
NAND2_X1 U722 ( .A1(KEYINPUT56), .A2(G107), .ZN(n1010) );
NAND3_X1 U723 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(G75) );
NAND2_X1 U724 ( .A1(G952), .A2(n1014), .ZN(n1013) );
NAND3_X1 U725 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND2_X1 U726 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NAND2_X1 U727 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND3_X1 U728 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NAND2_X1 U729 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND2_X1 U730 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
OR2_X1 U731 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U732 ( .A1(n1031), .A2(n1032), .ZN(n1025) );
NAND2_X1 U733 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U734 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND3_X1 U735 ( .A1(n1031), .A2(n1037), .A3(n1027), .ZN(n1020) );
NAND2_X1 U736 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U737 ( .A1(n1024), .A2(n1040), .ZN(n1039) );
OR2_X1 U738 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U739 ( .A1(n1022), .A2(n1043), .ZN(n1038) );
NAND2_X1 U740 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U741 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XNOR2_X1 U742 ( .A(n1048), .B(KEYINPUT58), .ZN(n1046) );
INV_X1 U743 ( .A(n1049), .ZN(n1018) );
NAND2_X1 U744 ( .A1(KEYINPUT0), .A2(n1050), .ZN(n1015) );
NAND2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(n1011) );
NAND2_X1 U746 ( .A1(KEYINPUT0), .A2(G952), .ZN(n1052) );
INV_X1 U747 ( .A(n1050), .ZN(n1051) );
NAND4_X1 U748 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1050) );
NOR4_X1 U749 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
XNOR2_X1 U750 ( .A(KEYINPUT60), .B(n1061), .ZN(n1060) );
XOR2_X1 U751 ( .A(KEYINPUT27), .B(n1062), .Z(n1059) );
NOR2_X1 U752 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U753 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XNOR2_X1 U754 ( .A(KEYINPUT55), .B(n1067), .ZN(n1066) );
XNOR2_X1 U755 ( .A(n1068), .B(n1069), .ZN(n1058) );
NAND2_X1 U756 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NAND2_X1 U757 ( .A1(KEYINPUT2), .A2(n1072), .ZN(n1071) );
NAND2_X1 U758 ( .A1(KEYINPUT18), .A2(n1073), .ZN(n1070) );
NOR3_X1 U759 ( .A1(n1074), .A2(n1035), .A3(n1075), .ZN(n1055) );
INV_X1 U760 ( .A(n1076), .ZN(n1075) );
XNOR2_X1 U761 ( .A(n1077), .B(n1078), .ZN(n1074) );
NAND2_X1 U762 ( .A1(KEYINPUT63), .A2(n1079), .ZN(n1077) );
XOR2_X1 U763 ( .A(G475), .B(n1080), .Z(n1054) );
NOR2_X1 U764 ( .A1(KEYINPUT35), .A2(n1081), .ZN(n1080) );
XNOR2_X1 U765 ( .A(KEYINPUT49), .B(n1082), .ZN(n1081) );
XOR2_X1 U766 ( .A(KEYINPUT36), .B(n1047), .Z(n1053) );
NAND2_X1 U767 ( .A1(n1083), .A2(n1084), .ZN(G72) );
NAND2_X1 U768 ( .A1(n1085), .A2(n1012), .ZN(n1084) );
XNOR2_X1 U769 ( .A(n1086), .B(n1087), .ZN(n1085) );
NOR2_X1 U770 ( .A1(n1088), .A2(KEYINPUT53), .ZN(n1087) );
INV_X1 U771 ( .A(n1089), .ZN(n1088) );
NAND2_X1 U772 ( .A1(n1090), .A2(G953), .ZN(n1083) );
XOR2_X1 U773 ( .A(n1086), .B(n1091), .Z(n1090) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1091) );
NAND2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1086) );
NAND2_X1 U776 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U777 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U778 ( .A(KEYINPUT40), .B(n1097), .Z(n1096) );
XOR2_X1 U779 ( .A(KEYINPUT8), .B(KEYINPUT57), .Z(n1097) );
XNOR2_X1 U780 ( .A(n1098), .B(n1099), .ZN(n1095) );
XOR2_X1 U781 ( .A(n1100), .B(n1101), .Z(n1098) );
XOR2_X1 U782 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND3_X1 U784 ( .A1(n1106), .A2(n1107), .A3(KEYINPUT48), .ZN(n1105) );
NAND2_X1 U785 ( .A1(n1108), .A2(G953), .ZN(n1107) );
XNOR2_X1 U786 ( .A(G898), .B(KEYINPUT44), .ZN(n1108) );
NAND2_X1 U787 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
XNOR2_X1 U788 ( .A(KEYINPUT10), .B(n1012), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1111), .A2(n1012), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XOR2_X1 U792 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U793 ( .A1(n1118), .A2(G217), .ZN(n1116) );
NOR2_X1 U794 ( .A1(n1119), .A2(n1120), .ZN(G63) );
XOR2_X1 U795 ( .A(KEYINPUT13), .B(n1114), .Z(n1120) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1119) );
NAND2_X1 U797 ( .A1(n1118), .A2(G478), .ZN(n1121) );
NOR3_X1 U798 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(G60) );
AND2_X1 U799 ( .A1(KEYINPUT6), .A2(n1114), .ZN(n1125) );
NOR3_X1 U800 ( .A1(KEYINPUT6), .A2(G953), .A3(G952), .ZN(n1124) );
XOR2_X1 U801 ( .A(n1126), .B(n1127), .Z(n1123) );
NAND2_X1 U802 ( .A1(n1118), .A2(G475), .ZN(n1126) );
XOR2_X1 U803 ( .A(G104), .B(n1128), .Z(G6) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1129), .ZN(G57) );
XNOR2_X1 U805 ( .A(n1130), .B(n1131), .ZN(n1129) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U807 ( .A1(KEYINPUT1), .A2(n1134), .ZN(n1133) );
XOR2_X1 U808 ( .A(KEYINPUT54), .B(n1135), .Z(n1134) );
NAND2_X1 U809 ( .A1(n1118), .A2(G472), .ZN(n1132) );
NOR2_X1 U810 ( .A1(n1114), .A2(n1136), .ZN(G54) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR3_X1 U813 ( .A1(n1079), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR2_X1 U814 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
INV_X1 U815 ( .A(KEYINPUT4), .ZN(n1144) );
NOR2_X1 U816 ( .A1(n1017), .A2(G902), .ZN(n1143) );
NOR2_X1 U817 ( .A1(KEYINPUT4), .A2(n1118), .ZN(n1141) );
INV_X1 U818 ( .A(G469), .ZN(n1079) );
NOR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
XOR2_X1 U820 ( .A(KEYINPUT5), .B(n1147), .Z(n1146) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
AND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
XNOR2_X1 U823 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1114), .A2(n1152), .ZN(G51) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U826 ( .A(KEYINPUT28), .B(n1155), .Z(n1154) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
AND2_X1 U828 ( .A1(n1157), .A2(n1156), .ZN(n1153) );
XOR2_X1 U829 ( .A(n1106), .B(n1158), .Z(n1156) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
INV_X1 U831 ( .A(n1161), .ZN(n1160) );
NAND2_X1 U832 ( .A1(n1118), .A2(n1073), .ZN(n1157) );
INV_X1 U833 ( .A(n1072), .ZN(n1073) );
NOR2_X1 U834 ( .A1(n1162), .A2(n1017), .ZN(n1118) );
NOR2_X1 U835 ( .A1(n1110), .A2(n1089), .ZN(n1017) );
NAND4_X1 U836 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1089) );
NOR4_X1 U837 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
NOR2_X1 U839 ( .A1(n1033), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U840 ( .A(KEYINPUT42), .B(n1174), .ZN(n1173) );
INV_X1 U841 ( .A(n1175), .ZN(n1171) );
NAND4_X1 U842 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1110) );
AND4_X1 U843 ( .A1(n1009), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1179) );
NAND3_X1 U844 ( .A1(n1031), .A2(n1042), .A3(n1183), .ZN(n1009) );
NOR2_X1 U845 ( .A1(n1128), .A2(n1184), .ZN(n1178) );
NOR2_X1 U846 ( .A1(n1033), .A2(n1185), .ZN(n1184) );
AND3_X1 U847 ( .A1(n1183), .A2(n1031), .A3(n1041), .ZN(n1128) );
NAND3_X1 U848 ( .A1(n1029), .A2(n1183), .A3(n1186), .ZN(n1176) );
XNOR2_X1 U849 ( .A(KEYINPUT21), .B(n1022), .ZN(n1186) );
NOR2_X1 U850 ( .A1(n1012), .A2(G952), .ZN(n1114) );
XOR2_X1 U851 ( .A(G146), .B(n1187), .Z(G48) );
NOR3_X1 U852 ( .A1(n1174), .A2(KEYINPUT34), .A3(n1033), .ZN(n1187) );
NAND2_X1 U853 ( .A1(n1188), .A2(n1041), .ZN(n1174) );
NAND2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(G45) );
NAND2_X1 U855 ( .A1(G143), .A2(n1175), .ZN(n1190) );
XOR2_X1 U856 ( .A(n1191), .B(KEYINPUT16), .Z(n1189) );
OR2_X1 U857 ( .A1(n1175), .A2(G143), .ZN(n1191) );
NAND2_X1 U858 ( .A1(n1192), .A2(n1193), .ZN(n1175) );
XOR2_X1 U859 ( .A(G140), .B(n1169), .Z(G42) );
AND4_X1 U860 ( .A1(n1027), .A2(n1029), .A3(n1194), .A4(n1041), .ZN(n1169) );
NOR2_X1 U861 ( .A1(n1195), .A2(n1044), .ZN(n1194) );
XNOR2_X1 U862 ( .A(G137), .B(n1196), .ZN(G39) );
NOR2_X1 U863 ( .A1(n1168), .A2(KEYINPUT46), .ZN(n1196) );
AND3_X1 U864 ( .A1(n1188), .A2(n1022), .A3(n1027), .ZN(n1168) );
XNOR2_X1 U865 ( .A(G134), .B(n1163), .ZN(G36) );
NAND3_X1 U866 ( .A1(n1027), .A2(n1042), .A3(n1192), .ZN(n1163) );
XOR2_X1 U867 ( .A(n1164), .B(n1197), .Z(G33) );
NOR2_X1 U868 ( .A1(G131), .A2(KEYINPUT25), .ZN(n1197) );
NAND3_X1 U869 ( .A1(n1027), .A2(n1041), .A3(n1192), .ZN(n1164) );
NOR3_X1 U870 ( .A1(n1044), .A2(n1195), .A3(n1198), .ZN(n1192) );
INV_X1 U871 ( .A(n1199), .ZN(n1195) );
AND2_X1 U872 ( .A1(n1200), .A2(n1036), .ZN(n1027) );
XOR2_X1 U873 ( .A(KEYINPUT20), .B(n1035), .Z(n1200) );
XOR2_X1 U874 ( .A(G128), .B(n1167), .Z(G30) );
AND3_X1 U875 ( .A1(n1201), .A2(n1042), .A3(n1188), .ZN(n1167) );
AND4_X1 U876 ( .A1(n1202), .A2(n1057), .A3(n1199), .A4(n1203), .ZN(n1188) );
XNOR2_X1 U877 ( .A(G101), .B(n1177), .ZN(G3) );
NAND3_X1 U878 ( .A1(n1183), .A2(n1022), .A3(n1030), .ZN(n1177) );
XOR2_X1 U879 ( .A(G125), .B(n1170), .Z(G27) );
AND4_X1 U880 ( .A1(n1201), .A2(n1029), .A3(n1204), .A4(n1041), .ZN(n1170) );
AND2_X1 U881 ( .A1(n1199), .A2(n1024), .ZN(n1204) );
NAND2_X1 U882 ( .A1(n1049), .A2(n1205), .ZN(n1199) );
NAND4_X1 U883 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1094), .ZN(n1205) );
INV_X1 U884 ( .A(G900), .ZN(n1094) );
XNOR2_X1 U885 ( .A(G122), .B(n1182), .ZN(G24) );
NAND3_X1 U886 ( .A1(n1207), .A2(n1031), .A3(n1193), .ZN(n1182) );
AND3_X1 U887 ( .A1(n1208), .A2(n1209), .A3(n1201), .ZN(n1193) );
NOR2_X1 U888 ( .A1(n1203), .A2(n1057), .ZN(n1031) );
XNOR2_X1 U889 ( .A(G119), .B(n1210), .ZN(G21) );
NAND2_X1 U890 ( .A1(n1211), .A2(n1201), .ZN(n1210) );
XOR2_X1 U891 ( .A(n1185), .B(KEYINPUT11), .Z(n1211) );
NAND4_X1 U892 ( .A1(n1207), .A2(n1022), .A3(n1057), .A4(n1203), .ZN(n1185) );
NAND2_X1 U893 ( .A1(n1212), .A2(n1213), .ZN(G18) );
OR2_X1 U894 ( .A1(n1181), .A2(G116), .ZN(n1213) );
XOR2_X1 U895 ( .A(n1214), .B(KEYINPUT26), .Z(n1212) );
NAND2_X1 U896 ( .A1(G116), .A2(n1181), .ZN(n1214) );
NAND4_X1 U897 ( .A1(n1201), .A2(n1030), .A3(n1207), .A4(n1042), .ZN(n1181) );
AND2_X1 U898 ( .A1(n1208), .A2(n1215), .ZN(n1042) );
XNOR2_X1 U899 ( .A(n1216), .B(n1209), .ZN(n1215) );
INV_X1 U900 ( .A(n1033), .ZN(n1201) );
XOR2_X1 U901 ( .A(n1217), .B(KEYINPUT61), .Z(n1033) );
XNOR2_X1 U902 ( .A(G113), .B(n1180), .ZN(G15) );
NAND4_X1 U903 ( .A1(n1030), .A2(n1207), .A3(n1041), .A4(n1217), .ZN(n1180) );
AND2_X1 U904 ( .A1(n1024), .A2(n1218), .ZN(n1207) );
NOR2_X1 U905 ( .A1(n1048), .A2(n1047), .ZN(n1024) );
INV_X1 U906 ( .A(n1198), .ZN(n1030) );
NAND2_X1 U907 ( .A1(n1219), .A2(n1057), .ZN(n1198) );
XNOR2_X1 U908 ( .A(G110), .B(n1220), .ZN(G12) );
NAND3_X1 U909 ( .A1(n1221), .A2(n1022), .A3(n1183), .ZN(n1220) );
AND3_X1 U910 ( .A1(n1217), .A2(n1218), .A3(n1202), .ZN(n1183) );
INV_X1 U911 ( .A(n1044), .ZN(n1202) );
NAND2_X1 U912 ( .A1(n1222), .A2(n1048), .ZN(n1044) );
XNOR2_X1 U913 ( .A(n1078), .B(G469), .ZN(n1048) );
NAND2_X1 U914 ( .A1(n1223), .A2(n1224), .ZN(n1078) );
XOR2_X1 U915 ( .A(n1137), .B(n1225), .Z(n1223) );
NOR2_X1 U916 ( .A1(KEYINPUT43), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U917 ( .A(n1227), .B(n1148), .ZN(n1226) );
NAND2_X1 U918 ( .A1(n1228), .A2(KEYINPUT24), .ZN(n1227) );
XOR2_X1 U919 ( .A(n1229), .B(n1151), .Z(n1228) );
XNOR2_X1 U920 ( .A(n1099), .B(KEYINPUT14), .ZN(n1151) );
NAND2_X1 U921 ( .A1(KEYINPUT19), .A2(n1150), .ZN(n1229) );
NAND3_X1 U922 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1150) );
NAND3_X1 U923 ( .A1(KEYINPUT33), .A2(n1233), .A3(n1234), .ZN(n1231) );
OR2_X1 U924 ( .A1(n1234), .A2(KEYINPUT33), .ZN(n1230) );
XOR2_X1 U925 ( .A(n1235), .B(n1236), .Z(n1137) );
XNOR2_X1 U926 ( .A(G140), .B(n1237), .ZN(n1236) );
NAND2_X1 U927 ( .A1(G227), .A2(n1012), .ZN(n1235) );
XOR2_X1 U928 ( .A(KEYINPUT9), .B(n1047), .Z(n1222) );
AND2_X1 U929 ( .A1(G221), .A2(n1238), .ZN(n1047) );
NAND2_X1 U930 ( .A1(n1049), .A2(n1239), .ZN(n1218) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1113), .ZN(n1239) );
INV_X1 U932 ( .A(G898), .ZN(n1113) );
NAND3_X1 U933 ( .A1(n1206), .A2(n1012), .A3(G952), .ZN(n1049) );
NAND2_X1 U934 ( .A1(G237), .A2(G234), .ZN(n1206) );
NOR2_X1 U935 ( .A1(n1036), .A2(n1035), .ZN(n1217) );
AND2_X1 U936 ( .A1(G214), .A2(n1240), .ZN(n1035) );
XOR2_X1 U937 ( .A(n1241), .B(n1072), .Z(n1036) );
NAND2_X1 U938 ( .A1(G210), .A2(n1240), .ZN(n1072) );
NAND2_X1 U939 ( .A1(n1162), .A2(n1242), .ZN(n1240) );
INV_X1 U940 ( .A(G237), .ZN(n1242) );
NAND2_X1 U941 ( .A1(KEYINPUT39), .A2(n1069), .ZN(n1241) );
NAND2_X1 U942 ( .A1(n1224), .A2(n1243), .ZN(n1069) );
XNOR2_X1 U943 ( .A(n1106), .B(n1244), .ZN(n1243) );
NAND3_X1 U944 ( .A1(n1245), .A2(n1246), .A3(n1161), .ZN(n1244) );
NAND2_X1 U945 ( .A1(n1247), .A2(n1248), .ZN(n1161) );
NAND2_X1 U946 ( .A1(G224), .A2(n1012), .ZN(n1248) );
NAND2_X1 U947 ( .A1(n1159), .A2(n1249), .ZN(n1246) );
INV_X1 U948 ( .A(KEYINPUT50), .ZN(n1249) );
NOR3_X1 U949 ( .A1(n1112), .A2(G953), .A3(n1247), .ZN(n1159) );
INV_X1 U950 ( .A(G224), .ZN(n1112) );
NAND2_X1 U951 ( .A1(KEYINPUT50), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U952 ( .A(G125), .B(n1099), .ZN(n1247) );
AND2_X1 U953 ( .A1(n1250), .A2(n1251), .ZN(n1106) );
NAND3_X1 U954 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
XOR2_X1 U955 ( .A(n1255), .B(n1256), .Z(n1252) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1258), .ZN(n1250) );
NAND2_X1 U957 ( .A1(n1254), .A2(n1253), .ZN(n1258) );
NAND2_X1 U958 ( .A1(n1259), .A2(n1260), .ZN(n1253) );
XNOR2_X1 U959 ( .A(KEYINPUT38), .B(n1237), .ZN(n1259) );
XOR2_X1 U960 ( .A(n1261), .B(KEYINPUT32), .Z(n1254) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U962 ( .A(KEYINPUT38), .B(G110), .ZN(n1263) );
XNOR2_X1 U963 ( .A(G122), .B(KEYINPUT22), .ZN(n1262) );
XNOR2_X1 U964 ( .A(n1255), .B(n1256), .ZN(n1257) );
XNOR2_X1 U965 ( .A(n1264), .B(n1265), .ZN(n1256) );
NOR2_X1 U966 ( .A1(KEYINPUT37), .A2(n1266), .ZN(n1265) );
INV_X1 U967 ( .A(n1267), .ZN(n1266) );
NAND2_X1 U968 ( .A1(n1268), .A2(n1232), .ZN(n1255) );
OR2_X1 U969 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U970 ( .A1(n1269), .A2(n1233), .ZN(n1268) );
INV_X1 U971 ( .A(G107), .ZN(n1233) );
XNOR2_X1 U972 ( .A(KEYINPUT12), .B(n1234), .ZN(n1269) );
XOR2_X1 U973 ( .A(G104), .B(n1270), .Z(n1234) );
NAND2_X1 U974 ( .A1(n1271), .A2(n1272), .ZN(n1022) );
NAND2_X1 U975 ( .A1(n1041), .A2(n1216), .ZN(n1272) );
NOR2_X1 U976 ( .A1(n1208), .A2(n1273), .ZN(n1041) );
INV_X1 U977 ( .A(n1209), .ZN(n1273) );
OR3_X1 U978 ( .A1(n1208), .A2(n1209), .A3(n1216), .ZN(n1271) );
INV_X1 U979 ( .A(KEYINPUT51), .ZN(n1216) );
XNOR2_X1 U980 ( .A(n1082), .B(G475), .ZN(n1209) );
NAND2_X1 U981 ( .A1(n1224), .A2(n1127), .ZN(n1082) );
XNOR2_X1 U982 ( .A(n1274), .B(n1275), .ZN(n1127) );
XOR2_X1 U983 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U984 ( .A(n1278), .B(G104), .ZN(n1277) );
INV_X1 U985 ( .A(G113), .ZN(n1278) );
XNOR2_X1 U986 ( .A(G131), .B(n1260), .ZN(n1276) );
XOR2_X1 U987 ( .A(n1279), .B(n1280), .Z(n1274) );
XOR2_X1 U988 ( .A(n1281), .B(n1101), .Z(n1279) );
NAND2_X1 U989 ( .A1(n1282), .A2(G214), .ZN(n1281) );
NAND2_X1 U990 ( .A1(n1283), .A2(n1284), .ZN(n1208) );
NAND2_X1 U991 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
INV_X1 U992 ( .A(KEYINPUT52), .ZN(n1286) );
NAND2_X1 U993 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
NAND2_X1 U994 ( .A1(n1289), .A2(n1067), .ZN(n1288) );
INV_X1 U995 ( .A(n1063), .ZN(n1287) );
NOR2_X1 U996 ( .A1(n1067), .A2(n1289), .ZN(n1063) );
NAND2_X1 U997 ( .A1(KEYINPUT52), .A2(n1290), .ZN(n1283) );
XNOR2_X1 U998 ( .A(n1067), .B(n1065), .ZN(n1290) );
INV_X1 U999 ( .A(n1289), .ZN(n1065) );
XOR2_X1 U1000 ( .A(G478), .B(KEYINPUT30), .Z(n1289) );
NAND2_X1 U1001 ( .A1(n1291), .A2(n1224), .ZN(n1067) );
XOR2_X1 U1002 ( .A(n1122), .B(KEYINPUT59), .Z(n1291) );
XOR2_X1 U1003 ( .A(n1292), .B(n1293), .Z(n1122) );
XOR2_X1 U1004 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1005 ( .A1(G128), .A2(KEYINPUT41), .ZN(n1295) );
AND3_X1 U1006 ( .A1(G217), .A2(n1012), .A3(G234), .ZN(n1294) );
XOR2_X1 U1007 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U1008 ( .A(G143), .B(G134), .Z(n1297) );
NAND2_X1 U1009 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
NAND2_X1 U1010 ( .A1(G107), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1011 ( .A(KEYINPUT62), .B(n1301), .Z(n1298) );
NOR2_X1 U1012 ( .A1(G107), .A2(n1300), .ZN(n1301) );
XNOR2_X1 U1013 ( .A(n1260), .B(n1302), .ZN(n1300) );
NOR2_X1 U1014 ( .A1(KEYINPUT15), .A2(n1303), .ZN(n1302) );
INV_X1 U1015 ( .A(G122), .ZN(n1260) );
XOR2_X1 U1016 ( .A(KEYINPUT23), .B(n1029), .Z(n1221) );
NOR2_X1 U1017 ( .A1(n1057), .A2(n1219), .ZN(n1029) );
INV_X1 U1018 ( .A(n1203), .ZN(n1219) );
NAND2_X1 U1019 ( .A1(n1076), .A2(n1061), .ZN(n1203) );
NAND3_X1 U1020 ( .A1(n1224), .A2(n1304), .A3(n1117), .ZN(n1061) );
NAND2_X1 U1021 ( .A1(G217), .A2(n1238), .ZN(n1304) );
NAND3_X1 U1022 ( .A1(n1238), .A2(n1305), .A3(G217), .ZN(n1076) );
NAND2_X1 U1023 ( .A1(n1117), .A2(n1224), .ZN(n1305) );
XOR2_X1 U1024 ( .A(n1306), .B(n1307), .Z(n1117) );
XOR2_X1 U1025 ( .A(G137), .B(n1308), .Z(n1307) );
AND3_X1 U1026 ( .A1(G221), .A2(n1012), .A3(G234), .ZN(n1308) );
INV_X1 U1027 ( .A(G953), .ZN(n1012) );
NAND2_X1 U1028 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
NAND2_X1 U1029 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1030 ( .A(KEYINPUT3), .B(n1313), .Z(n1309) );
NOR2_X1 U1031 ( .A1(n1311), .A2(n1312), .ZN(n1313) );
XOR2_X1 U1032 ( .A(G146), .B(n1101), .Z(n1312) );
XOR2_X1 U1033 ( .A(G125), .B(G140), .Z(n1101) );
XOR2_X1 U1034 ( .A(n1314), .B(n1315), .Z(n1311) );
XNOR2_X1 U1035 ( .A(G128), .B(n1237), .ZN(n1315) );
INV_X1 U1036 ( .A(G110), .ZN(n1237) );
NAND2_X1 U1037 ( .A1(KEYINPUT47), .A2(G119), .ZN(n1314) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1162), .ZN(n1238) );
INV_X1 U1039 ( .A(G902), .ZN(n1162) );
XNOR2_X1 U1040 ( .A(n1316), .B(G472), .ZN(n1057) );
NAND2_X1 U1041 ( .A1(n1317), .A2(n1224), .ZN(n1316) );
XNOR2_X1 U1042 ( .A(G902), .B(KEYINPUT29), .ZN(n1224) );
XNOR2_X1 U1043 ( .A(n1318), .B(n1135), .ZN(n1317) );
XOR2_X1 U1044 ( .A(n1319), .B(n1099), .Z(n1135) );
XNOR2_X1 U1045 ( .A(G128), .B(n1280), .ZN(n1099) );
XOR2_X1 U1046 ( .A(G143), .B(G146), .Z(n1280) );
XNOR2_X1 U1047 ( .A(n1148), .B(n1320), .ZN(n1319) );
NOR2_X1 U1048 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1049 ( .A(n1323), .B(KEYINPUT17), .Z(n1322) );
NAND2_X1 U1050 ( .A1(n1264), .A2(n1267), .ZN(n1323) );
NOR2_X1 U1051 ( .A1(n1267), .A2(n1264), .ZN(n1321) );
XNOR2_X1 U1052 ( .A(G113), .B(KEYINPUT45), .ZN(n1264) );
XOR2_X1 U1053 ( .A(G119), .B(n1303), .Z(n1267) );
INV_X1 U1054 ( .A(G116), .ZN(n1303) );
XNOR2_X1 U1055 ( .A(n1100), .B(KEYINPUT7), .ZN(n1148) );
XNOR2_X1 U1056 ( .A(G131), .B(n1324), .ZN(n1100) );
XOR2_X1 U1057 ( .A(G137), .B(G134), .Z(n1324) );
NAND2_X1 U1058 ( .A1(n1325), .A2(n1326), .ZN(n1318) );
NAND3_X1 U1059 ( .A1(n1327), .A2(n1270), .A3(n1328), .ZN(n1326) );
INV_X1 U1060 ( .A(KEYINPUT31), .ZN(n1328) );
NAND2_X1 U1061 ( .A1(n1130), .A2(KEYINPUT31), .ZN(n1325) );
XOR2_X1 U1062 ( .A(n1327), .B(n1270), .Z(n1130) );
INV_X1 U1063 ( .A(G101), .ZN(n1270) );
NAND2_X1 U1064 ( .A1(n1282), .A2(G210), .ZN(n1327) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1282) );
endmodule


