//Key = 1001110100100110000011011001101111000110100110011001111101110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358;

XNOR2_X1 U753 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U754 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U755 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
NOR2_X1 U756 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U757 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U758 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
INV_X1 U759 ( .A(n1040), .ZN(n1039) );
NOR2_X1 U760 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
NOR2_X1 U761 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U762 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1041) );
NOR2_X1 U763 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U764 ( .A1(n1045), .A2(n1050), .A3(n1044), .ZN(n1036) );
NOR2_X1 U765 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U766 ( .A1(n1053), .A2(n1047), .ZN(n1052) );
NOR2_X1 U767 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U768 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
XNOR2_X1 U769 ( .A(KEYINPUT19), .B(n1058), .ZN(n1057) );
NOR3_X1 U770 ( .A1(n1059), .A2(KEYINPUT33), .A3(n1043), .ZN(n1051) );
AND4_X1 U771 ( .A1(n1040), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1043) );
NAND3_X1 U772 ( .A1(n1063), .A2(n1064), .A3(n1045), .ZN(n1062) );
NAND2_X1 U773 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U774 ( .A1(KEYINPUT33), .A2(n1067), .A3(n1068), .ZN(n1061) );
NAND2_X1 U775 ( .A1(n1068), .A2(n1069), .ZN(n1060) );
NOR3_X1 U776 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U777 ( .A1(n1070), .A2(n1063), .A3(n1071), .A4(n1072), .ZN(n1031) );
NOR4_X1 U778 ( .A1(n1065), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XNOR2_X1 U779 ( .A(n1076), .B(KEYINPUT47), .ZN(n1074) );
XNOR2_X1 U780 ( .A(n1077), .B(n1078), .ZN(n1071) );
XNOR2_X1 U781 ( .A(n1066), .B(KEYINPUT25), .ZN(n1070) );
XOR2_X1 U782 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U783 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XOR2_X1 U785 ( .A(KEYINPUT43), .B(G227), .Z(n1084) );
INV_X1 U786 ( .A(G900), .ZN(n1083) );
NOR2_X1 U787 ( .A1(KEYINPUT34), .A2(n1085), .ZN(n1079) );
XOR2_X1 U788 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U789 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U790 ( .A(n1090), .B(n1091), .Z(n1089) );
XNOR2_X1 U791 ( .A(n1092), .B(KEYINPUT29), .ZN(n1091) );
NAND2_X1 U792 ( .A1(n1093), .A2(KEYINPUT28), .ZN(n1092) );
XNOR2_X1 U793 ( .A(G134), .B(G137), .ZN(n1093) );
XOR2_X1 U794 ( .A(n1094), .B(n1095), .Z(n1090) );
NAND2_X1 U795 ( .A1(n1082), .A2(n1096), .ZN(n1086) );
XOR2_X1 U796 ( .A(n1097), .B(n1098), .Z(G69) );
NOR2_X1 U797 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U798 ( .A(n1101), .B(KEYINPUT14), .Z(n1100) );
NAND2_X1 U799 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR3_X1 U800 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1099) );
NOR2_X1 U801 ( .A1(G898), .A2(n1082), .ZN(n1104) );
AND2_X1 U802 ( .A1(n1105), .A2(n1082), .ZN(n1103) );
NAND2_X1 U803 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U804 ( .A(n1108), .B(n1109), .Z(n1102) );
NAND3_X1 U805 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1108) );
OR2_X1 U806 ( .A1(n1113), .A2(KEYINPUT23), .ZN(n1112) );
NAND3_X1 U807 ( .A1(KEYINPUT23), .A2(n1114), .A3(n1115), .ZN(n1111) );
OR2_X1 U808 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
NOR2_X1 U809 ( .A1(KEYINPUT15), .A2(n1116), .ZN(n1114) );
NAND2_X1 U810 ( .A1(G953), .A2(n1117), .ZN(n1097) );
NAND2_X1 U811 ( .A1(G898), .A2(G224), .ZN(n1117) );
NOR2_X1 U812 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U813 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U814 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR2_X1 U815 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U816 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U817 ( .A(n1127), .B(KEYINPUT1), .Z(n1125) );
NAND2_X1 U818 ( .A1(n1128), .A2(G478), .ZN(n1127) );
NOR2_X1 U819 ( .A1(n1118), .A2(n1129), .ZN(G60) );
NOR2_X1 U820 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U821 ( .A(n1132), .B(n1133), .Z(n1131) );
AND2_X1 U822 ( .A1(G475), .A2(n1128), .ZN(n1133) );
AND2_X1 U823 ( .A1(n1134), .A2(KEYINPUT58), .ZN(n1132) );
NOR2_X1 U824 ( .A1(KEYINPUT58), .A2(n1134), .ZN(n1130) );
XOR2_X1 U825 ( .A(n1135), .B(n1136), .Z(G6) );
NAND2_X1 U826 ( .A1(KEYINPUT7), .A2(n1137), .ZN(n1135) );
INV_X1 U827 ( .A(G104), .ZN(n1137) );
NOR2_X1 U828 ( .A1(n1118), .A2(n1138), .ZN(G57) );
XOR2_X1 U829 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U830 ( .A(n1141), .B(n1142), .Z(n1140) );
AND2_X1 U831 ( .A1(G472), .A2(n1128), .ZN(n1141) );
XOR2_X1 U832 ( .A(n1143), .B(n1144), .Z(n1139) );
NOR3_X1 U833 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
NOR2_X1 U834 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U835 ( .A1(KEYINPUT46), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U836 ( .A(G101), .B(KEYINPUT17), .ZN(n1150) );
NOR3_X1 U837 ( .A1(n1151), .A2(KEYINPUT46), .A3(n1152), .ZN(n1146) );
AND2_X1 U838 ( .A1(n1152), .A2(KEYINPUT46), .ZN(n1145) );
NAND2_X1 U839 ( .A1(n1153), .A2(n1154), .ZN(n1143) );
NAND2_X1 U840 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U841 ( .A(KEYINPUT31), .B(n1157), .Z(n1153) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1156), .ZN(n1157) );
NOR2_X1 U843 ( .A1(n1118), .A2(n1158), .ZN(G54) );
XOR2_X1 U844 ( .A(n1159), .B(n1160), .Z(n1158) );
XNOR2_X1 U845 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U846 ( .A(G140), .B(G110), .Z(n1162) );
XOR2_X1 U847 ( .A(n1163), .B(n1164), .Z(n1159) );
AND2_X1 U848 ( .A1(G469), .A2(n1128), .ZN(n1164) );
NAND3_X1 U849 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1163) );
OR2_X1 U850 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U851 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
INV_X1 U852 ( .A(KEYINPUT40), .ZN(n1171) );
NAND2_X1 U853 ( .A1(n1172), .A2(n1169), .ZN(n1170) );
XNOR2_X1 U854 ( .A(KEYINPUT59), .B(n1168), .ZN(n1172) );
NAND2_X1 U855 ( .A1(KEYINPUT40), .A2(n1173), .ZN(n1165) );
NAND2_X1 U856 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
OR2_X1 U857 ( .A1(n1168), .A2(KEYINPUT59), .ZN(n1175) );
NAND3_X1 U858 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT59), .ZN(n1174) );
XNOR2_X1 U859 ( .A(n1176), .B(KEYINPUT35), .ZN(n1169) );
NOR2_X1 U860 ( .A1(n1118), .A2(n1177), .ZN(G51) );
XOR2_X1 U861 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U862 ( .A(n1180), .B(n1181), .ZN(n1179) );
XNOR2_X1 U863 ( .A(n1182), .B(n1183), .ZN(n1178) );
XOR2_X1 U864 ( .A(n1184), .B(KEYINPUT26), .Z(n1183) );
NAND2_X1 U865 ( .A1(n1128), .A2(n1185), .ZN(n1184) );
INV_X1 U866 ( .A(n1123), .ZN(n1128) );
NAND2_X1 U867 ( .A1(G902), .A2(n1033), .ZN(n1123) );
NAND3_X1 U868 ( .A1(n1106), .A2(n1186), .A3(n1187), .ZN(n1033) );
INV_X1 U869 ( .A(n1096), .ZN(n1187) );
NAND4_X1 U870 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1096) );
NOR4_X1 U871 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NAND2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
NAND2_X1 U873 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U874 ( .A1(n1049), .A2(n1067), .ZN(n1199) );
INV_X1 U875 ( .A(n1200), .ZN(n1049) );
XNOR2_X1 U876 ( .A(KEYINPUT38), .B(n1107), .ZN(n1186) );
AND4_X1 U877 ( .A1(n1201), .A2(n1028), .A3(n1202), .A4(n1203), .ZN(n1106) );
NOR3_X1 U878 ( .A1(n1204), .A2(n1136), .A3(n1205), .ZN(n1203) );
NOR3_X1 U879 ( .A1(n1206), .A2(n1207), .A3(n1047), .ZN(n1205) );
AND2_X1 U880 ( .A1(n1067), .A2(n1208), .ZN(n1136) );
NOR2_X1 U881 ( .A1(n1209), .A2(n1210), .ZN(n1204) );
NOR2_X1 U882 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
XOR2_X1 U883 ( .A(n1213), .B(KEYINPUT24), .Z(n1212) );
NOR2_X1 U884 ( .A1(n1214), .A2(n1198), .ZN(n1211) );
NAND2_X1 U885 ( .A1(n1069), .A2(n1208), .ZN(n1028) );
NOR2_X1 U886 ( .A1(n1207), .A2(n1044), .ZN(n1208) );
INV_X1 U887 ( .A(n1215), .ZN(n1044) );
NOR2_X1 U888 ( .A1(n1082), .A2(G952), .ZN(n1118) );
XNOR2_X1 U889 ( .A(G146), .B(n1188), .ZN(G48) );
NAND2_X1 U890 ( .A1(n1216), .A2(n1067), .ZN(n1188) );
XNOR2_X1 U891 ( .A(G143), .B(n1189), .ZN(G45) );
NAND3_X1 U892 ( .A1(n1048), .A2(n1217), .A3(n1218), .ZN(n1189) );
XOR2_X1 U893 ( .A(G140), .B(n1219), .Z(G42) );
NOR3_X1 U894 ( .A1(n1220), .A2(n1200), .A3(n1221), .ZN(n1219) );
XNOR2_X1 U895 ( .A(KEYINPUT52), .B(n1059), .ZN(n1220) );
XOR2_X1 U896 ( .A(n1222), .B(n1223), .Z(G39) );
XNOR2_X1 U897 ( .A(G137), .B(KEYINPUT45), .ZN(n1223) );
NAND3_X1 U898 ( .A1(n1224), .A2(n1196), .A3(KEYINPUT63), .ZN(n1222) );
INV_X1 U899 ( .A(n1198), .ZN(n1224) );
XOR2_X1 U900 ( .A(G134), .B(n1195), .Z(G36) );
AND3_X1 U901 ( .A1(n1196), .A2(n1069), .A3(n1048), .ZN(n1195) );
INV_X1 U902 ( .A(n1221), .ZN(n1196) );
XNOR2_X1 U903 ( .A(n1194), .B(n1225), .ZN(G33) );
NAND2_X1 U904 ( .A1(KEYINPUT48), .A2(G131), .ZN(n1225) );
NOR3_X1 U905 ( .A1(n1221), .A2(n1059), .A3(n1206), .ZN(n1194) );
NAND2_X1 U906 ( .A1(n1040), .A2(n1217), .ZN(n1221) );
NOR2_X1 U907 ( .A1(n1076), .A2(n1073), .ZN(n1040) );
XOR2_X1 U908 ( .A(G128), .B(n1193), .Z(G30) );
AND2_X1 U909 ( .A1(n1216), .A2(n1069), .ZN(n1193) );
AND4_X1 U910 ( .A1(n1217), .A2(n1055), .A3(n1075), .A4(n1226), .ZN(n1216) );
AND3_X1 U911 ( .A1(n1227), .A2(n1228), .A3(n1066), .ZN(n1217) );
NAND2_X1 U912 ( .A1(n1229), .A2(n1230), .ZN(G3) );
OR2_X1 U913 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U914 ( .A1(n1232), .A2(n1233), .ZN(n1229) );
NAND2_X1 U915 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U916 ( .A1(KEYINPUT57), .A2(n1231), .ZN(n1235) );
OR2_X1 U917 ( .A1(KEYINPUT9), .A2(n1236), .ZN(n1231) );
OR2_X1 U918 ( .A1(n1236), .A2(KEYINPUT57), .ZN(n1234) );
XOR2_X1 U919 ( .A(G101), .B(KEYINPUT30), .Z(n1236) );
NOR3_X1 U920 ( .A1(n1047), .A2(n1207), .A3(n1237), .ZN(n1232) );
XNOR2_X1 U921 ( .A(n1206), .B(KEYINPUT4), .ZN(n1237) );
INV_X1 U922 ( .A(n1048), .ZN(n1206) );
XNOR2_X1 U923 ( .A(n1238), .B(n1192), .ZN(G27) );
AND4_X1 U924 ( .A1(n1055), .A2(n1227), .A3(n1067), .A4(n1239), .ZN(n1192) );
NOR2_X1 U925 ( .A1(n1045), .A2(n1200), .ZN(n1239) );
INV_X1 U926 ( .A(n1068), .ZN(n1045) );
NAND2_X1 U927 ( .A1(n1240), .A2(n1035), .ZN(n1227) );
NAND3_X1 U928 ( .A1(G902), .A2(n1241), .A3(n1088), .ZN(n1240) );
NOR2_X1 U929 ( .A1(n1082), .A2(G900), .ZN(n1088) );
NAND2_X1 U930 ( .A1(n1242), .A2(n1243), .ZN(G24) );
OR2_X1 U931 ( .A1(n1202), .A2(G122), .ZN(n1243) );
XOR2_X1 U932 ( .A(n1244), .B(KEYINPUT60), .Z(n1242) );
NAND2_X1 U933 ( .A1(G122), .A2(n1202), .ZN(n1244) );
NAND3_X1 U934 ( .A1(n1218), .A2(n1215), .A3(n1245), .ZN(n1202) );
NOR2_X1 U935 ( .A1(n1226), .A2(n1075), .ZN(n1215) );
AND3_X1 U936 ( .A1(n1246), .A2(n1247), .A3(n1055), .ZN(n1218) );
XOR2_X1 U937 ( .A(G119), .B(n1248), .Z(G21) );
NOR3_X1 U938 ( .A1(n1249), .A2(n1214), .A3(n1198), .ZN(n1248) );
NAND3_X1 U939 ( .A1(n1075), .A2(n1226), .A3(n1063), .ZN(n1198) );
XNOR2_X1 U940 ( .A(KEYINPUT10), .B(n1210), .ZN(n1249) );
XNOR2_X1 U941 ( .A(n1250), .B(n1251), .ZN(G18) );
NOR3_X1 U942 ( .A1(n1213), .A2(KEYINPUT6), .A3(n1210), .ZN(n1251) );
INV_X1 U943 ( .A(n1055), .ZN(n1210) );
NAND3_X1 U944 ( .A1(n1048), .A2(n1069), .A3(n1245), .ZN(n1213) );
NOR2_X1 U945 ( .A1(n1246), .A2(n1252), .ZN(n1069) );
XNOR2_X1 U946 ( .A(G113), .B(n1201), .ZN(G15) );
NAND4_X1 U947 ( .A1(n1245), .A2(n1048), .A3(n1067), .A4(n1055), .ZN(n1201) );
INV_X1 U948 ( .A(n1059), .ZN(n1067) );
NAND2_X1 U949 ( .A1(n1252), .A2(n1246), .ZN(n1059) );
INV_X1 U950 ( .A(n1247), .ZN(n1252) );
NOR2_X1 U951 ( .A1(n1226), .A2(n1253), .ZN(n1048) );
INV_X1 U952 ( .A(n1214), .ZN(n1245) );
NAND2_X1 U953 ( .A1(n1068), .A2(n1254), .ZN(n1214) );
NOR2_X1 U954 ( .A1(n1066), .A2(n1065), .ZN(n1068) );
INV_X1 U955 ( .A(n1228), .ZN(n1065) );
XNOR2_X1 U956 ( .A(G110), .B(n1107), .ZN(G12) );
OR3_X1 U957 ( .A1(n1047), .A2(n1207), .A3(n1200), .ZN(n1107) );
NAND2_X1 U958 ( .A1(n1253), .A2(n1226), .ZN(n1200) );
NAND3_X1 U959 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1226) );
NAND2_X1 U960 ( .A1(KEYINPUT8), .A2(n1077), .ZN(n1257) );
NAND3_X1 U961 ( .A1(n1258), .A2(n1259), .A3(n1078), .ZN(n1256) );
INV_X1 U962 ( .A(n1122), .ZN(n1078) );
NAND2_X1 U963 ( .A1(n1260), .A2(n1122), .ZN(n1255) );
NAND2_X1 U964 ( .A1(G217), .A2(n1261), .ZN(n1122) );
NAND2_X1 U965 ( .A1(n1262), .A2(n1259), .ZN(n1260) );
INV_X1 U966 ( .A(KEYINPUT8), .ZN(n1259) );
XNOR2_X1 U967 ( .A(n1077), .B(KEYINPUT16), .ZN(n1262) );
INV_X1 U968 ( .A(n1258), .ZN(n1077) );
NAND2_X1 U969 ( .A1(n1263), .A2(n1264), .ZN(n1258) );
XNOR2_X1 U970 ( .A(n1121), .B(KEYINPUT61), .ZN(n1263) );
XNOR2_X1 U971 ( .A(n1265), .B(n1266), .ZN(n1121) );
XOR2_X1 U972 ( .A(G137), .B(n1267), .Z(n1266) );
NOR2_X1 U973 ( .A1(KEYINPUT36), .A2(n1268), .ZN(n1267) );
XOR2_X1 U974 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U975 ( .A(G110), .B(n1271), .Z(n1270) );
XOR2_X1 U976 ( .A(G119), .B(n1272), .Z(n1269) );
XOR2_X1 U977 ( .A(G146), .B(G128), .Z(n1272) );
NAND3_X1 U978 ( .A1(G234), .A2(n1082), .A3(G221), .ZN(n1265) );
INV_X1 U979 ( .A(n1075), .ZN(n1253) );
XNOR2_X1 U980 ( .A(n1273), .B(G472), .ZN(n1075) );
NAND2_X1 U981 ( .A1(n1274), .A2(n1264), .ZN(n1273) );
XOR2_X1 U982 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U983 ( .A(n1277), .B(n1156), .ZN(n1276) );
INV_X1 U984 ( .A(n1182), .ZN(n1156) );
XNOR2_X1 U985 ( .A(n1142), .B(n1148), .ZN(n1277) );
INV_X1 U986 ( .A(n1151), .ZN(n1148) );
NAND2_X1 U987 ( .A1(G210), .A2(n1278), .ZN(n1151) );
XNOR2_X1 U988 ( .A(n1279), .B(n1280), .ZN(n1142) );
XOR2_X1 U989 ( .A(KEYINPUT51), .B(G119), .Z(n1280) );
XNOR2_X1 U990 ( .A(G116), .B(n1281), .ZN(n1279) );
XOR2_X1 U991 ( .A(n1282), .B(n1283), .Z(n1275) );
XNOR2_X1 U992 ( .A(KEYINPUT27), .B(n1152), .ZN(n1283) );
NAND2_X1 U993 ( .A1(KEYINPUT5), .A2(n1155), .ZN(n1282) );
NAND4_X1 U994 ( .A1(n1055), .A2(n1066), .A3(n1254), .A4(n1228), .ZN(n1207) );
NAND2_X1 U995 ( .A1(G221), .A2(n1261), .ZN(n1228) );
NAND2_X1 U996 ( .A1(G234), .A2(n1264), .ZN(n1261) );
NAND2_X1 U997 ( .A1(n1035), .A2(n1284), .ZN(n1254) );
NAND4_X1 U998 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1285), .ZN(n1284) );
INV_X1 U999 ( .A(G898), .ZN(n1285) );
NAND3_X1 U1000 ( .A1(n1241), .A2(n1082), .A3(G952), .ZN(n1035) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1241) );
XNOR2_X1 U1002 ( .A(n1286), .B(G469), .ZN(n1066) );
NAND3_X1 U1003 ( .A1(n1287), .A2(n1288), .A3(n1264), .ZN(n1286) );
NAND2_X1 U1004 ( .A1(n1289), .A2(n1161), .ZN(n1288) );
XOR2_X1 U1005 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U1006 ( .A1(KEYINPUT3), .A2(n1292), .ZN(n1291) );
NAND2_X1 U1007 ( .A1(n1293), .A2(n1294), .ZN(n1287) );
INV_X1 U1008 ( .A(n1161), .ZN(n1294) );
NAND2_X1 U1009 ( .A1(G227), .A2(n1082), .ZN(n1161) );
XOR2_X1 U1010 ( .A(n1290), .B(n1295), .Z(n1293) );
NAND2_X1 U1011 ( .A1(KEYINPUT3), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U1012 ( .A(KEYINPUT42), .B(n1292), .ZN(n1296) );
XNOR2_X1 U1013 ( .A(G140), .B(n1297), .ZN(n1292) );
NOR2_X1 U1014 ( .A1(G110), .A2(KEYINPUT22), .ZN(n1297) );
NAND3_X1 U1015 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1290) );
OR2_X1 U1016 ( .A1(n1301), .A2(KEYINPUT13), .ZN(n1300) );
INV_X1 U1017 ( .A(n1176), .ZN(n1301) );
NAND3_X1 U1018 ( .A1(KEYINPUT13), .A2(n1302), .A3(n1155), .ZN(n1299) );
OR2_X1 U1019 ( .A1(n1155), .A2(n1302), .ZN(n1298) );
NOR2_X1 U1020 ( .A1(KEYINPUT2), .A2(n1176), .ZN(n1302) );
XNOR2_X1 U1021 ( .A(n1303), .B(n1095), .ZN(n1176) );
XNOR2_X1 U1022 ( .A(n1304), .B(n1305), .ZN(n1095) );
NAND3_X1 U1023 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1303) );
NAND2_X1 U1024 ( .A1(n1309), .A2(G101), .ZN(n1307) );
NAND2_X1 U1025 ( .A1(n1310), .A2(n1152), .ZN(n1306) );
XNOR2_X1 U1026 ( .A(G104), .B(G107), .ZN(n1310) );
INV_X1 U1027 ( .A(n1168), .ZN(n1155) );
XNOR2_X1 U1028 ( .A(n1311), .B(n1312), .ZN(n1168) );
XOR2_X1 U1029 ( .A(KEYINPUT21), .B(G131), .Z(n1312) );
NAND2_X1 U1030 ( .A1(KEYINPUT55), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1031 ( .A(G137), .B(G134), .Z(n1313) );
NOR2_X1 U1032 ( .A1(n1058), .A2(n1073), .ZN(n1055) );
INV_X1 U1033 ( .A(n1056), .ZN(n1073) );
NAND2_X1 U1034 ( .A1(G214), .A2(n1314), .ZN(n1056) );
INV_X1 U1035 ( .A(n1076), .ZN(n1058) );
XNOR2_X1 U1036 ( .A(n1315), .B(n1185), .ZN(n1076) );
AND2_X1 U1037 ( .A1(G210), .A2(n1314), .ZN(n1185) );
NAND2_X1 U1038 ( .A1(n1316), .A2(n1264), .ZN(n1314) );
XNOR2_X1 U1039 ( .A(G237), .B(KEYINPUT50), .ZN(n1316) );
NAND2_X1 U1040 ( .A1(n1317), .A2(n1264), .ZN(n1315) );
XOR2_X1 U1041 ( .A(n1318), .B(n1180), .Z(n1317) );
XOR2_X1 U1042 ( .A(n1319), .B(n1320), .Z(n1180) );
XNOR2_X1 U1043 ( .A(n1115), .B(n1321), .ZN(n1320) );
NAND2_X1 U1044 ( .A1(G224), .A2(n1082), .ZN(n1321) );
INV_X1 U1045 ( .A(G953), .ZN(n1082) );
AND3_X1 U1046 ( .A1(n1322), .A2(n1323), .A3(n1308), .ZN(n1115) );
NAND3_X1 U1047 ( .A1(G104), .A2(n1324), .A3(G101), .ZN(n1308) );
NAND3_X1 U1048 ( .A1(n1325), .A2(n1326), .A3(n1152), .ZN(n1323) );
INV_X1 U1049 ( .A(G101), .ZN(n1152) );
NAND2_X1 U1050 ( .A1(G104), .A2(n1324), .ZN(n1326) );
XNOR2_X1 U1051 ( .A(n1309), .B(KEYINPUT39), .ZN(n1325) );
NAND2_X1 U1052 ( .A1(n1327), .A2(G101), .ZN(n1322) );
XNOR2_X1 U1053 ( .A(KEYINPUT39), .B(n1328), .ZN(n1327) );
INV_X1 U1054 ( .A(n1309), .ZN(n1328) );
NOR2_X1 U1055 ( .A1(n1324), .A2(G104), .ZN(n1309) );
XNOR2_X1 U1056 ( .A(n1116), .B(n1109), .ZN(n1319) );
XOR2_X1 U1057 ( .A(G110), .B(n1329), .Z(n1109) );
XOR2_X1 U1058 ( .A(KEYINPUT41), .B(G122), .Z(n1329) );
INV_X1 U1059 ( .A(n1113), .ZN(n1116) );
NAND2_X1 U1060 ( .A1(n1330), .A2(n1331), .ZN(n1113) );
NAND2_X1 U1061 ( .A1(n1332), .A2(n1250), .ZN(n1331) );
XOR2_X1 U1062 ( .A(KEYINPUT11), .B(n1333), .Z(n1332) );
NAND2_X1 U1063 ( .A1(n1334), .A2(G116), .ZN(n1330) );
XOR2_X1 U1064 ( .A(KEYINPUT20), .B(n1333), .Z(n1334) );
XOR2_X1 U1065 ( .A(G119), .B(n1281), .Z(n1333) );
NAND2_X1 U1066 ( .A1(n1335), .A2(KEYINPUT62), .ZN(n1318) );
XNOR2_X1 U1067 ( .A(n1182), .B(n1336), .ZN(n1335) );
XOR2_X1 U1068 ( .A(KEYINPUT0), .B(n1337), .Z(n1336) );
NOR2_X1 U1069 ( .A1(KEYINPUT56), .A2(n1181), .ZN(n1337) );
XOR2_X1 U1070 ( .A(G125), .B(KEYINPUT18), .Z(n1181) );
XNOR2_X1 U1071 ( .A(n1338), .B(n1305), .ZN(n1182) );
XOR2_X1 U1072 ( .A(G128), .B(KEYINPUT12), .Z(n1305) );
NAND2_X1 U1073 ( .A1(KEYINPUT32), .A2(n1304), .ZN(n1338) );
INV_X1 U1074 ( .A(n1063), .ZN(n1047) );
NOR2_X1 U1075 ( .A1(n1247), .A2(n1246), .ZN(n1063) );
XNOR2_X1 U1076 ( .A(n1339), .B(G475), .ZN(n1246) );
NAND2_X1 U1077 ( .A1(n1134), .A2(n1264), .ZN(n1339) );
XOR2_X1 U1078 ( .A(n1340), .B(n1341), .Z(n1134) );
XOR2_X1 U1079 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1080 ( .A(G122), .B(G104), .ZN(n1343) );
NAND2_X1 U1081 ( .A1(G214), .A2(n1278), .ZN(n1342) );
NOR2_X1 U1082 ( .A1(G953), .A2(G237), .ZN(n1278) );
XOR2_X1 U1083 ( .A(n1094), .B(n1344), .Z(n1340) );
XNOR2_X1 U1084 ( .A(n1281), .B(n1304), .ZN(n1344) );
XNOR2_X1 U1085 ( .A(G143), .B(G146), .ZN(n1304) );
XOR2_X1 U1086 ( .A(G113), .B(KEYINPUT53), .Z(n1281) );
XNOR2_X1 U1087 ( .A(G131), .B(n1271), .ZN(n1094) );
XNOR2_X1 U1088 ( .A(n1238), .B(G140), .ZN(n1271) );
INV_X1 U1089 ( .A(G125), .ZN(n1238) );
XNOR2_X1 U1090 ( .A(n1345), .B(G478), .ZN(n1247) );
NAND2_X1 U1091 ( .A1(n1126), .A2(n1264), .ZN(n1345) );
INV_X1 U1092 ( .A(G902), .ZN(n1264) );
XNOR2_X1 U1093 ( .A(n1346), .B(n1347), .ZN(n1126) );
NOR3_X1 U1094 ( .A1(n1348), .A2(G953), .A3(n1349), .ZN(n1347) );
INV_X1 U1095 ( .A(G217), .ZN(n1349) );
XOR2_X1 U1096 ( .A(KEYINPUT44), .B(G234), .Z(n1348) );
NAND2_X1 U1097 ( .A1(n1350), .A2(KEYINPUT54), .ZN(n1346) );
XOR2_X1 U1098 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1099 ( .A(G122), .B(n1250), .ZN(n1352) );
INV_X1 U1100 ( .A(G116), .ZN(n1250) );
XNOR2_X1 U1101 ( .A(n1353), .B(n1324), .ZN(n1351) );
INV_X1 U1102 ( .A(G107), .ZN(n1324) );
NAND3_X1 U1103 ( .A1(n1354), .A2(n1355), .A3(KEYINPUT37), .ZN(n1353) );
NAND2_X1 U1104 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1105 ( .A(G134), .B(n1358), .Z(n1356) );
OR3_X1 U1106 ( .A1(n1358), .A2(G134), .A3(n1357), .ZN(n1354) );
INV_X1 U1107 ( .A(KEYINPUT49), .ZN(n1357) );
XOR2_X1 U1108 ( .A(G143), .B(G128), .Z(n1358) );
endmodule


