//Key = 1111111111111111011011111010110110111110011111
module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, 
        G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, 
        G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, 
        KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, 
        KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, 
        KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, 
        KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, 
        KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, 
        KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, 
        KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, 
        KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, G3, G6, G9, G12, G30, 
        G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
        G60, G63, G66, G69, G72, G57 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
         KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
         KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
         KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
         KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
         KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
         KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
         KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
         KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
         KEYINPUT43, KEYINPUT44, KEYINPUT45;
         
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932;

  NAND2_X1 U520 ( .A1(n707), .A2(KEYINPUT10), .ZN(G9) );
  XNOR2_X1 U521 ( .A(n708), .B(G107), .ZN(n707) );
  NOR2_X1 U522 ( .A1(n709), .A2(n710), .ZN(G75) );
  NOR2_X1 U523 ( .A1(G952), .A2(n711), .ZN(n710) );
  NOR2_X1 U524 ( .A1(n712), .A2(n713), .ZN(n709) );
  NAND4_X1 U525 ( .A1(KEYINPUT43), .A2(KEYINPUT36), .A3(KEYINPUT26), .A4(KEYINPUT22), .ZN(n713) );
  NAND4_X1 U526 ( .A1(n714), .A2(n715), .A3(n716), .A4(n717), .ZN(n712) );
  NAND2_X1 U527 ( .A1(n718), .A2(n719), .ZN(n717) );
  NAND2_X1 U528 ( .A1(n720), .A2(n721), .ZN(n719) );
  NAND3_X1 U529 ( .A1(n722), .A2(n723), .A3(n724), .ZN(n721) );
  NAND2_X1 U530 ( .A1(n725), .A2(n726), .ZN(n723) );
  NAND2_X1 U531 ( .A1(n727), .A2(n728), .ZN(n726) );
  NAND2_X1 U532 ( .A1(n729), .A2(n730), .ZN(n728) );
  NAND2_X1 U533 ( .A1(n731), .A2(n732), .ZN(n725) );
  NAND3_X1 U534 ( .A1(n727), .A2(n733), .A3(n731), .ZN(n720) );
  NAND2_X1 U535 ( .A1(n734), .A2(n735), .ZN(n733) );
  NAND2_X1 U536 ( .A1(n724), .A2(n736), .ZN(n735) );
  OR2_X1 U537 ( .A1(n737), .A2(n738), .ZN(n736) );
  NAND2_X1 U538 ( .A1(n722), .A2(n739), .ZN(n734) );
  NAND2_X1 U539 ( .A1(n740), .A2(n741), .ZN(n739) );
  INV_X1 U540 ( .A(n742), .ZN(n718) );
  INV_X1 U541 ( .A(n711), .ZN(n716) );
  NAND2_X1 U542 ( .A1(n743), .A2(n744), .ZN(n711) );
  NAND4_X1 U543 ( .A1(n724), .A2(n731), .A3(n727), .A4(n722), .ZN(n744) );
  XOR2_X1 U544 ( .A(n745), .B(n746), .Z(G72) );
  NOR2_X1 U545 ( .A1(n747), .A2(n743), .ZN(n746) );
  NOR2_X1 U546 ( .A1(n748), .A2(n749), .ZN(n747) );
  NAND2_X1 U547 ( .A1(n750), .A2(n751), .ZN(n745) );
  NAND2_X1 U548 ( .A1(n752), .A2(n743), .ZN(n751) );
  XOR2_X1 U549 ( .A(n715), .B(n753), .Z(n752) );
  OR3_X1 U550 ( .A1(n749), .A2(n753), .A3(n743), .ZN(n750) );
  XOR2_X1 U551 ( .A(n754), .B(n755), .Z(n753) );
  XOR2_X1 U552 ( .A(n756), .B(n757), .Z(G69) );
  NOR2_X1 U553 ( .A1(n758), .A2(n743), .ZN(n757) );
  NOR2_X1 U554 ( .A1(n759), .A2(n760), .ZN(n758) );
  NAND2_X1 U555 ( .A1(n761), .A2(n762), .ZN(n756) );
  NAND2_X1 U556 ( .A1(n763), .A2(n743), .ZN(n762) );
  XNOR2_X1 U557 ( .A(n714), .B(n764), .ZN(n763) );
  NAND3_X1 U558 ( .A1(G898), .A2(n764), .A3(G953), .ZN(n761) );
  NOR2_X1 U559 ( .A1(n765), .A2(n766), .ZN(G66) );
  XNOR2_X1 U560 ( .A(n767), .B(n768), .ZN(n766) );
  NOR2_X1 U561 ( .A1(n769), .A2(n770), .ZN(n768) );
  NOR2_X1 U562 ( .A1(n765), .A2(n771), .ZN(G63) );
  XNOR2_X1 U563 ( .A(n772), .B(n773), .ZN(n771) );
  NOR2_X1 U564 ( .A1(n774), .A2(n770), .ZN(n773) );
  NOR2_X1 U565 ( .A1(n765), .A2(n775), .ZN(G60) );
  XNOR2_X1 U566 ( .A(n776), .B(n777), .ZN(n775) );
  NOR2_X1 U567 ( .A1(n778), .A2(n770), .ZN(n777) );
  NAND2_X1 U568 ( .A1(n779), .A2(KEYINPUT9), .ZN(G6) );
  XOR2_X1 U569 ( .A(n780), .B(G104), .Z(n779) );
  NOR2_X1 U570 ( .A1(n765), .A2(n781), .ZN(G57) );
  XNOR2_X1 U571 ( .A(n782), .B(n783), .ZN(n781) );
  NOR2_X1 U572 ( .A1(n784), .A2(n770), .ZN(n783) );
  NOR2_X1 U573 ( .A1(n765), .A2(n785), .ZN(G54) );
  XNOR2_X1 U574 ( .A(n786), .B(n787), .ZN(n785) );
  NOR2_X1 U575 ( .A1(n788), .A2(n770), .ZN(n787) );
  NOR2_X1 U576 ( .A1(n765), .A2(n789), .ZN(G51) );
  XNOR2_X1 U577 ( .A(n790), .B(n791), .ZN(n789) );
  NOR2_X1 U578 ( .A1(n792), .A2(n770), .ZN(n791) );
  NAND2_X1 U579 ( .A1(G902), .A2(n793), .ZN(n770) );
  NAND2_X1 U580 ( .A1(n714), .A2(n715), .ZN(n793) );
  NOR4_X1 U581 ( .A1(n794), .A2(n795), .A3(n796), .A4(n797), .ZN(n715) );
  NAND3_X1 U582 ( .A1(n798), .A2(n799), .A3(n800), .ZN(n797) );
  NAND2_X1 U583 ( .A1(n801), .A2(n732), .ZN(n800) );
  NAND2_X1 U584 ( .A1(n802), .A2(n803), .ZN(n732) );
  INV_X1 U585 ( .A(n804), .ZN(n801) );
  NAND4_X1 U586 ( .A1(n805), .A2(n806), .A3(n807), .A4(n808), .ZN(n796) );
  NAND3_X1 U587 ( .A1(KEYINPUT37), .A2(KEYINPUT34), .A3(KEYINPUT41), .ZN(n795) );
  NAND3_X1 U588 ( .A1(KEYINPUT20), .A2(KEYINPUT17), .A3(KEYINPUT23), .ZN(n794) );
  AND4_X1 U589 ( .A1(KEYINPUT44), .A2(KEYINPUT31), .A3(n809), .A4(n810), .ZN(n714) );
  NOR4_X1 U590 ( .A1(n811), .A2(n708), .A3(n812), .A4(n813), .ZN(n810) );
  AND3_X1 U591 ( .A1(n814), .A2(n722), .A3(n815), .ZN(n708) );
  NAND3_X1 U592 ( .A1(n816), .A2(n817), .A3(n818), .ZN(n811) );
  AND3_X1 U593 ( .A1(n780), .A2(n819), .A3(KEYINPUT28), .ZN(n809) );
  NAND3_X1 U594 ( .A1(n815), .A2(n722), .A3(n820), .ZN(n780) );
  NOR2_X1 U595 ( .A1(n743), .A2(G952), .ZN(n765) );
  NAND3_X1 U596 ( .A1(n821), .A2(n822), .A3(KEYINPUT0), .ZN(G48) );
  OR2_X1 U597 ( .A1(n823), .A2(G146), .ZN(n822) );
  NAND3_X1 U598 ( .A1(KEYINPUT18), .A2(n823), .A3(G146), .ZN(n821) );
  NOR2_X1 U599 ( .A1(n824), .A2(KEYINPUT16), .ZN(n823) );
  NOR2_X1 U600 ( .A1(n802), .A2(n804), .ZN(n824) );
  NAND3_X1 U601 ( .A1(n825), .A2(n826), .A3(KEYINPUT2), .ZN(G45) );
  OR2_X1 U602 ( .A1(n827), .A2(G143), .ZN(n826) );
  NAND3_X1 U603 ( .A1(KEYINPUT24), .A2(n827), .A3(G143), .ZN(n825) );
  NOR2_X1 U604 ( .A1(n828), .A2(KEYINPUT25), .ZN(n827) );
  INV_X1 U605 ( .A(n798), .ZN(n828) );
  NAND4_X1 U606 ( .A1(n829), .A2(n830), .A3(n737), .A4(n831), .ZN(n798) );
  AND3_X1 U607 ( .A1(n832), .A2(n833), .A3(n834), .ZN(n831) );
  NAND3_X1 U608 ( .A1(n835), .A2(n836), .A3(KEYINPUT7), .ZN(G42) );
  OR2_X1 U609 ( .A1(n837), .A2(G140), .ZN(n836) );
  NAND3_X1 U610 ( .A1(KEYINPUT42), .A2(n837), .A3(G140), .ZN(n835) );
  NOR2_X1 U611 ( .A1(n838), .A2(KEYINPUT40), .ZN(n837) );
  INV_X1 U612 ( .A(n808), .ZN(n838) );
  NAND3_X1 U613 ( .A1(n820), .A2(n738), .A3(n839), .ZN(n808) );
  NAND3_X1 U614 ( .A1(n840), .A2(n841), .A3(KEYINPUT6), .ZN(G39) );
  OR2_X1 U615 ( .A1(n842), .A2(G137), .ZN(n841) );
  NAND3_X1 U616 ( .A1(KEYINPUT38), .A2(n842), .A3(G137), .ZN(n840) );
  NOR2_X1 U617 ( .A1(n843), .A2(KEYINPUT39), .ZN(n842) );
  INV_X1 U618 ( .A(n807), .ZN(n843) );
  NAND2_X1 U619 ( .A1(n839), .A2(n844), .ZN(n807) );
  NAND2_X1 U620 ( .A1(n845), .A2(KEYINPUT15), .ZN(G36) );
  XOR2_X1 U621 ( .A(G134), .B(n799), .Z(n845) );
  NAND3_X1 U622 ( .A1(n737), .A2(n814), .A3(n839), .ZN(n799) );
  NAND2_X1 U623 ( .A1(n846), .A2(KEYINPUT14), .ZN(G33) );
  XOR2_X1 U624 ( .A(G131), .B(n805), .Z(n846) );
  NAND3_X1 U625 ( .A1(n737), .A2(n820), .A3(n839), .ZN(n805) );
  AND3_X1 U626 ( .A1(n829), .A2(n833), .A3(n724), .ZN(n839) );
  NOR2_X1 U627 ( .A1(n740), .A2(n847), .ZN(n724) );
  AND2_X1 U628 ( .A1(G214), .A2(n848), .ZN(n847) );
  NAND3_X1 U629 ( .A1(n849), .A2(n850), .A3(KEYINPUT1), .ZN(G30) );
  OR2_X1 U630 ( .A1(n851), .A2(G128), .ZN(n850) );
  NAND3_X1 U631 ( .A1(KEYINPUT21), .A2(n851), .A3(G128), .ZN(n849) );
  NOR2_X1 U632 ( .A1(n852), .A2(KEYINPUT19), .ZN(n851) );
  NOR2_X1 U633 ( .A1(n803), .A2(n804), .ZN(n852) );
  NAND3_X1 U634 ( .A1(n829), .A2(n853), .A3(n854), .ZN(n804) );
  INV_X1 U635 ( .A(n814), .ZN(n803) );
  NAND3_X1 U636 ( .A1(n855), .A2(n856), .A3(KEYINPUT8), .ZN(G3) );
  NAND3_X1 U637 ( .A1(KEYINPUT45), .A2(G101), .A3(n819), .ZN(n856) );
  OR2_X1 U638 ( .A1(n819), .A2(G101), .ZN(n855) );
  NAND3_X1 U639 ( .A1(n727), .A2(n815), .A3(n737), .ZN(n819) );
  NAND3_X1 U640 ( .A1(n857), .A2(n858), .A3(KEYINPUT5), .ZN(G27) );
  OR2_X1 U641 ( .A1(n859), .A2(G125), .ZN(n858) );
  NAND3_X1 U642 ( .A1(KEYINPUT35), .A2(n859), .A3(G125), .ZN(n857) );
  NOR2_X1 U643 ( .A1(n860), .A2(KEYINPUT33), .ZN(n859) );
  INV_X1 U644 ( .A(n806), .ZN(n860) );
  NAND4_X1 U645 ( .A1(n854), .A2(n820), .A3(n861), .A4(n731), .ZN(n806) );
  AND3_X1 U646 ( .A1(n862), .A2(n833), .A3(n830), .ZN(n854) );
  NAND2_X1 U647 ( .A1(n742), .A2(n863), .ZN(n833) );
  NAND4_X1 U648 ( .A1(G953), .A2(G902), .A3(n864), .A4(n749), .ZN(n863) );
  INV_X1 U649 ( .A(G900), .ZN(n749) );
  NAND2_X1 U650 ( .A1(n865), .A2(KEYINPUT13), .ZN(G24) );
  XOR2_X1 U651 ( .A(n818), .B(G122), .Z(n865) );
  NAND4_X1 U652 ( .A1(n866), .A2(n722), .A3(n832), .A4(n834), .ZN(n818) );
  NOR2_X1 U653 ( .A1(n862), .A2(n853), .ZN(n722) );
  NAND3_X1 U654 ( .A1(n867), .A2(n868), .A3(KEYINPUT4), .ZN(G21) );
  OR2_X1 U655 ( .A1(n869), .A2(G119), .ZN(n868) );
  NAND3_X1 U656 ( .A1(KEYINPUT32), .A2(n869), .A3(G119), .ZN(n867) );
  NOR2_X1 U657 ( .A1(n870), .A2(KEYINPUT30), .ZN(n869) );
  INV_X1 U658 ( .A(n817), .ZN(n870) );
  NAND2_X1 U659 ( .A1(n844), .A2(n866), .ZN(n817) );
  AND3_X1 U660 ( .A1(n853), .A2(n862), .A3(n727), .ZN(n844) );
  NAND2_X1 U661 ( .A1(n871), .A2(KEYINPUT12), .ZN(G18) );
  XOR2_X1 U662 ( .A(n816), .B(G116), .Z(n871) );
  NAND3_X1 U663 ( .A1(n737), .A2(n814), .A3(n866), .ZN(n816) );
  NOR2_X1 U664 ( .A1(n832), .A2(n872), .ZN(n814) );
  NAND2_X1 U665 ( .A1(n873), .A2(KEYINPUT11), .ZN(G15) );
  XNOR2_X1 U666 ( .A(n813), .B(G113), .ZN(n873) );
  AND3_X1 U667 ( .A1(n737), .A2(n820), .A3(n866), .ZN(n813) );
  AND3_X1 U668 ( .A1(n830), .A2(n874), .A3(n731), .ZN(n866) );
  NOR2_X1 U669 ( .A1(n729), .A2(n875), .ZN(n731) );
  AND2_X1 U670 ( .A1(G221), .A2(n876), .ZN(n875) );
  INV_X1 U671 ( .A(n802), .ZN(n820) );
  NAND2_X1 U672 ( .A1(n872), .A2(n832), .ZN(n802) );
  INV_X1 U673 ( .A(n834), .ZN(n872) );
  NOR2_X1 U674 ( .A1(n862), .A2(n861), .ZN(n737) );
  NAND3_X1 U675 ( .A1(n877), .A2(n878), .A3(KEYINPUT3), .ZN(G12) );
  OR2_X1 U676 ( .A1(n879), .A2(G110), .ZN(n878) );
  NAND3_X1 U677 ( .A1(KEYINPUT29), .A2(n879), .A3(G110), .ZN(n877) );
  NOR2_X1 U678 ( .A1(n812), .A2(KEYINPUT27), .ZN(n879) );
  AND3_X1 U679 ( .A1(n738), .A2(n815), .A3(n727), .ZN(n812) );
  NOR2_X1 U680 ( .A1(n834), .A2(n832), .ZN(n727) );
  XOR2_X1 U681 ( .A(n880), .B(n778), .Z(n832) );
  INV_X1 U682 ( .A(G475), .ZN(n778) );
  NAND2_X1 U683 ( .A1(n776), .A2(n881), .ZN(n880) );
  XNOR2_X1 U684 ( .A(n882), .B(n883), .ZN(n776) );
  XOR2_X1 U685 ( .A(n884), .B(n885), .Z(n883) );
  XOR2_X1 U686 ( .A(G122), .B(G113), .Z(n885) );
  XOR2_X1 U687 ( .A(G143), .B(G131), .Z(n884) );
  XNOR2_X1 U688 ( .A(n754), .B(n886), .ZN(n882) );
  XNOR2_X1 U689 ( .A(G104), .B(n887), .ZN(n886) );
  NAND2_X1 U690 ( .A1(n888), .A2(G214), .ZN(n887) );
  XOR2_X1 U691 ( .A(n889), .B(n774), .Z(n834) );
  INV_X1 U692 ( .A(G478), .ZN(n774) );
  NAND2_X1 U693 ( .A1(n772), .A2(n881), .ZN(n889) );
  XNOR2_X1 U694 ( .A(n890), .B(n891), .ZN(n772) );
  XOR2_X1 U695 ( .A(G107), .B(n892), .Z(n891) );
  XOR2_X1 U696 ( .A(G122), .B(G116), .Z(n892) );
  XOR2_X1 U697 ( .A(n893), .B(n894), .Z(n890) );
  NOR2_X1 U698 ( .A1(n895), .A2(n769), .ZN(n894) );
  INV_X1 U699 ( .A(G217), .ZN(n769) );
  AND3_X1 U700 ( .A1(n830), .A2(n874), .A3(n829), .ZN(n815) );
  INV_X1 U701 ( .A(n730), .ZN(n829) );
  NAND2_X1 U702 ( .A1(n729), .A2(n896), .ZN(n730) );
  NAND2_X1 U703 ( .A1(G221), .A2(n876), .ZN(n896) );
  XOR2_X1 U704 ( .A(n897), .B(n788), .Z(n729) );
  INV_X1 U705 ( .A(G469), .ZN(n788) );
  NAND2_X1 U706 ( .A1(n786), .A2(n881), .ZN(n897) );
  XNOR2_X1 U707 ( .A(n898), .B(n899), .ZN(n786) );
  XOR2_X1 U708 ( .A(G140), .B(n900), .Z(n899) );
  NOR2_X1 U709 ( .A1(G953), .A2(n748), .ZN(n900) );
  INV_X1 U710 ( .A(G227), .ZN(n748) );
  XOR2_X1 U711 ( .A(n901), .B(n902), .Z(n898) );
  NAND2_X1 U712 ( .A1(n742), .A2(n903), .ZN(n874) );
  NAND4_X1 U713 ( .A1(G953), .A2(G902), .A3(n864), .A4(n760), .ZN(n903) );
  INV_X1 U714 ( .A(G898), .ZN(n760) );
  NAND3_X1 U715 ( .A1(n864), .A2(n743), .A3(G952), .ZN(n742) );
  NAND2_X1 U716 ( .A1(G237), .A2(G234), .ZN(n864) );
  INV_X1 U717 ( .A(n741), .ZN(n830) );
  NAND2_X1 U718 ( .A1(n740), .A2(n904), .ZN(n741) );
  NAND2_X1 U719 ( .A1(G214), .A2(n848), .ZN(n904) );
  INV_X1 U720 ( .A(n905), .ZN(n848) );
  XNOR2_X1 U721 ( .A(n906), .B(n907), .ZN(n740) );
  NOR2_X1 U722 ( .A1(n905), .A2(n792), .ZN(n907) );
  INV_X1 U723 ( .A(G210), .ZN(n792) );
  NOR2_X1 U724 ( .A1(G902), .A2(G237), .ZN(n905) );
  NAND2_X1 U725 ( .A1(n790), .A2(n881), .ZN(n906) );
  XNOR2_X1 U726 ( .A(n908), .B(n909), .ZN(n790) );
  XOR2_X1 U727 ( .A(n910), .B(n911), .Z(n909) );
  NOR2_X1 U728 ( .A1(G953), .A2(n759), .ZN(n910) );
  INV_X1 U729 ( .A(G224), .ZN(n759) );
  XOR2_X1 U730 ( .A(n764), .B(n912), .Z(n908) );
  XOR2_X1 U731 ( .A(n913), .B(n902), .Z(n764) );
  XNOR2_X1 U732 ( .A(n914), .B(n915), .ZN(n902) );
  XOR2_X1 U733 ( .A(G110), .B(G107), .Z(n915) );
  XNOR2_X1 U734 ( .A(G104), .B(G101), .ZN(n914) );
  XNOR2_X1 U735 ( .A(n916), .B(G122), .ZN(n913) );
  AND2_X1 U736 ( .A1(n861), .A2(n862), .ZN(n738) );
  XNOR2_X1 U737 ( .A(n917), .B(n918), .ZN(n862) );
  AND2_X1 U738 ( .A1(n876), .A2(G217), .ZN(n918) );
  NAND2_X1 U739 ( .A1(G234), .A2(n881), .ZN(n876) );
  NAND2_X1 U740 ( .A1(n767), .A2(n881), .ZN(n917) );
  XNOR2_X1 U741 ( .A(n919), .B(n920), .ZN(n767) );
  XOR2_X1 U742 ( .A(G119), .B(n921), .Z(n920) );
  XOR2_X1 U743 ( .A(G137), .B(G128), .Z(n921) );
  XNOR2_X1 U744 ( .A(n922), .B(n923), .ZN(n919) );
  INV_X1 U745 ( .A(n754), .ZN(n923) );
  XOR2_X1 U746 ( .A(G140), .B(n912), .Z(n754) );
  XOR2_X1 U747 ( .A(G125), .B(G146), .Z(n912) );
  XOR2_X1 U748 ( .A(n924), .B(G110), .Z(n922) );
  NAND2_X1 U749 ( .A1(n925), .A2(G221), .ZN(n924) );
  INV_X1 U750 ( .A(n895), .ZN(n925) );
  NAND2_X1 U751 ( .A1(G234), .A2(n743), .ZN(n895) );
  INV_X1 U752 ( .A(G953), .ZN(n743) );
  INV_X1 U753 ( .A(n853), .ZN(n861) );
  XOR2_X1 U754 ( .A(n926), .B(n784), .Z(n853) );
  INV_X1 U755 ( .A(G472), .ZN(n784) );
  NAND2_X1 U756 ( .A1(n782), .A2(n881), .ZN(n926) );
  INV_X1 U757 ( .A(G902), .ZN(n881) );
  XNOR2_X1 U758 ( .A(n927), .B(n928), .ZN(n782) );
  XNOR2_X1 U759 ( .A(G101), .B(n929), .ZN(n928) );
  NAND2_X1 U760 ( .A1(n888), .A2(G210), .ZN(n929) );
  NOR2_X1 U761 ( .A1(G953), .A2(G237), .ZN(n888) );
  XNOR2_X1 U762 ( .A(n901), .B(n930), .ZN(n927) );
  INV_X1 U763 ( .A(n916), .ZN(n930) );
  XOR2_X1 U764 ( .A(G113), .B(n931), .Z(n916) );
  XOR2_X1 U765 ( .A(G119), .B(G116), .Z(n931) );
  XNOR2_X1 U766 ( .A(G146), .B(n755), .ZN(n901) );
  XNOR2_X1 U767 ( .A(n893), .B(n932), .ZN(n755) );
  XOR2_X1 U768 ( .A(G137), .B(G131), .Z(n932) );
  XNOR2_X1 U769 ( .A(G134), .B(n911), .ZN(n893) );
  XOR2_X1 U770 ( .A(G128), .B(G143), .Z(n911) );
endmodule

