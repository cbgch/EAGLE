//Key = 1101101100111001100101111010110000001101110101111000000100011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;

XOR2_X1 U737 ( .A(G107), .B(n1016), .Z(G9) );
NOR4_X1 U738 ( .A1(KEYINPUT33), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1016) );
NOR2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND4_X1 U741 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(G952), .ZN(n1023) );
XOR2_X1 U742 ( .A(n1027), .B(KEYINPUT41), .Z(n1024) );
NAND2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
XOR2_X1 U747 ( .A(KEYINPUT53), .B(n1037), .Z(n1035) );
NAND2_X1 U748 ( .A1(n1038), .A2(n1039), .ZN(n1032) );
NAND4_X1 U749 ( .A1(n1040), .A2(n1038), .A3(n1034), .A4(n1041), .ZN(n1028) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U751 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1042) );
NAND4_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1022) );
NAND3_X1 U754 ( .A1(n1038), .A2(n1053), .A3(n1040), .ZN(n1050) );
INV_X1 U755 ( .A(n1054), .ZN(n1040) );
NAND2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NAND3_X1 U757 ( .A1(n1047), .A2(n1034), .A3(n1057), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1045), .A2(n1058), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1034), .A2(n1061), .ZN(n1060) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1047), .ZN(n1059) );
NAND3_X1 U762 ( .A1(n1034), .A2(n1063), .A3(n1030), .ZN(n1049) );
NOR3_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1054), .ZN(n1030) );
NOR3_X1 U764 ( .A1(n1066), .A2(G953), .A3(n1067), .ZN(n1020) );
INV_X1 U765 ( .A(n1051), .ZN(n1067) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1051) );
NOR4_X1 U767 ( .A1(n1070), .A2(n1036), .A3(n1071), .A4(n1072), .ZN(n1069) );
XOR2_X1 U768 ( .A(n1073), .B(n1074), .Z(n1072) );
XOR2_X1 U769 ( .A(KEYINPUT47), .B(KEYINPUT46), .Z(n1074) );
XOR2_X1 U770 ( .A(n1075), .B(n1076), .Z(n1073) );
NOR2_X1 U771 ( .A1(G472), .A2(KEYINPUT32), .ZN(n1076) );
NOR2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1071) );
NOR2_X1 U773 ( .A1(G902), .A2(n1079), .ZN(n1077) );
NOR4_X1 U774 ( .A1(n1080), .A2(n1081), .A3(n1065), .A4(n1082), .ZN(n1068) );
XNOR2_X1 U775 ( .A(n1083), .B(KEYINPUT6), .ZN(n1080) );
XNOR2_X1 U776 ( .A(G952), .B(KEYINPUT1), .ZN(n1066) );
XOR2_X1 U777 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U778 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U779 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1088) );
NAND3_X1 U781 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1086) );
XOR2_X1 U782 ( .A(n1092), .B(KEYINPUT25), .Z(n1091) );
NAND2_X1 U783 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
XOR2_X1 U785 ( .A(KEYINPUT16), .B(n1093), .Z(n1096) );
XNOR2_X1 U786 ( .A(n1097), .B(n1098), .ZN(n1093) );
XOR2_X1 U787 ( .A(KEYINPUT61), .B(n1094), .Z(n1095) );
NAND2_X1 U788 ( .A1(G953), .A2(n1099), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1026), .A2(G953), .ZN(n1084) );
XOR2_X1 U790 ( .A(n1100), .B(n1101), .Z(G69) );
XOR2_X1 U791 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U793 ( .A1(G953), .A2(n1106), .ZN(n1105) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(n1104) );
XNOR2_X1 U795 ( .A(n1109), .B(n1110), .ZN(n1108) );
NAND2_X1 U796 ( .A1(KEYINPUT29), .A2(n1111), .ZN(n1109) );
XOR2_X1 U797 ( .A(G110), .B(n1112), .Z(n1107) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1102) );
XOR2_X1 U799 ( .A(KEYINPUT60), .B(n1025), .Z(n1114) );
XNOR2_X1 U800 ( .A(G953), .B(KEYINPUT8), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1052), .ZN(n1100) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1106), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XNOR2_X1 U804 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U806 ( .A1(n1117), .A2(n1123), .ZN(G63) );
XOR2_X1 U807 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U808 ( .A1(KEYINPUT18), .A2(n1126), .ZN(n1125) );
NAND2_X1 U809 ( .A1(n1127), .A2(G478), .ZN(n1124) );
NOR2_X1 U810 ( .A1(n1117), .A2(n1128), .ZN(G60) );
XOR2_X1 U811 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U812 ( .A(KEYINPUT37), .B(n1131), .Z(n1130) );
AND2_X1 U813 ( .A1(G475), .A2(n1127), .ZN(n1131) );
XNOR2_X1 U814 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(G57) );
XOR2_X1 U816 ( .A(KEYINPUT27), .B(n1117), .Z(n1134) );
XOR2_X1 U817 ( .A(n1135), .B(n1136), .Z(n1133) );
XOR2_X1 U818 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
AND2_X1 U820 ( .A1(G472), .A2(n1127), .ZN(n1140) );
NOR2_X1 U821 ( .A1(KEYINPUT42), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U822 ( .A(n1142), .B(G128), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1143), .A2(n1144), .ZN(n1137) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1135) );
NAND2_X1 U825 ( .A1(KEYINPUT3), .A2(n1147), .ZN(n1145) );
NOR2_X1 U826 ( .A1(n1117), .A2(n1148), .ZN(G54) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U828 ( .A(n1151), .B(KEYINPUT19), .Z(n1150) );
NAND2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
AND2_X1 U831 ( .A1(n1127), .A2(G469), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1117), .A2(n1154), .ZN(G51) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND3_X1 U834 ( .A1(n1127), .A2(n1157), .A3(KEYINPUT15), .ZN(n1155) );
XNOR2_X1 U835 ( .A(KEYINPUT50), .B(n1078), .ZN(n1157) );
INV_X1 U836 ( .A(n1122), .ZN(n1127) );
NAND2_X1 U837 ( .A1(G902), .A2(n1158), .ZN(n1122) );
NAND2_X1 U838 ( .A1(n1025), .A2(n1026), .ZN(n1158) );
AND4_X1 U839 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1026) );
NOR4_X1 U840 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NOR2_X1 U841 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U842 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1062), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U845 ( .A(KEYINPUT52), .B(n1174), .ZN(n1173) );
NOR3_X1 U846 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1164) );
AND2_X1 U847 ( .A1(n1175), .A2(n1178), .ZN(n1163) );
INV_X1 U848 ( .A(KEYINPUT31), .ZN(n1175) );
INV_X1 U849 ( .A(n1179), .ZN(n1161) );
AND4_X1 U850 ( .A1(n1132), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1025) );
NOR4_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NOR2_X1 U852 ( .A1(KEYINPUT34), .A2(n1187), .ZN(n1186) );
NOR2_X1 U853 ( .A1(n1188), .A2(n1018), .ZN(n1185) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR2_X1 U855 ( .A1(n1064), .A2(n1191), .ZN(n1190) );
NOR2_X1 U856 ( .A1(n1017), .A2(n1019), .ZN(n1189) );
AND3_X1 U857 ( .A1(KEYINPUT24), .A2(n1192), .A3(n1193), .ZN(n1184) );
NOR4_X1 U858 ( .A1(n1063), .A2(n1194), .A3(n1195), .A4(n1065), .ZN(n1183) );
NOR2_X1 U859 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
AND2_X1 U860 ( .A1(n1170), .A2(KEYINPUT34), .ZN(n1197) );
NOR2_X1 U861 ( .A1(KEYINPUT24), .A2(n1198), .ZN(n1196) );
INV_X1 U862 ( .A(n1193), .ZN(n1198) );
NOR2_X1 U863 ( .A1(n1199), .A2(n1200), .ZN(n1181) );
NAND3_X1 U864 ( .A1(n1201), .A2(n1034), .A3(n1057), .ZN(n1132) );
NOR2_X1 U865 ( .A1(n1052), .A2(G952), .ZN(n1117) );
XOR2_X1 U866 ( .A(G146), .B(n1165), .Z(G48) );
AND3_X1 U867 ( .A1(n1057), .A2(n1202), .A3(n1203), .ZN(n1165) );
XOR2_X1 U868 ( .A(G143), .B(n1178), .Z(G45) );
NOR2_X1 U869 ( .A1(n1177), .A2(n1204), .ZN(n1178) );
NAND4_X1 U870 ( .A1(n1205), .A2(n1062), .A3(n1082), .A4(n1083), .ZN(n1177) );
XNOR2_X1 U871 ( .A(n1206), .B(n1207), .ZN(G42) );
NOR3_X1 U872 ( .A1(n1168), .A2(n1174), .A3(n1172), .ZN(n1207) );
XNOR2_X1 U873 ( .A(n1208), .B(n1209), .ZN(G39) );
NOR2_X1 U874 ( .A1(n1210), .A2(n1168), .ZN(n1209) );
XNOR2_X1 U875 ( .A(G134), .B(n1211), .ZN(G36) );
NAND2_X1 U876 ( .A1(KEYINPUT7), .A2(n1179), .ZN(n1211) );
NOR3_X1 U877 ( .A1(n1191), .A2(n1019), .A3(n1168), .ZN(n1179) );
INV_X1 U878 ( .A(n1048), .ZN(n1019) );
XOR2_X1 U879 ( .A(G131), .B(n1212), .Z(G33) );
NOR3_X1 U880 ( .A1(n1168), .A2(n1213), .A3(n1191), .ZN(n1212) );
XNOR2_X1 U881 ( .A(n1057), .B(KEYINPUT9), .ZN(n1213) );
NAND3_X1 U882 ( .A1(n1061), .A2(n1176), .A3(n1038), .ZN(n1168) );
AND2_X1 U883 ( .A1(n1037), .A2(n1214), .ZN(n1038) );
XNOR2_X1 U884 ( .A(G128), .B(n1159), .ZN(G30) );
NAND3_X1 U885 ( .A1(n1048), .A2(n1202), .A3(n1203), .ZN(n1159) );
AND3_X1 U886 ( .A1(n1215), .A2(n1176), .A3(n1205), .ZN(n1203) );
AND2_X1 U887 ( .A1(n1063), .A2(n1061), .ZN(n1205) );
XOR2_X1 U888 ( .A(G101), .B(n1216), .Z(G3) );
NOR4_X1 U889 ( .A1(n1217), .A2(n1218), .A3(n1064), .A4(n1191), .ZN(n1216) );
XNOR2_X1 U890 ( .A(n1063), .B(KEYINPUT62), .ZN(n1217) );
XNOR2_X1 U891 ( .A(G125), .B(n1160), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1057), .A2(n1039), .A3(n1219), .A4(n1047), .ZN(n1160) );
INV_X1 U893 ( .A(n1065), .ZN(n1047) );
NOR2_X1 U894 ( .A1(n1204), .A2(n1220), .ZN(n1219) );
INV_X1 U895 ( .A(n1176), .ZN(n1204) );
NAND2_X1 U896 ( .A1(n1054), .A2(n1221), .ZN(n1176) );
NAND4_X1 U897 ( .A1(n1222), .A2(G953), .A3(n1223), .A4(n1099), .ZN(n1221) );
INV_X1 U898 ( .A(G900), .ZN(n1099) );
XNOR2_X1 U899 ( .A(G902), .B(KEYINPUT40), .ZN(n1222) );
INV_X1 U900 ( .A(n1174), .ZN(n1039) );
INV_X1 U901 ( .A(n1172), .ZN(n1057) );
XNOR2_X1 U902 ( .A(G122), .B(n1180), .ZN(G24) );
NAND4_X1 U903 ( .A1(n1192), .A2(n1034), .A3(n1082), .A4(n1083), .ZN(n1180) );
INV_X1 U904 ( .A(n1017), .ZN(n1034) );
NAND2_X1 U905 ( .A1(n1224), .A2(n1225), .ZN(n1017) );
XNOR2_X1 U906 ( .A(n1226), .B(n1227), .ZN(G21) );
NOR2_X1 U907 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NOR2_X1 U908 ( .A1(KEYINPUT56), .A2(n1230), .ZN(n1229) );
INV_X1 U909 ( .A(n1187), .ZN(n1230) );
NOR2_X1 U910 ( .A1(KEYINPUT4), .A2(n1187), .ZN(n1228) );
NAND2_X1 U911 ( .A1(n1170), .A2(n1192), .ZN(n1187) );
INV_X1 U912 ( .A(n1210), .ZN(n1170) );
NAND3_X1 U913 ( .A1(n1202), .A2(n1215), .A3(n1045), .ZN(n1210) );
XOR2_X1 U914 ( .A(G116), .B(n1200), .Z(G18) );
AND3_X1 U915 ( .A1(n1062), .A2(n1048), .A3(n1192), .ZN(n1200) );
NOR2_X1 U916 ( .A1(n1083), .A2(n1231), .ZN(n1048) );
INV_X1 U917 ( .A(n1082), .ZN(n1231) );
INV_X1 U918 ( .A(n1191), .ZN(n1062) );
XOR2_X1 U919 ( .A(n1232), .B(G113), .Z(G15) );
NAND2_X1 U920 ( .A1(KEYINPUT59), .A2(n1233), .ZN(n1232) );
NAND2_X1 U921 ( .A1(n1193), .A2(n1192), .ZN(n1233) );
NOR3_X1 U922 ( .A1(n1220), .A2(n1194), .A3(n1065), .ZN(n1192) );
NAND2_X1 U923 ( .A1(n1044), .A2(n1234), .ZN(n1065) );
INV_X1 U924 ( .A(n1235), .ZN(n1194) );
NOR2_X1 U925 ( .A1(n1172), .A2(n1191), .ZN(n1193) );
NAND2_X1 U926 ( .A1(n1202), .A2(n1225), .ZN(n1191) );
XOR2_X1 U927 ( .A(n1215), .B(KEYINPUT39), .Z(n1225) );
NAND2_X1 U928 ( .A1(n1236), .A2(n1237), .ZN(n1172) );
XOR2_X1 U929 ( .A(KEYINPUT38), .B(n1083), .Z(n1237) );
XOR2_X1 U930 ( .A(G110), .B(n1199), .Z(G12) );
NOR3_X1 U931 ( .A1(n1174), .A2(n1018), .A3(n1064), .ZN(n1199) );
INV_X1 U932 ( .A(n1045), .ZN(n1064) );
NOR2_X1 U933 ( .A1(n1238), .A2(n1083), .ZN(n1045) );
XNOR2_X1 U934 ( .A(n1239), .B(G475), .ZN(n1083) );
NAND2_X1 U935 ( .A1(n1129), .A2(n1240), .ZN(n1239) );
XNOR2_X1 U936 ( .A(n1241), .B(n1242), .ZN(n1129) );
XOR2_X1 U937 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U938 ( .A(G113), .B(G104), .Z(n1244) );
XOR2_X1 U939 ( .A(KEYINPUT0), .B(G131), .Z(n1243) );
XOR2_X1 U940 ( .A(n1245), .B(n1246), .Z(n1241) );
XOR2_X1 U941 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U942 ( .A1(G122), .A2(KEYINPUT2), .ZN(n1248) );
NOR3_X1 U943 ( .A1(n1249), .A2(G237), .A3(n1250), .ZN(n1247) );
XNOR2_X1 U944 ( .A(G953), .B(KEYINPUT36), .ZN(n1250) );
INV_X1 U945 ( .A(G214), .ZN(n1249) );
XOR2_X1 U946 ( .A(n1251), .B(n1252), .Z(n1245) );
NAND2_X1 U947 ( .A1(KEYINPUT28), .A2(n1206), .ZN(n1251) );
INV_X1 U948 ( .A(G140), .ZN(n1206) );
XNOR2_X1 U949 ( .A(n1236), .B(KEYINPUT57), .ZN(n1238) );
XNOR2_X1 U950 ( .A(n1082), .B(KEYINPUT58), .ZN(n1236) );
XOR2_X1 U951 ( .A(G478), .B(n1253), .Z(n1082) );
NOR2_X1 U952 ( .A1(G902), .A2(n1126), .ZN(n1253) );
NAND3_X1 U953 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1126) );
NAND2_X1 U954 ( .A1(KEYINPUT20), .A2(n1257), .ZN(n1256) );
NAND3_X1 U955 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1255) );
INV_X1 U956 ( .A(KEYINPUT20), .ZN(n1259) );
NAND2_X1 U957 ( .A1(G217), .A2(n1261), .ZN(n1258) );
NAND3_X1 U958 ( .A1(G217), .A2(n1261), .A3(n1262), .ZN(n1254) );
INV_X1 U959 ( .A(n1260), .ZN(n1262) );
NOR2_X1 U960 ( .A1(KEYINPUT63), .A2(n1257), .ZN(n1260) );
XOR2_X1 U961 ( .A(n1263), .B(n1264), .Z(n1257) );
XOR2_X1 U962 ( .A(G122), .B(n1265), .Z(n1264) );
XOR2_X1 U963 ( .A(G143), .B(G128), .Z(n1265) );
XOR2_X1 U964 ( .A(n1266), .B(n1267), .Z(n1263) );
XOR2_X1 U965 ( .A(G116), .B(G107), .Z(n1267) );
NAND2_X1 U966 ( .A1(KEYINPUT26), .A2(n1268), .ZN(n1266) );
INV_X1 U967 ( .A(G134), .ZN(n1268) );
INV_X1 U968 ( .A(n1201), .ZN(n1018) );
NOR2_X1 U969 ( .A1(n1220), .A2(n1218), .ZN(n1201) );
NAND2_X1 U970 ( .A1(n1061), .A2(n1235), .ZN(n1218) );
NAND2_X1 U971 ( .A1(n1054), .A2(n1269), .ZN(n1235) );
NAND4_X1 U972 ( .A1(G902), .A2(G953), .A3(n1223), .A4(n1106), .ZN(n1269) );
INV_X1 U973 ( .A(G898), .ZN(n1106) );
NAND3_X1 U974 ( .A1(n1223), .A2(n1052), .A3(G952), .ZN(n1054) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1223) );
NOR2_X1 U976 ( .A1(n1044), .A2(n1046), .ZN(n1061) );
INV_X1 U977 ( .A(n1234), .ZN(n1046) );
NAND2_X1 U978 ( .A1(G221), .A2(n1270), .ZN(n1234) );
XOR2_X1 U979 ( .A(n1271), .B(G469), .Z(n1044) );
OR2_X1 U980 ( .A1(n1153), .A2(G902), .ZN(n1271) );
XOR2_X1 U981 ( .A(n1272), .B(n1273), .Z(n1153) );
XNOR2_X1 U982 ( .A(n1146), .B(n1274), .ZN(n1273) );
XNOR2_X1 U983 ( .A(n1275), .B(n1276), .ZN(n1274) );
NOR2_X1 U984 ( .A1(KEYINPUT30), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U985 ( .A(n1278), .B(KEYINPUT22), .ZN(n1146) );
XOR2_X1 U986 ( .A(n1279), .B(n1280), .Z(n1272) );
XOR2_X1 U987 ( .A(n1097), .B(n1281), .Z(n1280) );
NAND2_X1 U988 ( .A1(G227), .A2(n1052), .ZN(n1281) );
NAND2_X1 U989 ( .A1(n1282), .A2(n1283), .ZN(n1097) );
NAND2_X1 U990 ( .A1(n1284), .A2(G143), .ZN(n1283) );
XOR2_X1 U991 ( .A(n1285), .B(KEYINPUT44), .Z(n1282) );
OR2_X1 U992 ( .A1(n1284), .A2(G143), .ZN(n1285) );
XOR2_X1 U993 ( .A(n1286), .B(KEYINPUT45), .Z(n1284) );
XNOR2_X1 U994 ( .A(G140), .B(G101), .ZN(n1279) );
INV_X1 U995 ( .A(n1063), .ZN(n1220) );
NOR2_X1 U996 ( .A1(n1036), .A2(n1037), .ZN(n1063) );
NOR2_X1 U997 ( .A1(n1287), .A2(n1070), .ZN(n1037) );
NOR3_X1 U998 ( .A1(n1288), .A2(G902), .A3(n1079), .ZN(n1070) );
INV_X1 U999 ( .A(n1078), .ZN(n1288) );
AND2_X1 U1000 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
OR2_X1 U1001 ( .A1(n1079), .A2(G902), .ZN(n1290) );
XOR2_X1 U1002 ( .A(n1156), .B(KEYINPUT23), .Z(n1079) );
XOR2_X1 U1003 ( .A(n1291), .B(n1292), .Z(n1156) );
XNOR2_X1 U1004 ( .A(n1293), .B(n1252), .ZN(n1292) );
XNOR2_X1 U1005 ( .A(n1294), .B(n1142), .ZN(n1252) );
INV_X1 U1006 ( .A(G125), .ZN(n1294) );
XOR2_X1 U1007 ( .A(n1295), .B(n1296), .Z(n1291) );
NOR2_X1 U1008 ( .A1(G953), .A2(n1116), .ZN(n1296) );
INV_X1 U1009 ( .A(G224), .ZN(n1116) );
XOR2_X1 U1010 ( .A(n1297), .B(n1112), .Z(n1295) );
NOR2_X1 U1011 ( .A1(KEYINPUT13), .A2(G122), .ZN(n1112) );
NAND2_X1 U1012 ( .A1(n1298), .A2(KEYINPUT55), .ZN(n1297) );
XNOR2_X1 U1013 ( .A(n1111), .B(n1110), .ZN(n1298) );
XOR2_X1 U1014 ( .A(G113), .B(n1299), .Z(n1110) );
NOR2_X1 U1015 ( .A1(KEYINPUT49), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U1016 ( .A(G101), .B(n1277), .ZN(n1111) );
XNOR2_X1 U1017 ( .A(G104), .B(G107), .ZN(n1277) );
XNOR2_X1 U1018 ( .A(KEYINPUT14), .B(n1078), .ZN(n1289) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1301), .ZN(n1078) );
INV_X1 U1020 ( .A(n1214), .ZN(n1036) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1301), .ZN(n1214) );
NAND2_X1 U1022 ( .A1(n1302), .A2(n1240), .ZN(n1301) );
NAND2_X1 U1023 ( .A1(n1224), .A2(n1215), .ZN(n1174) );
XOR2_X1 U1024 ( .A(n1081), .B(KEYINPUT51), .Z(n1215) );
XOR2_X1 U1025 ( .A(n1303), .B(n1121), .Z(n1081) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1270), .ZN(n1121) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1240), .ZN(n1270) );
NAND2_X1 U1028 ( .A1(n1119), .A2(n1240), .ZN(n1303) );
XNOR2_X1 U1029 ( .A(n1304), .B(n1305), .ZN(n1119) );
XNOR2_X1 U1030 ( .A(G119), .B(n1306), .ZN(n1305) );
NAND2_X1 U1031 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1032 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1261), .ZN(n1310) );
XOR2_X1 U1034 ( .A(n1311), .B(KEYINPUT5), .Z(n1307) );
NAND3_X1 U1035 ( .A1(G221), .A2(n1261), .A3(n1312), .ZN(n1311) );
INV_X1 U1036 ( .A(n1309), .ZN(n1312) );
XOR2_X1 U1037 ( .A(G137), .B(KEYINPUT43), .Z(n1309) );
AND2_X1 U1038 ( .A1(G234), .A2(n1052), .ZN(n1261) );
XNOR2_X1 U1039 ( .A(n1313), .B(n1293), .ZN(n1304) );
INV_X1 U1040 ( .A(n1275), .ZN(n1293) );
XOR2_X1 U1041 ( .A(G110), .B(G128), .Z(n1275) );
NAND3_X1 U1042 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1313) );
OR2_X1 U1043 ( .A1(n1094), .A2(KEYINPUT11), .ZN(n1316) );
NAND3_X1 U1044 ( .A1(KEYINPUT11), .A2(n1094), .A3(n1286), .ZN(n1315) );
NAND2_X1 U1045 ( .A1(n1317), .A2(n1318), .ZN(n1314) );
NAND2_X1 U1046 ( .A1(KEYINPUT11), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1047 ( .A(KEYINPUT17), .B(n1094), .Z(n1319) );
XOR2_X1 U1048 ( .A(G125), .B(G140), .Z(n1094) );
INV_X1 U1049 ( .A(n1202), .ZN(n1224) );
XNOR2_X1 U1050 ( .A(n1075), .B(G472), .ZN(n1202) );
NAND2_X1 U1051 ( .A1(n1320), .A2(n1240), .ZN(n1075) );
INV_X1 U1052 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1053 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1054 ( .A1(n1143), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1055 ( .A(n1144), .B(KEYINPUT12), .ZN(n1323) );
AND2_X1 U1056 ( .A1(n1324), .A2(G101), .ZN(n1144) );
NOR2_X1 U1057 ( .A1(G101), .A2(n1324), .ZN(n1143) );
AND3_X1 U1058 ( .A1(n1302), .A2(n1052), .A3(G210), .ZN(n1324) );
INV_X1 U1059 ( .A(G953), .ZN(n1052) );
INV_X1 U1060 ( .A(G237), .ZN(n1302) );
NAND2_X1 U1061 ( .A1(KEYINPUT10), .A2(n1325), .ZN(n1321) );
XOR2_X1 U1062 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1063 ( .A(n1098), .B(n1142), .Z(n1327) );
XNOR2_X1 U1064 ( .A(G143), .B(n1286), .ZN(n1142) );
INV_X1 U1065 ( .A(n1317), .ZN(n1286) );
XOR2_X1 U1066 ( .A(G146), .B(KEYINPUT48), .Z(n1317) );
XNOR2_X1 U1067 ( .A(n1278), .B(G128), .ZN(n1098) );
XNOR2_X1 U1068 ( .A(G131), .B(n1328), .ZN(n1278) );
XNOR2_X1 U1069 ( .A(n1208), .B(G134), .ZN(n1328) );
INV_X1 U1070 ( .A(G137), .ZN(n1208) );
XOR2_X1 U1071 ( .A(n1147), .B(n1329), .Z(n1326) );
XNOR2_X1 U1072 ( .A(KEYINPUT22), .B(KEYINPUT54), .ZN(n1329) );
NAND3_X1 U1073 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1147) );
OR2_X1 U1074 ( .A1(n1300), .A2(KEYINPUT21), .ZN(n1332) );
NAND3_X1 U1075 ( .A1(KEYINPUT21), .A2(n1333), .A3(G113), .ZN(n1331) );
OR2_X1 U1076 ( .A1(n1333), .A2(G113), .ZN(n1330) );
NOR2_X1 U1077 ( .A1(KEYINPUT35), .A2(n1334), .ZN(n1333) );
INV_X1 U1078 ( .A(n1300), .ZN(n1334) );
XOR2_X1 U1079 ( .A(G116), .B(n1226), .Z(n1300) );
INV_X1 U1080 ( .A(G119), .ZN(n1226) );
endmodule


