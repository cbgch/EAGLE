//Key = 1001001001010101001010010110101110010101110010001100010110011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300;

XOR2_X1 U716 ( .A(n988), .B(n989), .Z(G9) );
NAND2_X1 U717 ( .A1(KEYINPUT55), .A2(G107), .ZN(n989) );
NOR2_X1 U718 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR3_X1 U719 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NOR2_X1 U720 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U721 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U722 ( .A1(KEYINPUT56), .A2(n999), .ZN(n998) );
NOR4_X1 U723 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
NOR2_X1 U724 ( .A1(n1004), .A2(n1003), .ZN(n997) );
NOR2_X1 U725 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1007), .A2(n1002), .ZN(n1006) );
INV_X1 U727 ( .A(n1008), .ZN(n1002) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
AND3_X1 U730 ( .A1(KEYINPUT56), .A2(n1013), .A3(n1014), .ZN(n1009) );
NOR3_X1 U731 ( .A1(n1012), .A2(n1001), .A3(n1015), .ZN(n1005) );
NAND3_X1 U732 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n992) );
NAND3_X1 U733 ( .A1(n1014), .A2(n1019), .A3(n1020), .ZN(n1018) );
INV_X1 U734 ( .A(n1003), .ZN(n1020) );
NAND2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NAND3_X1 U736 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1008), .A2(n1026), .ZN(n1021) );
NAND2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1023), .ZN(n1028) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1031), .ZN(n1027) );
NAND2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR3_X1 U743 ( .A1(n1036), .A2(G953), .A3(G952), .ZN(n990) );
INV_X1 U744 ( .A(n1016), .ZN(n1036) );
NAND4_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1016) );
NOR4_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
XNOR2_X1 U747 ( .A(n1045), .B(n1046), .ZN(n1044) );
XOR2_X1 U748 ( .A(n1047), .B(n1048), .Z(n1043) );
XNOR2_X1 U749 ( .A(n1049), .B(KEYINPUT10), .ZN(n1048) );
NOR2_X1 U750 ( .A1(n1034), .A2(n1030), .ZN(n1039) );
XNOR2_X1 U751 ( .A(KEYINPUT11), .B(n1029), .ZN(n1038) );
INV_X1 U752 ( .A(n1050), .ZN(n1029) );
XOR2_X1 U753 ( .A(n1051), .B(n1052), .Z(G72) );
NOR2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
AND2_X1 U755 ( .A1(G227), .A2(G900), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1051) );
NAND2_X1 U757 ( .A1(n1057), .A2(n1017), .ZN(n1056) );
XNOR2_X1 U758 ( .A(n1058), .B(n1059), .ZN(n1057) );
NAND3_X1 U759 ( .A1(n1058), .A2(G900), .A3(G953), .ZN(n1055) );
XNOR2_X1 U760 ( .A(n1060), .B(n1061), .ZN(n1058) );
XNOR2_X1 U761 ( .A(n1062), .B(n1063), .ZN(n1061) );
XNOR2_X1 U762 ( .A(n1064), .B(n1065), .ZN(n1060) );
XOR2_X1 U763 ( .A(n1066), .B(n1067), .Z(G69) );
XOR2_X1 U764 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1054), .ZN(n1069) );
XNOR2_X1 U766 ( .A(G953), .B(KEYINPUT14), .ZN(n1054) );
AND2_X1 U767 ( .A1(G224), .A2(G898), .ZN(n1070) );
NAND3_X1 U768 ( .A1(n1071), .A2(n1017), .A3(KEYINPUT59), .ZN(n1068) );
OR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1066) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XOR2_X1 U771 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR2_X1 U772 ( .A1(KEYINPUT24), .A2(n1078), .ZN(n1077) );
NAND3_X1 U773 ( .A1(n1049), .A2(n994), .A3(n1079), .ZN(n1076) );
XNOR2_X1 U774 ( .A(G902), .B(KEYINPUT25), .ZN(n1079) );
NOR2_X1 U775 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XNOR2_X1 U776 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1074), .A2(n1085), .ZN(G60) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND3_X1 U780 ( .A1(G475), .A2(G902), .A3(n1088), .ZN(n1086) );
XOR2_X1 U781 ( .A(n994), .B(KEYINPUT17), .Z(n1088) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(G6) );
NAND2_X1 U783 ( .A1(G104), .A2(n1091), .ZN(n1090) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U785 ( .A(KEYINPUT61), .B(n1094), .Z(n1089) );
NOR3_X1 U786 ( .A1(n1095), .A2(n1032), .A3(n1096), .ZN(n1094) );
XOR2_X1 U787 ( .A(KEYINPUT58), .B(G104), .Z(n1095) );
NOR3_X1 U788 ( .A1(n1074), .A2(n1097), .A3(n1098), .ZN(G57) );
NOR3_X1 U789 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR2_X1 U790 ( .A1(KEYINPUT39), .A2(KEYINPUT51), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1102), .A2(n1103), .ZN(n1097) );
INV_X1 U792 ( .A(n1099), .ZN(n1103) );
XNOR2_X1 U793 ( .A(n1104), .B(n1105), .ZN(n1099) );
XNOR2_X1 U794 ( .A(n1106), .B(n1107), .ZN(n1105) );
NOR2_X1 U795 ( .A1(KEYINPUT19), .A2(n1108), .ZN(n1106) );
XOR2_X1 U796 ( .A(n1109), .B(n1110), .Z(n1104) );
NOR2_X1 U797 ( .A1(n1111), .A2(n1084), .ZN(n1110) );
NAND2_X1 U798 ( .A1(KEYINPUT6), .A2(n1112), .ZN(n1109) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1102) );
INV_X1 U800 ( .A(KEYINPUT39), .ZN(n1114) );
XNOR2_X1 U801 ( .A(n1115), .B(KEYINPUT51), .ZN(n1113) );
NOR2_X1 U802 ( .A1(n1074), .A2(n1116), .ZN(G54) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR3_X1 U804 ( .A1(n1084), .A2(KEYINPUT8), .A3(n1119), .ZN(n1118) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XOR2_X1 U806 ( .A(n1122), .B(KEYINPUT13), .Z(n1121) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U808 ( .A(KEYINPUT49), .B(n1125), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1124), .ZN(n1120) );
XOR2_X1 U810 ( .A(n1126), .B(n1112), .Z(n1125) );
NAND2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U812 ( .A1(n1074), .A2(n1129), .ZN(G51) );
XOR2_X1 U813 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U814 ( .A(n1072), .B(n1132), .ZN(n1131) );
XOR2_X1 U815 ( .A(n1133), .B(n1134), .Z(n1130) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1084), .ZN(n1133) );
NAND2_X1 U817 ( .A1(G902), .A2(n994), .ZN(n1084) );
NAND2_X1 U818 ( .A1(n1059), .A2(n1136), .ZN(n994) );
INV_X1 U819 ( .A(n1071), .ZN(n1136) );
NAND4_X1 U820 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1071) );
AND4_X1 U821 ( .A1(n988), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1140) );
NAND4_X1 U822 ( .A1(n1144), .A2(n1024), .A3(n1014), .A4(n1145), .ZN(n988) );
NAND2_X1 U823 ( .A1(n1093), .A2(n1146), .ZN(n1139) );
XNOR2_X1 U824 ( .A(KEYINPUT45), .B(n1096), .ZN(n1146) );
INV_X1 U825 ( .A(n1092), .ZN(n1096) );
NOR4_X1 U826 ( .A1(n1015), .A2(n1001), .A3(n1000), .A4(n1147), .ZN(n1092) );
INV_X1 U827 ( .A(n1014), .ZN(n1001) );
NAND4_X1 U828 ( .A1(n1008), .A2(n1144), .A3(n1148), .A4(n1145), .ZN(n1138) );
INV_X1 U829 ( .A(n1011), .ZN(n1148) );
NOR2_X1 U830 ( .A1(n1149), .A2(n1150), .ZN(n1011) );
NAND3_X1 U831 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1137) );
XNOR2_X1 U832 ( .A(n1014), .B(KEYINPUT15), .ZN(n1153) );
AND4_X1 U833 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1059) );
AND4_X1 U834 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1162), .A2(n1163), .ZN(n1156) );
AND3_X1 U836 ( .A1(n1164), .A2(n1165), .A3(KEYINPUT29), .ZN(n1163) );
NOR2_X1 U837 ( .A1(n1164), .A2(n1166), .ZN(n1162) );
NOR2_X1 U838 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U839 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1168) );
NOR4_X1 U840 ( .A1(n1000), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1167) );
XNOR2_X1 U841 ( .A(KEYINPUT37), .B(n1032), .ZN(n1172) );
XNOR2_X1 U842 ( .A(KEYINPUT7), .B(n1152), .ZN(n1170) );
NAND2_X1 U843 ( .A1(n1173), .A2(n1093), .ZN(n1155) );
XOR2_X1 U844 ( .A(n1174), .B(KEYINPUT20), .Z(n1173) );
NAND2_X1 U845 ( .A1(n1175), .A2(n1023), .ZN(n1154) );
INV_X1 U846 ( .A(n996), .ZN(n1023) );
XOR2_X1 U847 ( .A(n1176), .B(KEYINPUT41), .Z(n1175) );
NAND4_X1 U848 ( .A1(n1177), .A2(n1150), .A3(n1013), .A4(n1178), .ZN(n1176) );
INV_X1 U849 ( .A(n1000), .ZN(n1013) );
XNOR2_X1 U850 ( .A(n1179), .B(KEYINPUT31), .ZN(n1177) );
XNOR2_X1 U851 ( .A(n1045), .B(KEYINPUT47), .ZN(n1135) );
NOR2_X1 U852 ( .A1(n1017), .A2(G952), .ZN(n1074) );
XNOR2_X1 U853 ( .A(G146), .B(n1161), .ZN(G48) );
NAND3_X1 U854 ( .A1(n1179), .A2(n1178), .A3(n1180), .ZN(n1161) );
XNOR2_X1 U855 ( .A(G143), .B(n1181), .ZN(G45) );
NAND4_X1 U856 ( .A1(n1150), .A2(n1144), .A3(n1152), .A4(n1178), .ZN(n1181) );
XNOR2_X1 U857 ( .A(G140), .B(n1160), .ZN(G42) );
NAND3_X1 U858 ( .A1(n1179), .A2(n1182), .A3(n1149), .ZN(n1160) );
XNOR2_X1 U859 ( .A(G137), .B(n1159), .ZN(G39) );
NAND4_X1 U860 ( .A1(n1183), .A2(n1008), .A3(n1182), .A4(n1041), .ZN(n1159) );
XNOR2_X1 U861 ( .A(G134), .B(n1158), .ZN(G36) );
NAND3_X1 U862 ( .A1(n1150), .A2(n1024), .A3(n1182), .ZN(n1158) );
XNOR2_X1 U863 ( .A(G131), .B(n1184), .ZN(G33) );
NAND2_X1 U864 ( .A1(n1185), .A2(n1182), .ZN(n1184) );
NOR3_X1 U865 ( .A1(n1000), .A2(n1164), .A3(n996), .ZN(n1182) );
NAND2_X1 U866 ( .A1(n1035), .A2(n1186), .ZN(n996) );
INV_X1 U867 ( .A(n1178), .ZN(n1164) );
XNOR2_X1 U868 ( .A(G128), .B(n1187), .ZN(G30) );
NAND2_X1 U869 ( .A1(n1165), .A2(n1178), .ZN(n1187) );
INV_X1 U870 ( .A(n1169), .ZN(n1165) );
NAND2_X1 U871 ( .A1(n1180), .A2(n1024), .ZN(n1169) );
AND3_X1 U872 ( .A1(n1144), .A2(n1041), .A3(n1183), .ZN(n1180) );
XOR2_X1 U873 ( .A(n1188), .B(n1189), .Z(G3) );
NAND2_X1 U874 ( .A1(KEYINPUT44), .A2(G101), .ZN(n1189) );
NAND4_X1 U875 ( .A1(n1008), .A2(n1150), .A3(n1144), .A4(n1190), .ZN(n1188) );
XNOR2_X1 U876 ( .A(KEYINPUT28), .B(n1145), .ZN(n1190) );
XOR2_X1 U877 ( .A(G125), .B(n1191), .Z(G27) );
NOR2_X1 U878 ( .A1(n1032), .A2(n1174), .ZN(n1191) );
NAND4_X1 U879 ( .A1(n1025), .A2(n1149), .A3(n1179), .A4(n1178), .ZN(n1174) );
NAND2_X1 U880 ( .A1(n1003), .A2(n1192), .ZN(n1178) );
NAND4_X1 U881 ( .A1(G953), .A2(G902), .A3(n1193), .A4(n1194), .ZN(n1192) );
INV_X1 U882 ( .A(G900), .ZN(n1194) );
INV_X1 U883 ( .A(n1015), .ZN(n1179) );
XNOR2_X1 U884 ( .A(G122), .B(n1195), .ZN(G24) );
NAND3_X1 U885 ( .A1(n1014), .A2(n1152), .A3(n1151), .ZN(n1195) );
NAND2_X1 U886 ( .A1(n1196), .A2(n1197), .ZN(n1152) );
OR2_X1 U887 ( .A1(n1015), .A2(KEYINPUT60), .ZN(n1197) );
NAND3_X1 U888 ( .A1(n1042), .A2(n1198), .A3(KEYINPUT60), .ZN(n1196) );
NOR2_X1 U889 ( .A1(n1041), .A2(n1183), .ZN(n1014) );
XNOR2_X1 U890 ( .A(G119), .B(n1143), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1151), .A2(n1008), .A3(n1183), .A4(n1041), .ZN(n1143) );
INV_X1 U892 ( .A(n1199), .ZN(n1183) );
XNOR2_X1 U893 ( .A(G116), .B(n1142), .ZN(G18) );
NAND3_X1 U894 ( .A1(n1150), .A2(n1024), .A3(n1151), .ZN(n1142) );
NOR2_X1 U895 ( .A1(n1198), .A2(n1200), .ZN(n1024) );
INV_X1 U896 ( .A(n1171), .ZN(n1150) );
XOR2_X1 U897 ( .A(n1141), .B(n1201), .Z(G15) );
NOR2_X1 U898 ( .A1(G113), .A2(KEYINPUT54), .ZN(n1201) );
NAND2_X1 U899 ( .A1(n1151), .A2(n1185), .ZN(n1141) );
NOR2_X1 U900 ( .A1(n1015), .A2(n1171), .ZN(n1185) );
NAND2_X1 U901 ( .A1(n1199), .A2(n1041), .ZN(n1171) );
NAND2_X1 U902 ( .A1(n1200), .A2(n1198), .ZN(n1015) );
INV_X1 U903 ( .A(n1042), .ZN(n1200) );
NOR3_X1 U904 ( .A1(n1032), .A2(n1147), .A3(n1012), .ZN(n1151) );
INV_X1 U905 ( .A(n1025), .ZN(n1012) );
NOR2_X1 U906 ( .A1(n1050), .A2(n1030), .ZN(n1025) );
INV_X1 U907 ( .A(n1145), .ZN(n1147) );
XNOR2_X1 U908 ( .A(G110), .B(n1202), .ZN(G12) );
NAND4_X1 U909 ( .A1(n1203), .A2(n1008), .A3(n1144), .A4(n1145), .ZN(n1202) );
NAND2_X1 U910 ( .A1(n1003), .A2(n1204), .ZN(n1145) );
NAND3_X1 U911 ( .A1(G902), .A2(n1193), .A3(n1073), .ZN(n1204) );
NOR2_X1 U912 ( .A1(n1017), .A2(G898), .ZN(n1073) );
NAND3_X1 U913 ( .A1(n1193), .A2(n1017), .A3(G952), .ZN(n1003) );
NAND2_X1 U914 ( .A1(G237), .A2(G234), .ZN(n1193) );
NOR2_X1 U915 ( .A1(n1032), .A2(n1000), .ZN(n1144) );
NAND2_X1 U916 ( .A1(n1205), .A2(n1050), .ZN(n1000) );
XOR2_X1 U917 ( .A(n1206), .B(n1119), .Z(n1050) );
INV_X1 U918 ( .A(G469), .ZN(n1119) );
NAND2_X1 U919 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U920 ( .A(n1209), .B(n1210), .Z(n1207) );
XNOR2_X1 U921 ( .A(n1124), .B(n1112), .ZN(n1210) );
XNOR2_X1 U922 ( .A(n1211), .B(n1212), .ZN(n1124) );
XOR2_X1 U923 ( .A(G140), .B(G110), .Z(n1212) );
NAND2_X1 U924 ( .A1(G227), .A2(n1017), .ZN(n1211) );
XOR2_X1 U925 ( .A(n1213), .B(KEYINPUT27), .Z(n1209) );
NAND2_X1 U926 ( .A1(n1214), .A2(n1128), .ZN(n1213) );
NAND2_X1 U927 ( .A1(n1215), .A2(n1216), .ZN(n1128) );
XNOR2_X1 U928 ( .A(n1063), .B(n1217), .ZN(n1216) );
XNOR2_X1 U929 ( .A(G101), .B(n1218), .ZN(n1215) );
XOR2_X1 U930 ( .A(n1127), .B(KEYINPUT36), .Z(n1214) );
NAND2_X1 U931 ( .A1(n1219), .A2(n1220), .ZN(n1127) );
XNOR2_X1 U932 ( .A(n1221), .B(n1218), .ZN(n1220) );
NOR2_X1 U933 ( .A1(KEYINPUT21), .A2(n1222), .ZN(n1218) );
XNOR2_X1 U934 ( .A(G128), .B(n1063), .ZN(n1219) );
NAND2_X1 U935 ( .A1(n1223), .A2(n1224), .ZN(n1063) );
NAND2_X1 U936 ( .A1(KEYINPUT42), .A2(n1225), .ZN(n1224) );
NAND2_X1 U937 ( .A1(KEYINPUT32), .A2(n1226), .ZN(n1223) );
XNOR2_X1 U938 ( .A(n1030), .B(KEYINPUT38), .ZN(n1205) );
AND2_X1 U939 ( .A1(G221), .A2(n1227), .ZN(n1030) );
INV_X1 U940 ( .A(n1093), .ZN(n1032) );
NOR2_X1 U941 ( .A1(n1035), .A2(n1034), .ZN(n1093) );
INV_X1 U942 ( .A(n1186), .ZN(n1034) );
NAND2_X1 U943 ( .A1(G214), .A2(n1228), .ZN(n1186) );
XNOR2_X1 U944 ( .A(n1046), .B(n1229), .ZN(n1035) );
NOR2_X1 U945 ( .A1(n1045), .A2(KEYINPUT1), .ZN(n1229) );
AND2_X1 U946 ( .A1(G210), .A2(n1228), .ZN(n1045) );
NAND2_X1 U947 ( .A1(n1230), .A2(n1208), .ZN(n1228) );
INV_X1 U948 ( .A(G237), .ZN(n1230) );
NAND2_X1 U949 ( .A1(n1231), .A2(n1208), .ZN(n1046) );
XOR2_X1 U950 ( .A(n1232), .B(n1072), .Z(n1231) );
XNOR2_X1 U951 ( .A(n1233), .B(n1234), .ZN(n1072) );
XOR2_X1 U952 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U953 ( .A(n1237), .B(G113), .Z(n1233) );
NAND2_X1 U954 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
OR2_X1 U955 ( .A1(n1222), .A2(n1240), .ZN(n1239) );
XOR2_X1 U956 ( .A(n1241), .B(KEYINPUT16), .Z(n1238) );
NAND2_X1 U957 ( .A1(n1240), .A2(n1222), .ZN(n1241) );
XOR2_X1 U958 ( .A(G107), .B(G104), .Z(n1222) );
XOR2_X1 U959 ( .A(G101), .B(KEYINPUT63), .Z(n1240) );
NAND2_X1 U960 ( .A1(n1242), .A2(n1243), .ZN(n1232) );
NAND2_X1 U961 ( .A1(n1132), .A2(n1244), .ZN(n1243) );
XOR2_X1 U962 ( .A(KEYINPUT3), .B(n1245), .Z(n1242) );
NOR2_X1 U963 ( .A1(n1132), .A2(n1244), .ZN(n1245) );
XOR2_X1 U964 ( .A(KEYINPUT35), .B(n1134), .Z(n1244) );
AND2_X1 U965 ( .A1(G224), .A2(n1017), .ZN(n1134) );
XNOR2_X1 U966 ( .A(G125), .B(n1246), .ZN(n1132) );
NOR2_X1 U967 ( .A1(n1042), .A2(n1198), .ZN(n1008) );
XNOR2_X1 U968 ( .A(n1037), .B(KEYINPUT5), .ZN(n1198) );
XOR2_X1 U969 ( .A(n1247), .B(G475), .Z(n1037) );
NAND2_X1 U970 ( .A1(n1087), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U971 ( .A(KEYINPUT23), .B(n1208), .ZN(n1248) );
XOR2_X1 U972 ( .A(n1249), .B(n1250), .Z(n1087) );
XOR2_X1 U973 ( .A(G104), .B(n1251), .Z(n1250) );
NOR2_X1 U974 ( .A1(KEYINPUT43), .A2(n1252), .ZN(n1251) );
XOR2_X1 U975 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U976 ( .A(n1255), .B(n1256), .Z(n1254) );
NAND2_X1 U977 ( .A1(KEYINPUT30), .A2(n1065), .ZN(n1256) );
NAND2_X1 U978 ( .A1(n1257), .A2(G214), .ZN(n1255) );
XNOR2_X1 U979 ( .A(n1258), .B(n1226), .ZN(n1253) );
XNOR2_X1 U980 ( .A(G122), .B(G113), .ZN(n1249) );
XNOR2_X1 U981 ( .A(n1259), .B(n1260), .ZN(n1042) );
XNOR2_X1 U982 ( .A(KEYINPUT34), .B(n1083), .ZN(n1260) );
INV_X1 U983 ( .A(G478), .ZN(n1083) );
NAND2_X1 U984 ( .A1(n1081), .A2(n1208), .ZN(n1259) );
XNOR2_X1 U985 ( .A(n1261), .B(n1262), .ZN(n1081) );
XOR2_X1 U986 ( .A(n1062), .B(n1236), .Z(n1262) );
XOR2_X1 U987 ( .A(G116), .B(G122), .Z(n1236) );
XNOR2_X1 U988 ( .A(G134), .B(n1217), .ZN(n1062) );
XOR2_X1 U989 ( .A(n1263), .B(n1264), .Z(n1261) );
XNOR2_X1 U990 ( .A(n1265), .B(G107), .ZN(n1264) );
INV_X1 U991 ( .A(G143), .ZN(n1265) );
NAND2_X1 U992 ( .A1(G217), .A2(n1266), .ZN(n1263) );
XNOR2_X1 U993 ( .A(n1149), .B(KEYINPUT26), .ZN(n1203) );
NOR2_X1 U994 ( .A1(n1199), .A2(n1041), .ZN(n1149) );
XOR2_X1 U995 ( .A(n1267), .B(n1111), .Z(n1041) );
INV_X1 U996 ( .A(G472), .ZN(n1111) );
NAND2_X1 U997 ( .A1(n1268), .A2(n1208), .ZN(n1267) );
XOR2_X1 U998 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U999 ( .A(n1101), .B(n1108), .ZN(n1270) );
XNOR2_X1 U1000 ( .A(n1271), .B(n1272), .ZN(n1108) );
NOR2_X1 U1001 ( .A1(KEYINPUT46), .A2(G113), .ZN(n1272) );
XNOR2_X1 U1002 ( .A(G116), .B(G119), .ZN(n1271) );
INV_X1 U1003 ( .A(n1115), .ZN(n1101) );
XOR2_X1 U1004 ( .A(n1273), .B(n1221), .Z(n1115) );
INV_X1 U1005 ( .A(G101), .ZN(n1221) );
NAND2_X1 U1006 ( .A1(n1257), .A2(G210), .ZN(n1273) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1257) );
XOR2_X1 U1008 ( .A(n1274), .B(n1275), .Z(n1269) );
XOR2_X1 U1009 ( .A(KEYINPUT18), .B(KEYINPUT0), .Z(n1275) );
NAND3_X1 U1010 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1274) );
OR2_X1 U1011 ( .A1(n1112), .A2(n1107), .ZN(n1278) );
NAND2_X1 U1012 ( .A1(KEYINPUT12), .A2(n1279), .ZN(n1277) );
NAND2_X1 U1013 ( .A1(n1280), .A2(n1112), .ZN(n1279) );
XNOR2_X1 U1014 ( .A(KEYINPUT48), .B(n1107), .ZN(n1280) );
NAND2_X1 U1015 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
INV_X1 U1016 ( .A(KEYINPUT12), .ZN(n1282) );
NAND2_X1 U1017 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
NAND3_X1 U1018 ( .A1(KEYINPUT48), .A2(n1112), .A3(n1107), .ZN(n1284) );
XOR2_X1 U1019 ( .A(n1285), .B(n1065), .Z(n1112) );
INV_X1 U1020 ( .A(G131), .ZN(n1065) );
NAND2_X1 U1021 ( .A1(n1286), .A2(KEYINPUT62), .ZN(n1285) );
XOR2_X1 U1022 ( .A(n1287), .B(G134), .Z(n1286) );
NAND2_X1 U1023 ( .A1(n1288), .A2(KEYINPUT40), .ZN(n1287) );
XNOR2_X1 U1024 ( .A(G137), .B(KEYINPUT22), .ZN(n1288) );
OR2_X1 U1025 ( .A1(n1107), .A2(KEYINPUT48), .ZN(n1283) );
XNOR2_X1 U1026 ( .A(n1246), .B(KEYINPUT57), .ZN(n1107) );
XNOR2_X1 U1027 ( .A(n1225), .B(n1289), .ZN(n1246) );
NOR2_X1 U1028 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1289) );
INV_X1 U1029 ( .A(n1226), .ZN(n1225) );
XNOR2_X1 U1030 ( .A(G143), .B(n1290), .ZN(n1226) );
XNOR2_X1 U1031 ( .A(n1047), .B(n1291), .ZN(n1199) );
NOR2_X1 U1032 ( .A1(n1049), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1033 ( .A(KEYINPUT4), .B(KEYINPUT33), .Z(n1292) );
AND2_X1 U1034 ( .A1(G217), .A2(n1227), .ZN(n1049) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1208), .ZN(n1227) );
INV_X1 U1036 ( .A(G902), .ZN(n1208) );
OR2_X1 U1037 ( .A1(n1078), .A2(G902), .ZN(n1047) );
XOR2_X1 U1038 ( .A(n1293), .B(n1294), .Z(n1078) );
XOR2_X1 U1039 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1040 ( .A(n1297), .B(n1298), .ZN(n1296) );
NAND2_X1 U1041 ( .A1(KEYINPUT9), .A2(n1217), .ZN(n1298) );
INV_X1 U1042 ( .A(G128), .ZN(n1217) );
NAND2_X1 U1043 ( .A1(KEYINPUT53), .A2(n1290), .ZN(n1297) );
INV_X1 U1044 ( .A(G146), .ZN(n1290) );
XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(KEYINPUT50), .ZN(n1295) );
XOR2_X1 U1046 ( .A(n1064), .B(n1299), .Z(n1293) );
XNOR2_X1 U1047 ( .A(n1300), .B(n1235), .ZN(n1299) );
XOR2_X1 U1048 ( .A(G110), .B(G119), .Z(n1235) );
NAND2_X1 U1049 ( .A1(n1266), .A2(G221), .ZN(n1300) );
AND2_X1 U1050 ( .A1(G234), .A2(n1017), .ZN(n1266) );
INV_X1 U1051 ( .A(G953), .ZN(n1017) );
XNOR2_X1 U1052 ( .A(G137), .B(n1258), .ZN(n1064) );
XOR2_X1 U1053 ( .A(G125), .B(G140), .Z(n1258) );
endmodule


