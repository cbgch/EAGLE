//Key = 1110010011101100000101011101000010111101100001001101100010100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U769 ( .A(n1058), .B(n1059), .Z(G9) );
NAND2_X1 U770 ( .A1(KEYINPUT2), .A2(G107), .ZN(n1059) );
NOR2_X1 U771 ( .A1(n1060), .A2(n1061), .ZN(G75) );
NOR4_X1 U772 ( .A1(n1062), .A2(n1063), .A3(KEYINPUT44), .A4(G953), .ZN(n1061) );
NAND3_X1 U773 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NAND2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND4_X1 U776 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NAND2_X1 U777 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U778 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U779 ( .A1(n1079), .A2(n1080), .A3(n1078), .ZN(n1069) );
NAND2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1072), .A2(n1083), .ZN(n1082) );
NAND2_X1 U782 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U784 ( .A(n1071), .B(KEYINPUT25), .ZN(n1086) );
NAND2_X1 U785 ( .A1(n1071), .A2(n1088), .ZN(n1084) );
NAND2_X1 U786 ( .A1(n1073), .A2(n1089), .ZN(n1081) );
NAND2_X1 U787 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U788 ( .A1(n1072), .A2(n1092), .ZN(n1091) );
NAND2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U790 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U791 ( .A1(n1071), .A2(n1097), .ZN(n1090) );
INV_X1 U792 ( .A(n1098), .ZN(n1067) );
NOR3_X1 U793 ( .A1(n1063), .A2(G953), .A3(G952), .ZN(n1060) );
AND4_X1 U794 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1063) );
NOR4_X1 U795 ( .A1(n1095), .A2(n1103), .A3(n1077), .A4(n1104), .ZN(n1102) );
AND2_X1 U796 ( .A1(n1105), .A2(G469), .ZN(n1104) );
AND2_X1 U797 ( .A1(n1072), .A2(n1106), .ZN(n1101) );
XOR2_X1 U798 ( .A(n1107), .B(KEYINPUT4), .Z(n1099) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U801 ( .A(n1112), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
NAND2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U805 ( .A(n1064), .B(n1119), .ZN(n1117) );
NAND3_X1 U806 ( .A1(n1119), .A2(G900), .A3(G953), .ZN(n1115) );
XNOR2_X1 U807 ( .A(n1120), .B(n1121), .ZN(n1119) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U809 ( .A(G131), .B(n1124), .ZN(n1120) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U812 ( .A(KEYINPUT46), .B(n1129), .Z(n1128) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U814 ( .A(n1132), .B(KEYINPUT49), .Z(n1130) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1132), .ZN(n1127) );
NAND2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1118), .B(KEYINPUT16), .Z(n1134) );
INV_X1 U818 ( .A(n1131), .ZN(n1133) );
NAND2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
NAND2_X1 U820 ( .A1(G953), .A2(n1138), .ZN(n1137) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(n1136) );
NOR2_X1 U822 ( .A1(KEYINPUT31), .A2(n1141), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1112), .A2(n1142), .ZN(n1125) );
NAND2_X1 U824 ( .A1(G898), .A2(G224), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1118), .B(KEYINPUT27), .Z(n1112) );
NOR3_X1 U826 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(G66) );
NOR3_X1 U827 ( .A1(n1146), .A2(G953), .A3(G952), .ZN(n1145) );
AND2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
INV_X1 U829 ( .A(KEYINPUT7), .ZN(n1146) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1143) );
NAND2_X1 U831 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1147), .A2(n1152), .ZN(G63) );
XOR2_X1 U833 ( .A(n1153), .B(n1154), .Z(n1152) );
AND2_X1 U834 ( .A1(G478), .A2(n1150), .ZN(n1154) );
NAND2_X1 U835 ( .A1(KEYINPUT5), .A2(n1155), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1147), .A2(n1156), .ZN(G60) );
XOR2_X1 U837 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U838 ( .A1(n1150), .A2(G475), .ZN(n1157) );
XOR2_X1 U839 ( .A(n1159), .B(n1160), .Z(G6) );
NAND2_X1 U840 ( .A1(KEYINPUT34), .A2(G104), .ZN(n1160) );
NOR2_X1 U841 ( .A1(n1147), .A2(n1161), .ZN(G57) );
XOR2_X1 U842 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U843 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U844 ( .A(n1166), .B(n1167), .Z(n1162) );
XOR2_X1 U845 ( .A(n1168), .B(G101), .Z(n1167) );
NAND2_X1 U846 ( .A1(n1150), .A2(G472), .ZN(n1168) );
NAND2_X1 U847 ( .A1(KEYINPUT1), .A2(n1169), .ZN(n1166) );
NOR2_X1 U848 ( .A1(n1147), .A2(n1170), .ZN(G54) );
XOR2_X1 U849 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U850 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U851 ( .A1(KEYINPUT29), .A2(n1175), .ZN(n1174) );
XOR2_X1 U852 ( .A(n1176), .B(n1177), .Z(n1171) );
NOR2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U854 ( .A(KEYINPUT55), .B(n1180), .Z(n1179) );
AND2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U856 ( .A1(n1182), .A2(n1181), .ZN(n1178) );
NAND2_X1 U857 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NAND2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U859 ( .A(G140), .ZN(n1186) );
XNOR2_X1 U860 ( .A(G110), .B(KEYINPUT17), .ZN(n1185) );
NAND2_X1 U861 ( .A1(G140), .A2(n1187), .ZN(n1183) );
XNOR2_X1 U862 ( .A(G110), .B(KEYINPUT13), .ZN(n1187) );
NOR2_X1 U863 ( .A1(n1113), .A2(G953), .ZN(n1182) );
NAND2_X1 U864 ( .A1(n1150), .A2(G469), .ZN(n1176) );
NOR2_X1 U865 ( .A1(n1147), .A2(n1188), .ZN(G51) );
XOR2_X1 U866 ( .A(n1189), .B(n1190), .Z(n1188) );
NAND2_X1 U867 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U868 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U869 ( .A(n1195), .B(KEYINPUT38), .Z(n1191) );
OR2_X1 U870 ( .A1(n1194), .A2(n1193), .ZN(n1195) );
XNOR2_X1 U871 ( .A(n1196), .B(n1197), .ZN(n1194) );
XOR2_X1 U872 ( .A(G125), .B(n1198), .Z(n1197) );
NAND2_X1 U873 ( .A1(KEYINPUT23), .A2(n1164), .ZN(n1196) );
NAND2_X1 U874 ( .A1(n1150), .A2(n1199), .ZN(n1189) );
AND2_X1 U875 ( .A1(G902), .A2(n1200), .ZN(n1150) );
NAND2_X1 U876 ( .A1(n1066), .A2(n1064), .ZN(n1200) );
AND4_X1 U877 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1064) );
AND4_X1 U878 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NOR2_X1 U879 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NOR2_X1 U880 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND4_X1 U881 ( .A1(n1213), .A2(n1071), .A3(n1214), .A4(n1075), .ZN(n1212) );
INV_X1 U882 ( .A(KEYINPUT22), .ZN(n1211) );
NOR2_X1 U883 ( .A1(KEYINPUT22), .A2(n1215), .ZN(n1209) );
NAND2_X1 U884 ( .A1(n1216), .A2(n1217), .ZN(n1202) );
XNOR2_X1 U885 ( .A(n1218), .B(KEYINPUT36), .ZN(n1216) );
NAND2_X1 U886 ( .A1(n1219), .A2(n1220), .ZN(n1201) );
NAND2_X1 U887 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XOR2_X1 U888 ( .A(KEYINPUT21), .B(n1223), .Z(n1221) );
INV_X1 U889 ( .A(n1224), .ZN(n1219) );
INV_X1 U890 ( .A(n1135), .ZN(n1066) );
NAND4_X1 U891 ( .A1(n1225), .A2(n1159), .A3(n1226), .A4(n1227), .ZN(n1135) );
AND4_X1 U892 ( .A1(n1228), .A2(n1229), .A3(n1058), .A4(n1230), .ZN(n1227) );
NAND4_X1 U893 ( .A1(n1231), .A2(n1088), .A3(n1072), .A4(n1232), .ZN(n1058) );
NAND2_X1 U894 ( .A1(n1233), .A2(n1097), .ZN(n1226) );
NAND2_X1 U895 ( .A1(n1222), .A2(n1234), .ZN(n1097) );
NAND4_X1 U896 ( .A1(n1087), .A2(n1231), .A3(n1072), .A4(n1232), .ZN(n1159) );
NAND3_X1 U897 ( .A1(n1088), .A2(n1235), .A3(n1236), .ZN(n1225) );
XOR2_X1 U898 ( .A(KEYINPUT26), .B(n1223), .Z(n1235) );
NOR2_X1 U899 ( .A1(n1118), .A2(G952), .ZN(n1147) );
XOR2_X1 U900 ( .A(n1237), .B(n1238), .Z(G48) );
NAND2_X1 U901 ( .A1(n1218), .A2(n1217), .ZN(n1238) );
AND3_X1 U902 ( .A1(n1087), .A2(n1239), .A3(n1240), .ZN(n1218) );
XNOR2_X1 U903 ( .A(G143), .B(n1208), .ZN(G45) );
NAND3_X1 U904 ( .A1(n1241), .A2(n1223), .A3(n1242), .ZN(n1208) );
NOR3_X1 U905 ( .A1(n1093), .A2(n1106), .A3(n1100), .ZN(n1242) );
XOR2_X1 U906 ( .A(G140), .B(n1243), .Z(G42) );
NOR2_X1 U907 ( .A1(n1222), .A2(n1224), .ZN(n1243) );
NAND2_X1 U908 ( .A1(n1244), .A2(n1245), .ZN(G39) );
NAND2_X1 U909 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U910 ( .A(KEYINPUT3), .B(n1207), .ZN(n1246) );
NAND2_X1 U911 ( .A1(G137), .A2(n1248), .ZN(n1244) );
XOR2_X1 U912 ( .A(n1207), .B(KEYINPUT59), .Z(n1248) );
NAND4_X1 U913 ( .A1(n1071), .A2(n1240), .A3(n1239), .A4(n1073), .ZN(n1207) );
XNOR2_X1 U914 ( .A(G134), .B(n1215), .ZN(G36) );
NAND3_X1 U915 ( .A1(n1241), .A2(n1071), .A3(n1213), .ZN(n1215) );
XOR2_X1 U916 ( .A(G131), .B(n1249), .Z(G33) );
NOR2_X1 U917 ( .A1(n1234), .A2(n1224), .ZN(n1249) );
NAND3_X1 U918 ( .A1(n1071), .A2(n1087), .A3(n1241), .ZN(n1224) );
NOR2_X1 U919 ( .A1(n1075), .A2(n1250), .ZN(n1241) );
AND2_X1 U920 ( .A1(n1251), .A2(n1096), .ZN(n1071) );
XNOR2_X1 U921 ( .A(n1095), .B(KEYINPUT53), .ZN(n1251) );
INV_X1 U922 ( .A(n1223), .ZN(n1234) );
XNOR2_X1 U923 ( .A(G128), .B(n1206), .ZN(G30) );
NAND4_X1 U924 ( .A1(n1240), .A2(n1088), .A3(n1217), .A4(n1232), .ZN(n1206) );
AND3_X1 U925 ( .A1(n1252), .A2(n1214), .A3(n1253), .ZN(n1240) );
XOR2_X1 U926 ( .A(n1254), .B(G101), .Z(G3) );
NAND2_X1 U927 ( .A1(KEYINPUT61), .A2(n1255), .ZN(n1254) );
NAND2_X1 U928 ( .A1(n1233), .A2(n1223), .ZN(n1255) );
AND3_X1 U929 ( .A1(n1073), .A2(n1232), .A3(n1231), .ZN(n1233) );
XOR2_X1 U930 ( .A(n1256), .B(n1205), .Z(G27) );
NAND4_X1 U931 ( .A1(n1087), .A2(n1078), .A3(n1257), .A4(n1258), .ZN(n1205) );
NOR3_X1 U932 ( .A1(n1093), .A2(n1077), .A3(n1250), .ZN(n1258) );
INV_X1 U933 ( .A(n1214), .ZN(n1250) );
NAND2_X1 U934 ( .A1(n1098), .A2(n1259), .ZN(n1214) );
NAND4_X1 U935 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1114), .ZN(n1259) );
INV_X1 U936 ( .A(G900), .ZN(n1114) );
INV_X1 U937 ( .A(n1080), .ZN(n1077) );
INV_X1 U938 ( .A(n1217), .ZN(n1093) );
XOR2_X1 U939 ( .A(n1261), .B(n1230), .Z(G24) );
NAND4_X1 U940 ( .A1(n1236), .A2(n1072), .A3(n1262), .A4(n1263), .ZN(n1230) );
INV_X1 U941 ( .A(n1100), .ZN(n1262) );
NOR2_X1 U942 ( .A1(n1252), .A2(n1253), .ZN(n1072) );
XOR2_X1 U943 ( .A(n1264), .B(n1229), .Z(G21) );
NAND4_X1 U944 ( .A1(n1236), .A2(n1073), .A3(n1253), .A4(n1252), .ZN(n1229) );
INV_X1 U945 ( .A(n1265), .ZN(n1252) );
XNOR2_X1 U946 ( .A(G116), .B(n1266), .ZN(G18) );
NAND2_X1 U947 ( .A1(n1213), .A2(n1236), .ZN(n1266) );
AND2_X1 U948 ( .A1(n1223), .A2(n1088), .ZN(n1213) );
XNOR2_X1 U949 ( .A(G113), .B(n1267), .ZN(G15) );
NAND2_X1 U950 ( .A1(KEYINPUT58), .A2(n1268), .ZN(n1267) );
INV_X1 U951 ( .A(n1228), .ZN(n1268) );
NAND3_X1 U952 ( .A1(n1223), .A2(n1087), .A3(n1236), .ZN(n1228) );
AND3_X1 U953 ( .A1(n1078), .A2(n1080), .A3(n1231), .ZN(n1236) );
AND2_X1 U954 ( .A1(n1269), .A2(n1263), .ZN(n1087) );
XOR2_X1 U955 ( .A(n1270), .B(n1100), .Z(n1269) );
NOR2_X1 U956 ( .A1(n1253), .A2(n1265), .ZN(n1223) );
XNOR2_X1 U957 ( .A(G110), .B(n1271), .ZN(G12) );
NAND4_X1 U958 ( .A1(n1257), .A2(n1231), .A3(n1272), .A4(n1073), .ZN(n1271) );
NAND2_X1 U959 ( .A1(n1273), .A2(n1274), .ZN(n1073) );
NAND2_X1 U960 ( .A1(n1088), .A2(n1270), .ZN(n1274) );
INV_X1 U961 ( .A(KEYINPUT24), .ZN(n1270) );
NOR2_X1 U962 ( .A1(n1263), .A2(n1100), .ZN(n1088) );
INV_X1 U963 ( .A(n1106), .ZN(n1263) );
NAND3_X1 U964 ( .A1(n1106), .A2(n1100), .A3(KEYINPUT24), .ZN(n1273) );
XOR2_X1 U965 ( .A(n1275), .B(G478), .Z(n1100) );
NAND2_X1 U966 ( .A1(n1155), .A2(n1276), .ZN(n1275) );
XOR2_X1 U967 ( .A(n1277), .B(n1278), .Z(n1155) );
NOR3_X1 U968 ( .A1(n1279), .A2(KEYINPUT11), .A3(n1280), .ZN(n1278) );
NOR2_X1 U969 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U970 ( .A(KEYINPUT63), .B(n1283), .Z(n1279) );
AND2_X1 U971 ( .A1(n1282), .A2(n1281), .ZN(n1283) );
XNOR2_X1 U972 ( .A(n1284), .B(n1285), .ZN(n1281) );
NOR2_X1 U973 ( .A1(KEYINPUT6), .A2(n1261), .ZN(n1285) );
INV_X1 U974 ( .A(G122), .ZN(n1261) );
XNOR2_X1 U975 ( .A(G107), .B(G116), .ZN(n1284) );
XNOR2_X1 U976 ( .A(n1286), .B(n1287), .ZN(n1282) );
XOR2_X1 U977 ( .A(KEYINPUT8), .B(G134), .Z(n1287) );
NAND2_X1 U978 ( .A1(KEYINPUT12), .A2(n1288), .ZN(n1286) );
NAND2_X1 U979 ( .A1(G217), .A2(n1289), .ZN(n1277) );
XOR2_X1 U980 ( .A(n1290), .B(G475), .Z(n1106) );
NAND2_X1 U981 ( .A1(n1158), .A2(n1276), .ZN(n1290) );
XNOR2_X1 U982 ( .A(n1291), .B(n1292), .ZN(n1158) );
XOR2_X1 U983 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U984 ( .A(G122), .B(G113), .Z(n1294) );
XOR2_X1 U985 ( .A(G143), .B(G131), .Z(n1293) );
XOR2_X1 U986 ( .A(n1295), .B(n1296), .Z(n1291) );
AND2_X1 U987 ( .A1(G214), .A2(n1297), .ZN(n1296) );
XOR2_X1 U988 ( .A(n1298), .B(G104), .Z(n1295) );
NAND3_X1 U989 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1298) );
NAND2_X1 U990 ( .A1(KEYINPUT62), .A2(G146), .ZN(n1301) );
OR3_X1 U991 ( .A1(G146), .A2(KEYINPUT62), .A3(n1122), .ZN(n1300) );
NAND2_X1 U992 ( .A1(n1122), .A2(n1302), .ZN(n1299) );
NAND2_X1 U993 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U994 ( .A(KEYINPUT62), .ZN(n1304) );
XOR2_X1 U995 ( .A(n1237), .B(KEYINPUT50), .Z(n1303) );
XOR2_X1 U996 ( .A(KEYINPUT18), .B(n1232), .Z(n1272) );
XOR2_X1 U997 ( .A(n1239), .B(KEYINPUT43), .Z(n1232) );
INV_X1 U998 ( .A(n1075), .ZN(n1239) );
NAND2_X1 U999 ( .A1(n1305), .A2(n1080), .ZN(n1075) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1306), .ZN(n1080) );
XOR2_X1 U1001 ( .A(KEYINPUT40), .B(n1078), .Z(n1305) );
NOR2_X1 U1002 ( .A1(n1307), .A2(n1103), .ZN(n1078) );
NOR2_X1 U1003 ( .A1(n1105), .A2(G469), .ZN(n1103) );
AND2_X1 U1004 ( .A1(n1308), .A2(n1105), .ZN(n1307) );
NAND2_X1 U1005 ( .A1(n1309), .A2(n1276), .ZN(n1105) );
XOR2_X1 U1006 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1007 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1008 ( .A(G140), .B(G110), .Z(n1313) );
NOR2_X1 U1009 ( .A1(KEYINPUT47), .A2(n1173), .ZN(n1312) );
AND2_X1 U1010 ( .A1(n1314), .A2(n1315), .ZN(n1173) );
NAND2_X1 U1011 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1012 ( .A(n1318), .B(n1319), .Z(n1316) );
NAND2_X1 U1013 ( .A1(n1123), .A2(n1320), .ZN(n1314) );
XOR2_X1 U1014 ( .A(n1319), .B(G101), .Z(n1320) );
NAND2_X1 U1015 ( .A1(KEYINPUT39), .A2(n1321), .ZN(n1319) );
INV_X1 U1016 ( .A(n1317), .ZN(n1123) );
NAND2_X1 U1017 ( .A1(n1322), .A2(n1323), .ZN(n1317) );
NAND3_X1 U1018 ( .A1(G128), .A2(n1324), .A3(n1325), .ZN(n1323) );
INV_X1 U1019 ( .A(KEYINPUT48), .ZN(n1325) );
XOR2_X1 U1020 ( .A(G146), .B(G143), .Z(n1324) );
NAND2_X1 U1021 ( .A1(n1326), .A2(KEYINPUT48), .ZN(n1322) );
XOR2_X1 U1022 ( .A(n1175), .B(n1327), .Z(n1310) );
NOR2_X1 U1023 ( .A1(KEYINPUT54), .A2(n1113), .ZN(n1327) );
INV_X1 U1024 ( .A(G227), .ZN(n1113) );
XOR2_X1 U1025 ( .A(KEYINPUT15), .B(G469), .Z(n1308) );
AND2_X1 U1026 ( .A1(n1217), .A2(n1328), .ZN(n1231) );
NAND2_X1 U1027 ( .A1(n1098), .A2(n1329), .ZN(n1328) );
NAND4_X1 U1028 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1138), .ZN(n1329) );
INV_X1 U1029 ( .A(G898), .ZN(n1138) );
NAND3_X1 U1030 ( .A1(n1260), .A2(n1118), .A3(n1330), .ZN(n1098) );
XNOR2_X1 U1031 ( .A(G952), .B(KEYINPUT45), .ZN(n1330) );
NAND2_X1 U1032 ( .A1(G237), .A2(n1331), .ZN(n1260) );
XOR2_X1 U1033 ( .A(KEYINPUT42), .B(G234), .Z(n1331) );
NOR2_X1 U1034 ( .A1(n1096), .A2(n1332), .ZN(n1217) );
XNOR2_X1 U1035 ( .A(KEYINPUT19), .B(n1095), .ZN(n1332) );
AND2_X1 U1036 ( .A1(G214), .A2(n1333), .ZN(n1095) );
XNOR2_X1 U1037 ( .A(n1107), .B(KEYINPUT56), .ZN(n1096) );
XOR2_X1 U1038 ( .A(n1334), .B(n1199), .Z(n1107) );
AND2_X1 U1039 ( .A1(G210), .A2(n1333), .ZN(n1199) );
NAND2_X1 U1040 ( .A1(n1276), .A2(n1335), .ZN(n1333) );
INV_X1 U1041 ( .A(G237), .ZN(n1335) );
NAND2_X1 U1042 ( .A1(n1336), .A2(n1276), .ZN(n1334) );
XOR2_X1 U1043 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1044 ( .A(G125), .B(n1339), .Z(n1338) );
NOR2_X1 U1045 ( .A1(KEYINPUT41), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1046 ( .A(KEYINPUT52), .B(n1198), .Z(n1340) );
AND2_X1 U1047 ( .A1(G224), .A2(n1118), .ZN(n1198) );
XOR2_X1 U1048 ( .A(n1193), .B(n1326), .Z(n1337) );
INV_X1 U1049 ( .A(n1164), .ZN(n1326) );
XOR2_X1 U1050 ( .A(n1140), .B(n1141), .Z(n1193) );
XOR2_X1 U1051 ( .A(n1341), .B(n1342), .Z(n1141) );
XOR2_X1 U1052 ( .A(n1343), .B(KEYINPUT32), .Z(n1341) );
NAND2_X1 U1053 ( .A1(KEYINPUT9), .A2(G113), .ZN(n1343) );
XNOR2_X1 U1054 ( .A(n1344), .B(n1345), .ZN(n1140) );
XOR2_X1 U1055 ( .A(G110), .B(n1346), .Z(n1345) );
XOR2_X1 U1056 ( .A(KEYINPUT60), .B(G122), .Z(n1346) );
XOR2_X1 U1057 ( .A(n1318), .B(n1321), .Z(n1344) );
XOR2_X1 U1058 ( .A(G104), .B(G107), .Z(n1321) );
INV_X1 U1059 ( .A(G101), .ZN(n1318) );
INV_X1 U1060 ( .A(n1222), .ZN(n1257) );
NAND2_X1 U1061 ( .A1(n1265), .A2(n1253), .ZN(n1222) );
XNOR2_X1 U1062 ( .A(n1347), .B(n1151), .ZN(n1253) );
AND2_X1 U1063 ( .A1(G217), .A2(n1306), .ZN(n1151) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1276), .ZN(n1306) );
NAND2_X1 U1065 ( .A1(n1276), .A2(n1148), .ZN(n1347) );
NAND2_X1 U1066 ( .A1(n1348), .A2(n1349), .ZN(n1148) );
NAND2_X1 U1067 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
XOR2_X1 U1068 ( .A(KEYINPUT0), .B(n1352), .Z(n1348) );
NOR2_X1 U1069 ( .A1(n1350), .A2(n1351), .ZN(n1352) );
XOR2_X1 U1070 ( .A(n1353), .B(G137), .Z(n1351) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1289), .ZN(n1353) );
AND2_X1 U1072 ( .A1(G234), .A2(n1118), .ZN(n1289) );
INV_X1 U1073 ( .A(G953), .ZN(n1118) );
XOR2_X1 U1074 ( .A(n1354), .B(n1355), .Z(n1350) );
NOR2_X1 U1075 ( .A1(KEYINPUT30), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1076 ( .A(n1237), .B(n1122), .Z(n1356) );
XNOR2_X1 U1077 ( .A(n1256), .B(G140), .ZN(n1122) );
INV_X1 U1078 ( .A(G125), .ZN(n1256) );
XOR2_X1 U1079 ( .A(n1357), .B(G110), .Z(n1354) );
NAND3_X1 U1080 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1357) );
OR2_X1 U1081 ( .A1(n1264), .A2(G128), .ZN(n1360) );
NAND2_X1 U1082 ( .A1(KEYINPUT57), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1083 ( .A1(G128), .A2(n1362), .ZN(n1361) );
XOR2_X1 U1084 ( .A(KEYINPUT37), .B(G119), .Z(n1362) );
NAND2_X1 U1085 ( .A1(n1363), .A2(n1364), .ZN(n1358) );
INV_X1 U1086 ( .A(KEYINPUT57), .ZN(n1364) );
NAND2_X1 U1087 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
OR2_X1 U1088 ( .A1(n1264), .A2(KEYINPUT37), .ZN(n1366) );
NAND3_X1 U1089 ( .A1(G128), .A2(n1264), .A3(KEYINPUT37), .ZN(n1365) );
INV_X1 U1090 ( .A(G119), .ZN(n1264) );
INV_X1 U1091 ( .A(G902), .ZN(n1276) );
XNOR2_X1 U1092 ( .A(G472), .B(n1367), .ZN(n1265) );
NOR2_X1 U1093 ( .A1(G902), .A2(n1368), .ZN(n1367) );
NOR2_X1 U1094 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
XOR2_X1 U1095 ( .A(n1371), .B(KEYINPUT35), .Z(n1370) );
NAND2_X1 U1096 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
XNOR2_X1 U1097 ( .A(n1374), .B(KEYINPUT51), .ZN(n1372) );
NOR2_X1 U1098 ( .A1(n1374), .A2(n1373), .ZN(n1369) );
XOR2_X1 U1099 ( .A(G101), .B(n1375), .Z(n1373) );
NOR2_X1 U1100 ( .A1(KEYINPUT20), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1101 ( .A(n1169), .B(KEYINPUT14), .Z(n1376) );
NAND2_X1 U1102 ( .A1(n1297), .A2(G210), .ZN(n1169) );
NOR2_X1 U1103 ( .A1(G953), .A2(G237), .ZN(n1297) );
XNOR2_X1 U1104 ( .A(n1165), .B(n1377), .ZN(n1374) );
NOR2_X1 U1105 ( .A1(KEYINPUT33), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1106 ( .A(n1164), .B(KEYINPUT10), .Z(n1378) );
XOR2_X1 U1107 ( .A(n1237), .B(n1288), .Z(n1164) );
XOR2_X1 U1108 ( .A(G143), .B(G128), .Z(n1288) );
INV_X1 U1109 ( .A(G146), .ZN(n1237) );
XOR2_X1 U1110 ( .A(n1379), .B(n1342), .Z(n1165) );
XOR2_X1 U1111 ( .A(G116), .B(G119), .Z(n1342) );
XOR2_X1 U1112 ( .A(n1175), .B(G113), .Z(n1379) );
XNOR2_X1 U1113 ( .A(G131), .B(n1380), .ZN(n1175) );
NOR2_X1 U1114 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
AND3_X1 U1115 ( .A1(KEYINPUT28), .A2(n1247), .A3(G134), .ZN(n1382) );
INV_X1 U1116 ( .A(G137), .ZN(n1247) );
NOR2_X1 U1117 ( .A1(KEYINPUT28), .A2(n1124), .ZN(n1381) );
XOR2_X1 U1118 ( .A(G134), .B(G137), .Z(n1124) );
endmodule


