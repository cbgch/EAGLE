//Key = 0101101100111000101001000101110001001011010111111111000100100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316;

XNOR2_X1 U722 ( .A(G107), .B(n995), .ZN(G9) );
NOR2_X1 U723 ( .A1(n996), .A2(n997), .ZN(G75) );
XOR2_X1 U724 ( .A(KEYINPUT0), .B(n998), .Z(n997) );
NOR3_X1 U725 ( .A1(n999), .A2(G953), .A3(G952), .ZN(n998) );
NOR4_X1 U726 ( .A1(n1000), .A2(n1001), .A3(G953), .A4(n999), .ZN(n996) );
AND4_X1 U727 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n999) );
NOR4_X1 U728 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1005) );
XNOR2_X1 U729 ( .A(G478), .B(n1010), .ZN(n1009) );
XOR2_X1 U730 ( .A(KEYINPUT30), .B(n1011), .Z(n1008) );
XOR2_X1 U731 ( .A(KEYINPUT39), .B(n1012), .Z(n1007) );
NOR3_X1 U732 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U734 ( .A1(KEYINPUT63), .A2(n1018), .ZN(n1017) );
XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n1019), .ZN(n1018) );
INV_X1 U736 ( .A(n1020), .ZN(n1016) );
NOR3_X1 U737 ( .A1(n1020), .A2(KEYINPUT63), .A3(n1019), .ZN(n1014) );
AND2_X1 U738 ( .A1(n1019), .A2(KEYINPUT63), .ZN(n1013) );
XNOR2_X1 U739 ( .A(G469), .B(KEYINPUT33), .ZN(n1019) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1004) );
XOR2_X1 U741 ( .A(n1023), .B(n1024), .Z(n1003) );
NAND2_X1 U742 ( .A1(KEYINPUT28), .A2(n1025), .ZN(n1024) );
XOR2_X1 U743 ( .A(n1026), .B(KEYINPUT42), .Z(n1002) );
NAND2_X1 U744 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
OR2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U746 ( .A1(G472), .A2(n1031), .A3(n1029), .ZN(n1027) );
INV_X1 U747 ( .A(KEYINPUT29), .ZN(n1029) );
AND4_X1 U748 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1001) );
NAND3_X1 U749 ( .A1(G952), .A2(n1036), .A3(n1037), .ZN(n1000) );
INV_X1 U750 ( .A(n1038), .ZN(n1037) );
NAND3_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NAND3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1035), .ZN(n1043) );
INV_X1 U754 ( .A(KEYINPUT4), .ZN(n1045) );
INV_X1 U755 ( .A(n1032), .ZN(n1042) );
NAND3_X1 U756 ( .A1(n1046), .A2(n1047), .A3(n1032), .ZN(n1039) );
NAND2_X1 U757 ( .A1(n1035), .A2(n1048), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U759 ( .A1(KEYINPUT4), .A2(n1044), .ZN(n1050) );
INV_X1 U760 ( .A(n1051), .ZN(n1049) );
AND2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(n1035) );
NAND2_X1 U762 ( .A1(n1034), .A2(n1054), .ZN(n1046) );
NAND4_X1 U763 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND3_X1 U764 ( .A1(n1022), .A2(n1052), .A3(n1059), .ZN(n1057) );
XOR2_X1 U765 ( .A(KEYINPUT59), .B(n1060), .Z(n1059) );
NAND3_X1 U766 ( .A1(n1053), .A2(n1061), .A3(n1021), .ZN(n1056) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(n1055) );
XOR2_X1 U768 ( .A(n1053), .B(KEYINPUT54), .Z(n1063) );
XOR2_X1 U769 ( .A(n1064), .B(n1065), .Z(G72) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U772 ( .A(n1070), .ZN(n1069) );
XNOR2_X1 U773 ( .A(KEYINPUT8), .B(n1071), .ZN(n1068) );
NOR2_X1 U774 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NAND2_X1 U775 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
XNOR2_X1 U778 ( .A(n1078), .B(n1079), .ZN(n1076) );
XOR2_X1 U779 ( .A(n1080), .B(n1081), .Z(n1078) );
NOR2_X1 U780 ( .A1(KEYINPUT22), .A2(n1082), .ZN(n1081) );
XNOR2_X1 U781 ( .A(n1083), .B(n1084), .ZN(n1082) );
XOR2_X1 U782 ( .A(G137), .B(n1085), .Z(n1084) );
NAND2_X1 U783 ( .A1(G953), .A2(n1086), .ZN(n1064) );
NAND2_X1 U784 ( .A1(G900), .A2(G227), .ZN(n1086) );
XOR2_X1 U785 ( .A(n1087), .B(n1088), .Z(G69) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U787 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
NAND2_X1 U788 ( .A1(n1093), .A2(n1072), .ZN(n1092) );
NAND2_X1 U789 ( .A1(G953), .A2(n1094), .ZN(n1091) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1094) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1096), .ZN(G66) );
XNOR2_X1 U792 ( .A(n1097), .B(n1098), .ZN(n1096) );
NOR3_X1 U793 ( .A1(n1099), .A2(KEYINPUT31), .A3(n1100), .ZN(n1098) );
NOR2_X1 U794 ( .A1(n1095), .A2(n1101), .ZN(G63) );
XOR2_X1 U795 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U796 ( .A1(n1104), .A2(G478), .ZN(n1102) );
NOR2_X1 U797 ( .A1(n1095), .A2(n1105), .ZN(G60) );
XOR2_X1 U798 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U799 ( .A1(n1104), .A2(G475), .ZN(n1106) );
XNOR2_X1 U800 ( .A(G104), .B(n1108), .ZN(G6) );
NAND2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U802 ( .A(n1111), .B(KEYINPUT6), .Z(n1109) );
NOR2_X1 U803 ( .A1(n1095), .A2(n1112), .ZN(G57) );
XOR2_X1 U804 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U805 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND4_X1 U807 ( .A1(n1104), .A2(G472), .A3(n1119), .A4(n1120), .ZN(n1118) );
XOR2_X1 U808 ( .A(n1121), .B(KEYINPUT24), .Z(n1117) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U810 ( .A1(n1119), .A2(n1120), .ZN(n1123) );
NAND3_X1 U811 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1120) );
NAND3_X1 U812 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1125) );
OR2_X1 U813 ( .A1(n1129), .A2(n1128), .ZN(n1124) );
NAND2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1119) );
XOR2_X1 U815 ( .A(n1132), .B(n1128), .Z(n1131) );
NAND2_X1 U816 ( .A1(n1127), .A2(n1129), .ZN(n1132) );
INV_X1 U817 ( .A(KEYINPUT20), .ZN(n1129) );
NAND2_X1 U818 ( .A1(n1104), .A2(G472), .ZN(n1122) );
NAND2_X1 U819 ( .A1(KEYINPUT47), .A2(G101), .ZN(n1113) );
NOR2_X1 U820 ( .A1(n1095), .A2(n1133), .ZN(G54) );
XOR2_X1 U821 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U822 ( .A(n1136), .B(n1137), .ZN(n1135) );
XOR2_X1 U823 ( .A(n1138), .B(n1139), .Z(n1134) );
XOR2_X1 U824 ( .A(n1140), .B(KEYINPUT56), .Z(n1139) );
NAND2_X1 U825 ( .A1(KEYINPUT16), .A2(n1141), .ZN(n1140) );
XOR2_X1 U826 ( .A(KEYINPUT5), .B(G140), .Z(n1141) );
NAND2_X1 U827 ( .A1(n1104), .A2(G469), .ZN(n1138) );
NOR2_X1 U828 ( .A1(n1095), .A2(n1142), .ZN(G51) );
XOR2_X1 U829 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U830 ( .A(n1145), .B(n1146), .Z(n1143) );
NOR2_X1 U831 ( .A1(KEYINPUT52), .A2(n1128), .ZN(n1146) );
NAND2_X1 U832 ( .A1(n1104), .A2(n1147), .ZN(n1145) );
INV_X1 U833 ( .A(n1099), .ZN(n1104) );
NAND2_X1 U834 ( .A1(n1148), .A2(n1038), .ZN(n1099) );
NAND3_X1 U835 ( .A1(n1074), .A2(n1149), .A3(n1150), .ZN(n1038) );
INV_X1 U836 ( .A(n1093), .ZN(n1150) );
NAND4_X1 U837 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1093) );
AND3_X1 U838 ( .A1(n1155), .A2(n995), .A3(n1156), .ZN(n1154) );
NAND2_X1 U839 ( .A1(n1110), .A2(n1157), .ZN(n995) );
NAND2_X1 U840 ( .A1(n1158), .A2(n1110), .ZN(n1153) );
AND2_X1 U841 ( .A1(n1034), .A2(n1159), .ZN(n1110) );
NAND3_X1 U842 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1151) );
NAND2_X1 U843 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
NAND2_X1 U844 ( .A1(n1044), .A2(n1033), .ZN(n1164) );
OR2_X1 U845 ( .A1(n1158), .A2(n1157), .ZN(n1033) );
XOR2_X1 U846 ( .A(KEYINPUT15), .B(n1075), .Z(n1149) );
AND4_X1 U847 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1075) );
AND4_X1 U848 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1074) );
NAND4_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1053), .ZN(n1169) );
XNOR2_X1 U850 ( .A(n1062), .B(KEYINPUT18), .ZN(n1173) );
XOR2_X1 U851 ( .A(KEYINPUT19), .B(G902), .Z(n1148) );
NOR2_X1 U852 ( .A1(n1072), .A2(G952), .ZN(n1095) );
XOR2_X1 U853 ( .A(n1176), .B(n1177), .Z(G48) );
NAND2_X1 U854 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U855 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NAND2_X1 U856 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
OR2_X1 U857 ( .A1(n1171), .A2(n1182), .ZN(n1178) );
INV_X1 U858 ( .A(KEYINPUT49), .ZN(n1182) );
NAND3_X1 U859 ( .A1(n1184), .A2(n1180), .A3(n1183), .ZN(n1171) );
NOR3_X1 U860 ( .A1(n1111), .A2(n1185), .A3(n1186), .ZN(n1183) );
NAND2_X1 U861 ( .A1(KEYINPUT48), .A2(n1187), .ZN(n1176) );
XOR2_X1 U862 ( .A(n1188), .B(n1172), .Z(G45) );
NAND4_X1 U863 ( .A1(n1044), .A2(n1006), .A3(n1180), .A4(n1189), .ZN(n1172) );
NOR2_X1 U864 ( .A1(n1186), .A2(n1190), .ZN(n1189) );
XOR2_X1 U865 ( .A(n1191), .B(n1170), .Z(G42) );
NAND3_X1 U866 ( .A1(n1158), .A2(n1051), .A3(n1192), .ZN(n1170) );
NAND2_X1 U867 ( .A1(n1193), .A2(n1194), .ZN(G39) );
NAND4_X1 U868 ( .A1(n1174), .A2(n1192), .A3(n1195), .A4(n1196), .ZN(n1194) );
NAND2_X1 U869 ( .A1(G137), .A2(n1197), .ZN(n1196) );
NAND2_X1 U870 ( .A1(KEYINPUT2), .A2(n1198), .ZN(n1195) );
NAND3_X1 U871 ( .A1(n1199), .A2(n1197), .A3(G137), .ZN(n1193) );
INV_X1 U872 ( .A(KEYINPUT37), .ZN(n1197) );
NAND3_X1 U873 ( .A1(n1192), .A2(n1200), .A3(n1174), .ZN(n1199) );
INV_X1 U874 ( .A(KEYINPUT2), .ZN(n1200) );
XNOR2_X1 U875 ( .A(G134), .B(n1165), .ZN(G36) );
NAND3_X1 U876 ( .A1(n1157), .A2(n1044), .A3(n1192), .ZN(n1165) );
XOR2_X1 U877 ( .A(n1166), .B(n1201), .Z(G33) );
NAND2_X1 U878 ( .A1(KEYINPUT1), .A2(G131), .ZN(n1201) );
NAND3_X1 U879 ( .A1(n1158), .A2(n1044), .A3(n1192), .ZN(n1166) );
AND2_X1 U880 ( .A1(n1202), .A2(n1053), .ZN(n1192) );
NAND2_X1 U881 ( .A1(n1203), .A2(n1204), .ZN(n1053) );
OR3_X1 U882 ( .A1(n1205), .A2(n1022), .A3(KEYINPUT59), .ZN(n1204) );
INV_X1 U883 ( .A(n1060), .ZN(n1205) );
NAND2_X1 U884 ( .A1(KEYINPUT59), .A2(n1180), .ZN(n1203) );
XOR2_X1 U885 ( .A(n1206), .B(n1167), .Z(G30) );
NAND3_X1 U886 ( .A1(n1184), .A2(n1202), .A3(n1207), .ZN(n1167) );
AND3_X1 U887 ( .A1(n1157), .A2(n1011), .A3(n1180), .ZN(n1207) );
INV_X1 U888 ( .A(n1186), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1175), .A2(n1062), .ZN(n1186) );
XOR2_X1 U890 ( .A(n1208), .B(n1152), .Z(G3) );
NAND3_X1 U891 ( .A1(n1159), .A2(n1044), .A3(n1041), .ZN(n1152) );
NAND3_X1 U892 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(G27) );
NAND2_X1 U893 ( .A1(G125), .A2(n1212), .ZN(n1211) );
OR3_X1 U894 ( .A1(n1212), .A2(G125), .A3(n1168), .ZN(n1210) );
INV_X1 U895 ( .A(KEYINPUT7), .ZN(n1212) );
NAND2_X1 U896 ( .A1(n1213), .A2(n1168), .ZN(n1209) );
NAND4_X1 U897 ( .A1(n1175), .A2(n1158), .A3(n1162), .A4(n1051), .ZN(n1168) );
INV_X1 U898 ( .A(n1111), .ZN(n1158) );
AND2_X1 U899 ( .A1(n1032), .A2(n1214), .ZN(n1175) );
NAND2_X1 U900 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U901 ( .A1(n1077), .A2(G902), .ZN(n1215) );
NOR2_X1 U902 ( .A1(n1217), .A2(G900), .ZN(n1077) );
NAND2_X1 U903 ( .A1(n1218), .A2(KEYINPUT7), .ZN(n1213) );
XNOR2_X1 U904 ( .A(G125), .B(KEYINPUT34), .ZN(n1218) );
XOR2_X1 U905 ( .A(n1155), .B(n1219), .Z(G24) );
XOR2_X1 U906 ( .A(KEYINPUT51), .B(G122), .Z(n1219) );
NAND4_X1 U907 ( .A1(n1160), .A2(n1006), .A3(n1034), .A4(n1220), .ZN(n1155) );
NOR2_X1 U908 ( .A1(n1058), .A2(n1190), .ZN(n1220) );
XOR2_X1 U909 ( .A(n1221), .B(n1222), .Z(G21) );
NAND4_X1 U910 ( .A1(KEYINPUT61), .A2(n1174), .A3(n1162), .A4(n1160), .ZN(n1222) );
INV_X1 U911 ( .A(n1163), .ZN(n1174) );
NAND3_X1 U912 ( .A1(n1041), .A2(n1011), .A3(n1184), .ZN(n1163) );
XOR2_X1 U913 ( .A(n1223), .B(n1030), .Z(n1184) );
XOR2_X1 U914 ( .A(n1224), .B(n1225), .Z(G18) );
NAND4_X1 U915 ( .A1(n1162), .A2(n1157), .A3(n1226), .A4(n1044), .ZN(n1225) );
XOR2_X1 U916 ( .A(KEYINPUT17), .B(n1160), .Z(n1226) );
NOR2_X1 U917 ( .A1(n1190), .A2(n1006), .ZN(n1157) );
INV_X1 U918 ( .A(n1058), .ZN(n1162) );
NAND2_X1 U919 ( .A1(n1052), .A2(n1180), .ZN(n1058) );
INV_X1 U920 ( .A(n1227), .ZN(n1052) );
XOR2_X1 U921 ( .A(n1228), .B(n1229), .Z(G15) );
NAND4_X1 U922 ( .A1(n1230), .A2(n1044), .A3(n1160), .A4(n1231), .ZN(n1229) );
NOR2_X1 U923 ( .A1(n1227), .A2(n1111), .ZN(n1231) );
NAND2_X1 U924 ( .A1(n1006), .A2(n1190), .ZN(n1111) );
INV_X1 U925 ( .A(n1232), .ZN(n1190) );
NAND2_X1 U926 ( .A1(n1061), .A2(n1233), .ZN(n1227) );
NAND2_X1 U927 ( .A1(n1234), .A2(n1235), .ZN(n1044) );
NAND2_X1 U928 ( .A1(n1034), .A2(n1223), .ZN(n1235) );
INV_X1 U929 ( .A(KEYINPUT10), .ZN(n1223) );
NOR2_X1 U930 ( .A1(n1030), .A2(n1011), .ZN(n1034) );
INV_X1 U931 ( .A(n1185), .ZN(n1011) );
NAND3_X1 U932 ( .A1(n1030), .A2(n1185), .A3(KEYINPUT10), .ZN(n1234) );
XOR2_X1 U933 ( .A(KEYINPUT53), .B(n1180), .Z(n1230) );
XOR2_X1 U934 ( .A(n1156), .B(n1236), .Z(G12) );
XOR2_X1 U935 ( .A(n1237), .B(KEYINPUT57), .Z(n1236) );
NAND3_X1 U936 ( .A1(n1051), .A2(n1159), .A3(n1041), .ZN(n1156) );
NOR2_X1 U937 ( .A1(n1006), .A2(n1232), .ZN(n1041) );
XOR2_X1 U938 ( .A(n1010), .B(n1238), .Z(n1232) );
NOR2_X1 U939 ( .A1(G478), .A2(KEYINPUT9), .ZN(n1238) );
NAND2_X1 U940 ( .A1(n1103), .A2(n1239), .ZN(n1010) );
XOR2_X1 U941 ( .A(n1240), .B(n1241), .Z(n1103) );
XOR2_X1 U942 ( .A(G116), .B(n1242), .Z(n1241) );
XOR2_X1 U943 ( .A(G143), .B(G128), .Z(n1242) );
XOR2_X1 U944 ( .A(n1243), .B(n1085), .Z(n1240) );
XOR2_X1 U945 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND3_X1 U946 ( .A1(G217), .A2(n1072), .A3(n1246), .ZN(n1244) );
XNOR2_X1 U947 ( .A(G234), .B(KEYINPUT50), .ZN(n1246) );
XNOR2_X1 U948 ( .A(n1247), .B(G475), .ZN(n1006) );
NAND2_X1 U949 ( .A1(n1107), .A2(n1239), .ZN(n1247) );
XOR2_X1 U950 ( .A(n1248), .B(n1249), .Z(n1107) );
XOR2_X1 U951 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U952 ( .A(G131), .B(n1252), .Z(n1251) );
NOR3_X1 U953 ( .A1(n1253), .A2(KEYINPUT35), .A3(n1254), .ZN(n1252) );
NOR2_X1 U954 ( .A1(G104), .A2(n1255), .ZN(n1254) );
XOR2_X1 U955 ( .A(n1256), .B(KEYINPUT55), .Z(n1253) );
NAND2_X1 U956 ( .A1(G104), .A2(n1255), .ZN(n1256) );
XNOR2_X1 U957 ( .A(G122), .B(n1228), .ZN(n1255) );
AND2_X1 U958 ( .A1(n1257), .A2(G214), .ZN(n1250) );
XOR2_X1 U959 ( .A(n1258), .B(n1259), .Z(n1248) );
NOR2_X1 U960 ( .A1(G125), .A2(KEYINPUT26), .ZN(n1259) );
AND3_X1 U961 ( .A1(n1180), .A2(n1160), .A3(n1062), .ZN(n1159) );
NOR2_X1 U962 ( .A1(n1061), .A2(n1021), .ZN(n1062) );
INV_X1 U963 ( .A(n1233), .ZN(n1021) );
NAND2_X1 U964 ( .A1(G221), .A2(n1260), .ZN(n1233) );
XNOR2_X1 U965 ( .A(n1020), .B(n1261), .ZN(n1061) );
NOR2_X1 U966 ( .A1(G469), .A2(KEYINPUT32), .ZN(n1261) );
NAND2_X1 U967 ( .A1(n1262), .A2(n1239), .ZN(n1020) );
XOR2_X1 U968 ( .A(n1137), .B(n1263), .Z(n1262) );
INV_X1 U969 ( .A(n1080), .ZN(n1263) );
XOR2_X1 U970 ( .A(n1258), .B(KEYINPUT56), .Z(n1080) );
XOR2_X1 U971 ( .A(n1191), .B(n1136), .Z(n1258) );
INV_X1 U972 ( .A(G140), .ZN(n1191) );
XOR2_X1 U973 ( .A(n1264), .B(n1265), .Z(n1137) );
XOR2_X1 U974 ( .A(G101), .B(n1266), .Z(n1265) );
XOR2_X1 U975 ( .A(KEYINPUT25), .B(G107), .Z(n1266) );
XNOR2_X1 U976 ( .A(n1267), .B(n1268), .ZN(n1264) );
XOR2_X1 U977 ( .A(n1269), .B(n1270), .Z(n1268) );
AND2_X1 U978 ( .A1(n1072), .A2(G227), .ZN(n1269) );
AND2_X1 U979 ( .A1(n1271), .A2(n1032), .ZN(n1160) );
NAND2_X1 U980 ( .A1(n1272), .A2(G234), .ZN(n1032) );
XNOR2_X1 U981 ( .A(G237), .B(KEYINPUT44), .ZN(n1272) );
NAND2_X1 U982 ( .A1(n1216), .A2(n1273), .ZN(n1271) );
NAND2_X1 U983 ( .A1(G902), .A2(n1089), .ZN(n1273) );
NOR2_X1 U984 ( .A1(n1217), .A2(G898), .ZN(n1089) );
XOR2_X1 U985 ( .A(G953), .B(KEYINPUT43), .Z(n1217) );
NAND2_X1 U986 ( .A1(n1274), .A2(G952), .ZN(n1216) );
XOR2_X1 U987 ( .A(n1072), .B(KEYINPUT14), .Z(n1274) );
NOR2_X1 U988 ( .A1(n1060), .A2(n1022), .ZN(n1180) );
AND2_X1 U989 ( .A1(G214), .A2(n1275), .ZN(n1022) );
XOR2_X1 U990 ( .A(n1025), .B(n1147), .Z(n1060) );
INV_X1 U991 ( .A(n1023), .ZN(n1147) );
NAND2_X1 U992 ( .A1(G210), .A2(n1275), .ZN(n1023) );
NAND2_X1 U993 ( .A1(n1276), .A2(n1239), .ZN(n1275) );
XOR2_X1 U994 ( .A(KEYINPUT58), .B(G237), .Z(n1276) );
NAND2_X1 U995 ( .A1(n1277), .A2(n1239), .ZN(n1025) );
XOR2_X1 U996 ( .A(n1278), .B(n1144), .Z(n1277) );
XNOR2_X1 U997 ( .A(n1090), .B(n1279), .ZN(n1144) );
XOR2_X1 U998 ( .A(G125), .B(n1280), .Z(n1279) );
AND2_X1 U999 ( .A1(n1072), .A2(G224), .ZN(n1280) );
XOR2_X1 U1000 ( .A(n1281), .B(n1282), .Z(n1090) );
XOR2_X1 U1001 ( .A(n1245), .B(n1270), .Z(n1282) );
XOR2_X1 U1002 ( .A(G110), .B(G104), .Z(n1270) );
XOR2_X1 U1003 ( .A(G107), .B(G122), .Z(n1245) );
XOR2_X1 U1004 ( .A(n1283), .B(n1284), .Z(n1281) );
NOR2_X1 U1005 ( .A1(KEYINPUT23), .A2(n1208), .ZN(n1284) );
INV_X1 U1006 ( .A(G101), .ZN(n1208) );
XOR2_X1 U1007 ( .A(n1285), .B(G113), .Z(n1283) );
NAND3_X1 U1008 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1285) );
OR2_X1 U1009 ( .A1(G116), .A2(KEYINPUT27), .ZN(n1288) );
NAND3_X1 U1010 ( .A1(KEYINPUT27), .A2(G116), .A3(n1221), .ZN(n1287) );
NAND2_X1 U1011 ( .A1(G119), .A2(n1289), .ZN(n1286) );
NAND2_X1 U1012 ( .A1(n1290), .A2(KEYINPUT27), .ZN(n1289) );
XOR2_X1 U1013 ( .A(n1224), .B(KEYINPUT41), .Z(n1290) );
INV_X1 U1014 ( .A(G116), .ZN(n1224) );
NAND2_X1 U1015 ( .A1(KEYINPUT12), .A2(n1128), .ZN(n1278) );
NOR2_X1 U1016 ( .A1(n1030), .A2(n1185), .ZN(n1051) );
XNOR2_X1 U1017 ( .A(n1291), .B(n1100), .ZN(n1185) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1260), .ZN(n1100) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1239), .ZN(n1260) );
NAND2_X1 U1020 ( .A1(n1097), .A2(n1239), .ZN(n1291) );
XNOR2_X1 U1021 ( .A(n1292), .B(n1293), .ZN(n1097) );
XOR2_X1 U1022 ( .A(G137), .B(n1294), .Z(n1293) );
NOR2_X1 U1023 ( .A1(KEYINPUT40), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1024 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1025 ( .A(G119), .B(n1298), .Z(n1297) );
XOR2_X1 U1026 ( .A(G146), .B(G140), .Z(n1298) );
XOR2_X1 U1027 ( .A(n1237), .B(n1079), .Z(n1296) );
XOR2_X1 U1028 ( .A(G128), .B(G125), .Z(n1079) );
INV_X1 U1029 ( .A(G110), .ZN(n1237) );
NAND4_X1 U1030 ( .A1(KEYINPUT62), .A2(G221), .A3(G234), .A4(n1072), .ZN(n1292) );
INV_X1 U1031 ( .A(G953), .ZN(n1072) );
XNOR2_X1 U1032 ( .A(G472), .B(n1031), .ZN(n1030) );
NAND2_X1 U1033 ( .A1(n1239), .A2(n1299), .ZN(n1031) );
NAND2_X1 U1034 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U1035 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1036 ( .A(KEYINPUT11), .B(n1304), .Z(n1300) );
NOR2_X1 U1037 ( .A1(n1303), .A2(n1302), .ZN(n1304) );
XOR2_X1 U1038 ( .A(n1115), .B(G101), .Z(n1302) );
NAND2_X1 U1039 ( .A1(G210), .A2(n1257), .ZN(n1115) );
NOR2_X1 U1040 ( .A1(G953), .A2(G237), .ZN(n1257) );
AND2_X1 U1041 ( .A1(n1305), .A2(n1306), .ZN(n1303) );
NAND2_X1 U1042 ( .A1(n1130), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1043 ( .A(n1308), .B(n1267), .Z(n1307) );
XNOR2_X1 U1044 ( .A(n1127), .B(n1206), .ZN(n1267) );
NAND2_X1 U1045 ( .A1(n1126), .A2(n1309), .ZN(n1305) );
NAND2_X1 U1046 ( .A1(n1128), .A2(n1127), .ZN(n1309) );
NOR2_X1 U1047 ( .A1(n1130), .A2(n1310), .ZN(n1126) );
NOR2_X1 U1048 ( .A1(n1127), .A2(n1128), .ZN(n1310) );
XOR2_X1 U1049 ( .A(n1206), .B(n1308), .Z(n1128) );
XNOR2_X1 U1050 ( .A(n1311), .B(KEYINPUT3), .ZN(n1308) );
NAND2_X1 U1051 ( .A1(KEYINPUT38), .A2(n1136), .ZN(n1311) );
XOR2_X1 U1052 ( .A(n1188), .B(n1187), .Z(n1136) );
INV_X1 U1053 ( .A(G146), .ZN(n1187) );
INV_X1 U1054 ( .A(G143), .ZN(n1188) );
INV_X1 U1055 ( .A(G128), .ZN(n1206) );
XNOR2_X1 U1056 ( .A(n1312), .B(n1313), .ZN(n1127) );
XOR2_X1 U1057 ( .A(n1198), .B(n1314), .Z(n1313) );
NAND2_X1 U1058 ( .A1(KEYINPUT46), .A2(n1085), .ZN(n1314) );
XOR2_X1 U1059 ( .A(G134), .B(KEYINPUT36), .Z(n1085) );
INV_X1 U1060 ( .A(G137), .ZN(n1198) );
NAND2_X1 U1061 ( .A1(KEYINPUT45), .A2(n1083), .ZN(n1312) );
XNOR2_X1 U1062 ( .A(G131), .B(KEYINPUT13), .ZN(n1083) );
XOR2_X1 U1063 ( .A(n1315), .B(n1316), .Z(n1130) );
NOR2_X1 U1064 ( .A1(KEYINPUT60), .A2(n1228), .ZN(n1316) );
INV_X1 U1065 ( .A(G113), .ZN(n1228) );
XOR2_X1 U1066 ( .A(n1221), .B(G116), .Z(n1315) );
INV_X1 U1067 ( .A(G119), .ZN(n1221) );
INV_X1 U1068 ( .A(G902), .ZN(n1239) );
endmodule


