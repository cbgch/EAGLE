//Key = 1101100101011011010110001001001111000010000010010111110011111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;

XNOR2_X1 U719 ( .A(n1000), .B(n1001), .ZN(G9) );
NAND2_X1 U720 ( .A1(KEYINPUT11), .A2(n1002), .ZN(n1000) );
NOR2_X1 U721 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U722 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
XOR2_X1 U723 ( .A(n1009), .B(KEYINPUT56), .Z(n1008) );
NAND4_X1 U724 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
AND2_X1 U725 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U726 ( .A1(n1016), .A2(n1017), .ZN(n1007) );
INV_X1 U727 ( .A(n1018), .ZN(n1017) );
NOR3_X1 U728 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1016) );
NOR2_X1 U729 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
INV_X1 U730 ( .A(KEYINPUT5), .ZN(n1023) );
AND2_X1 U731 ( .A1(n1024), .A2(n1014), .ZN(n1022) );
NOR4_X1 U732 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1020) );
NOR2_X1 U733 ( .A1(n1029), .A2(n1030), .ZN(n1026) );
NOR2_X1 U734 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U735 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U736 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U737 ( .A1(n1037), .A2(KEYINPUT5), .A3(n1038), .ZN(n1029) );
XOR2_X1 U738 ( .A(KEYINPUT46), .B(n1039), .Z(n1019) );
AND2_X1 U739 ( .A1(n1040), .A2(n1014), .ZN(n1039) );
INV_X1 U740 ( .A(n1041), .ZN(n1006) );
NAND3_X1 U741 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1005) );
NAND2_X1 U742 ( .A1(n1014), .A2(n1045), .ZN(n1044) );
NAND2_X1 U743 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U744 ( .A1(n1010), .A2(n1048), .ZN(n1047) );
NAND2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U747 ( .A(KEYINPUT14), .B(n1011), .ZN(n1051) );
NAND2_X1 U748 ( .A1(n1018), .A2(n1053), .ZN(n1049) );
NAND2_X1 U749 ( .A1(n1054), .A2(n1011), .ZN(n1046) );
NOR3_X1 U750 ( .A1(n1037), .A2(n1025), .A3(n1028), .ZN(n1014) );
INV_X1 U751 ( .A(KEYINPUT50), .ZN(n1028) );
INV_X1 U752 ( .A(n1055), .ZN(n1037) );
NOR3_X1 U753 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1003) );
INV_X1 U754 ( .A(n1042), .ZN(n1056) );
NAND2_X1 U755 ( .A1(n1057), .A2(n1058), .ZN(n1042) );
NOR4_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
XNOR2_X1 U757 ( .A(n1012), .B(KEYINPUT9), .ZN(n1062) );
XOR2_X1 U758 ( .A(n1063), .B(n1064), .Z(n1061) );
NOR2_X1 U759 ( .A1(G472), .A2(KEYINPUT29), .ZN(n1064) );
XOR2_X1 U760 ( .A(n1065), .B(n1066), .Z(n1060) );
NAND2_X1 U761 ( .A1(KEYINPUT47), .A2(n1067), .ZN(n1065) );
NOR4_X1 U762 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1057) );
XOR2_X1 U763 ( .A(G469), .B(n1072), .Z(n1071) );
XNOR2_X1 U764 ( .A(n1073), .B(n1074), .ZN(n1070) );
XOR2_X1 U765 ( .A(n1075), .B(n1076), .Z(G72) );
NOR2_X1 U766 ( .A1(n1077), .A2(n1043), .ZN(n1076) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U770 ( .A(n1082), .B(KEYINPUT37), .Z(n1080) );
XOR2_X1 U771 ( .A(KEYINPUT52), .B(n1083), .Z(n1078) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1082), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U775 ( .A(n1089), .B(n1090), .Z(n1085) );
XNOR2_X1 U776 ( .A(n1091), .B(n1092), .ZN(n1090) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1089) );
XNOR2_X1 U778 ( .A(G134), .B(G128), .ZN(n1093) );
XNOR2_X1 U779 ( .A(n1081), .B(KEYINPUT24), .ZN(n1084) );
AND2_X1 U780 ( .A1(n1043), .A2(n1095), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1096), .B(n1097), .Z(G69) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(n1097) );
AND2_X1 U783 ( .A1(n1100), .A2(n1043), .ZN(n1099) );
NOR2_X1 U784 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
AND2_X1 U785 ( .A1(n1103), .A2(n1087), .ZN(n1101) );
NOR2_X1 U786 ( .A1(n1104), .A2(n1043), .ZN(n1096) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1103), .ZN(n1104) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U789 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U790 ( .A1(n1110), .A2(G217), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1106), .A2(n1111), .ZN(G63) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U793 ( .A(KEYINPUT40), .B(n1114), .Z(n1113) );
NOR2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n1117), .ZN(n1116) );
INV_X1 U796 ( .A(n1118), .ZN(n1115) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1110), .A2(G478), .ZN(n1117) );
NOR2_X1 U799 ( .A1(n1106), .A2(n1119), .ZN(G60) );
NOR3_X1 U800 ( .A1(n1066), .A2(n1120), .A3(n1121), .ZN(n1119) );
AND3_X1 U801 ( .A1(n1122), .A2(G475), .A3(n1110), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1122), .ZN(n1120) );
NOR2_X1 U803 ( .A1(n1041), .A2(n1067), .ZN(n1123) );
XOR2_X1 U804 ( .A(G104), .B(n1124), .Z(G6) );
NOR2_X1 U805 ( .A1(n1106), .A2(n1125), .ZN(G57) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U809 ( .A(n1132), .B(KEYINPUT7), .ZN(n1131) );
NAND2_X1 U810 ( .A1(KEYINPUT20), .A2(n1133), .ZN(n1128) );
XNOR2_X1 U811 ( .A(n1134), .B(n1135), .ZN(n1133) );
XNOR2_X1 U812 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND2_X1 U813 ( .A1(n1110), .A2(G472), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1106), .A2(n1138), .ZN(G54) );
XOR2_X1 U815 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U818 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U819 ( .A(KEYINPUT32), .B(n1147), .Z(n1143) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1147) );
XNOR2_X1 U821 ( .A(n1148), .B(KEYINPUT12), .ZN(n1145) );
NAND2_X1 U822 ( .A1(n1149), .A2(KEYINPUT30), .ZN(n1141) );
XNOR2_X1 U823 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U824 ( .A1(n1110), .A2(G469), .ZN(n1139) );
NOR2_X1 U825 ( .A1(n1043), .A2(G952), .ZN(n1106) );
NOR2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(G51) );
XOR2_X1 U827 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U828 ( .A(n1156), .B(n1102), .Z(n1155) );
XNOR2_X1 U829 ( .A(n1157), .B(G101), .ZN(n1102) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1154) );
NOR2_X1 U831 ( .A1(KEYINPUT25), .A2(n1160), .ZN(n1159) );
NAND2_X1 U832 ( .A1(n1110), .A2(n1161), .ZN(n1158) );
INV_X1 U833 ( .A(n1074), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1162), .A2(n1041), .ZN(n1110) );
NOR2_X1 U835 ( .A1(n1095), .A2(n1100), .ZN(n1041) );
NAND4_X1 U836 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1100) );
AND4_X1 U837 ( .A1(n1002), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1166) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1040), .ZN(n1002) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1032), .ZN(n1040) );
NOR2_X1 U840 ( .A1(n1124), .A2(n1172), .ZN(n1165) );
NOR2_X1 U841 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
AND3_X1 U842 ( .A1(n1170), .A2(n1010), .A3(n1053), .ZN(n1124) );
NAND4_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1095) );
NOR4_X1 U844 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
INV_X1 U845 ( .A(n1183), .ZN(n1181) );
INV_X1 U846 ( .A(n1184), .ZN(n1179) );
OR2_X1 U847 ( .A1(n1185), .A2(n1173), .ZN(n1177) );
NAND2_X1 U848 ( .A1(n1186), .A2(n1187), .ZN(n1175) );
NAND2_X1 U849 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
NAND3_X1 U850 ( .A1(n1190), .A2(n1191), .A3(n1054), .ZN(n1189) );
INV_X1 U851 ( .A(n1192), .ZN(n1054) );
XOR2_X1 U852 ( .A(KEYINPUT13), .B(n1034), .Z(n1191) );
NAND2_X1 U853 ( .A1(n1193), .A2(n1194), .ZN(n1188) );
XOR2_X1 U854 ( .A(KEYINPUT10), .B(n1034), .Z(n1194) );
INV_X1 U855 ( .A(n1195), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1196), .A2(n1043), .ZN(n1152) );
XNOR2_X1 U857 ( .A(G952), .B(KEYINPUT58), .ZN(n1196) );
XOR2_X1 U858 ( .A(n1197), .B(n1198), .Z(G48) );
NOR2_X1 U859 ( .A1(KEYINPUT45), .A2(n1199), .ZN(n1198) );
NOR2_X1 U860 ( .A1(n1200), .A2(n1195), .ZN(n1197) );
NAND3_X1 U861 ( .A1(n1201), .A2(n1052), .A3(n1053), .ZN(n1195) );
XNOR2_X1 U862 ( .A(G143), .B(n1176), .ZN(G45) );
NAND4_X1 U863 ( .A1(n1202), .A2(n1052), .A3(n1203), .A4(n1204), .ZN(n1176) );
AND2_X1 U864 ( .A1(n1069), .A2(n1205), .ZN(n1203) );
XOR2_X1 U865 ( .A(G140), .B(n1182), .Z(G42) );
AND2_X1 U866 ( .A1(n1206), .A2(n1207), .ZN(n1182) );
XOR2_X1 U867 ( .A(n1208), .B(G137), .Z(G39) );
NAND2_X1 U868 ( .A1(KEYINPUT62), .A2(n1183), .ZN(n1208) );
NAND3_X1 U869 ( .A1(n1202), .A2(n1018), .A3(n1209), .ZN(n1183) );
XOR2_X1 U870 ( .A(n1210), .B(n1211), .Z(G36) );
NOR3_X1 U871 ( .A1(n1192), .A2(n1171), .A3(n1200), .ZN(n1211) );
NAND2_X1 U872 ( .A1(n1018), .A2(n1204), .ZN(n1192) );
XNOR2_X1 U873 ( .A(G134), .B(KEYINPUT31), .ZN(n1210) );
XOR2_X1 U874 ( .A(G131), .B(n1180), .Z(G33) );
AND2_X1 U875 ( .A1(n1206), .A2(n1204), .ZN(n1180) );
AND3_X1 U876 ( .A1(n1018), .A2(n1053), .A3(n1202), .ZN(n1206) );
NOR2_X1 U877 ( .A1(n1212), .A2(n1012), .ZN(n1018) );
XOR2_X1 U878 ( .A(n1213), .B(n1214), .Z(G30) );
NOR2_X1 U879 ( .A1(KEYINPUT43), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U880 ( .A(G128), .B(KEYINPUT42), .ZN(n1215) );
NOR2_X1 U881 ( .A1(n1216), .A2(n1173), .ZN(n1213) );
INV_X1 U882 ( .A(n1052), .ZN(n1173) );
XOR2_X1 U883 ( .A(n1185), .B(KEYINPUT54), .Z(n1216) );
NAND3_X1 U884 ( .A1(n1201), .A2(n1190), .A3(n1202), .ZN(n1185) );
INV_X1 U885 ( .A(n1200), .ZN(n1202) );
NAND2_X1 U886 ( .A1(n1034), .A2(n1187), .ZN(n1200) );
XNOR2_X1 U887 ( .A(G101), .B(n1217), .ZN(G3) );
NAND3_X1 U888 ( .A1(KEYINPUT44), .A2(n1052), .A3(n1218), .ZN(n1217) );
XOR2_X1 U889 ( .A(n1174), .B(KEYINPUT27), .Z(n1218) );
NAND4_X1 U890 ( .A1(n1034), .A2(n1011), .A3(n1204), .A4(n1219), .ZN(n1174) );
XNOR2_X1 U891 ( .A(G125), .B(n1184), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1207), .A2(n1187), .A3(n1052), .A4(n1220), .ZN(n1184) );
AND2_X1 U893 ( .A1(n1055), .A2(n1053), .ZN(n1220) );
NAND2_X1 U894 ( .A1(n1221), .A2(n1222), .ZN(n1187) );
NAND4_X1 U895 ( .A1(G902), .A2(n1087), .A3(n1223), .A4(n1088), .ZN(n1222) );
INV_X1 U896 ( .A(G900), .ZN(n1088) );
XNOR2_X1 U897 ( .A(G122), .B(n1163), .ZN(G24) );
NAND4_X1 U898 ( .A1(n1224), .A2(n1010), .A3(n1205), .A4(n1069), .ZN(n1163) );
INV_X1 U899 ( .A(n1032), .ZN(n1010) );
NAND2_X1 U900 ( .A1(n1225), .A2(n1226), .ZN(n1032) );
XNOR2_X1 U901 ( .A(KEYINPUT6), .B(n1068), .ZN(n1226) );
XNOR2_X1 U902 ( .A(n1227), .B(n1228), .ZN(n1225) );
XNOR2_X1 U903 ( .A(G119), .B(n1164), .ZN(G21) );
NAND2_X1 U904 ( .A1(n1224), .A2(n1209), .ZN(n1164) );
AND2_X1 U905 ( .A1(n1201), .A2(n1011), .ZN(n1209) );
XNOR2_X1 U906 ( .A(G116), .B(n1169), .ZN(G18) );
NAND3_X1 U907 ( .A1(n1190), .A2(n1204), .A3(n1224), .ZN(n1169) );
INV_X1 U908 ( .A(n1171), .ZN(n1190) );
NAND2_X1 U909 ( .A1(n1229), .A2(n1069), .ZN(n1171) );
XNOR2_X1 U910 ( .A(n1205), .B(KEYINPUT22), .ZN(n1229) );
NAND2_X1 U911 ( .A1(n1230), .A2(n1231), .ZN(G15) );
NAND2_X1 U912 ( .A1(G113), .A2(n1168), .ZN(n1231) );
XOR2_X1 U913 ( .A(n1232), .B(KEYINPUT36), .Z(n1230) );
OR2_X1 U914 ( .A1(n1168), .A2(G113), .ZN(n1232) );
NAND3_X1 U915 ( .A1(n1053), .A2(n1204), .A3(n1224), .ZN(n1168) );
AND3_X1 U916 ( .A1(n1052), .A2(n1219), .A3(n1055), .ZN(n1224) );
NOR2_X1 U917 ( .A1(n1035), .A2(n1059), .ZN(n1055) );
INV_X1 U918 ( .A(n1036), .ZN(n1059) );
NAND2_X1 U919 ( .A1(n1233), .A2(n1234), .ZN(n1204) );
OR3_X1 U920 ( .A1(n1068), .A2(n1228), .A3(KEYINPUT6), .ZN(n1234) );
NAND2_X1 U921 ( .A1(KEYINPUT6), .A2(n1201), .ZN(n1233) );
XNOR2_X1 U922 ( .A(G110), .B(n1167), .ZN(G12) );
NAND2_X1 U923 ( .A1(n1024), .A2(n1170), .ZN(n1167) );
AND3_X1 U924 ( .A1(n1052), .A2(n1219), .A3(n1034), .ZN(n1170) );
AND2_X1 U925 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U926 ( .A1(G221), .A2(n1235), .ZN(n1036) );
NAND2_X1 U927 ( .A1(G234), .A2(n1162), .ZN(n1235) );
XNOR2_X1 U928 ( .A(G469), .B(n1236), .ZN(n1035) );
NOR2_X1 U929 ( .A1(n1072), .A2(KEYINPUT41), .ZN(n1236) );
AND2_X1 U930 ( .A1(n1237), .A2(n1162), .ZN(n1072) );
XOR2_X1 U931 ( .A(n1150), .B(n1238), .Z(n1237) );
XNOR2_X1 U932 ( .A(n1239), .B(n1240), .ZN(n1238) );
NOR2_X1 U933 ( .A1(KEYINPUT8), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U934 ( .A(n1146), .B(n1242), .ZN(n1241) );
INV_X1 U935 ( .A(n1148), .ZN(n1242) );
XOR2_X1 U936 ( .A(G110), .B(G140), .Z(n1148) );
NAND2_X1 U937 ( .A1(G227), .A2(n1043), .ZN(n1146) );
NAND2_X1 U938 ( .A1(KEYINPUT1), .A2(n1151), .ZN(n1239) );
XOR2_X1 U939 ( .A(n1243), .B(n1244), .Z(n1150) );
XNOR2_X1 U940 ( .A(n1001), .B(G104), .ZN(n1244) );
XOR2_X1 U941 ( .A(n1245), .B(n1092), .Z(n1243) );
XNOR2_X1 U942 ( .A(n1246), .B(KEYINPUT59), .ZN(n1092) );
NAND2_X1 U943 ( .A1(KEYINPUT57), .A2(n1247), .ZN(n1246) );
NAND2_X1 U944 ( .A1(n1221), .A2(n1248), .ZN(n1219) );
NAND4_X1 U945 ( .A1(G902), .A2(n1087), .A3(n1223), .A4(n1103), .ZN(n1248) );
INV_X1 U946 ( .A(G898), .ZN(n1103) );
XOR2_X1 U947 ( .A(G953), .B(KEYINPUT16), .Z(n1087) );
NAND3_X1 U948 ( .A1(n1223), .A2(n1043), .A3(G952), .ZN(n1221) );
INV_X1 U949 ( .A(n1025), .ZN(n1223) );
NOR2_X1 U950 ( .A1(n1249), .A2(n1250), .ZN(n1025) );
NOR2_X1 U951 ( .A1(n1015), .A2(n1012), .ZN(n1052) );
AND2_X1 U952 ( .A1(G214), .A2(n1251), .ZN(n1012) );
INV_X1 U953 ( .A(n1212), .ZN(n1015) );
NAND2_X1 U954 ( .A1(n1252), .A2(n1253), .ZN(n1212) );
NAND2_X1 U955 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XNOR2_X1 U956 ( .A(KEYINPUT21), .B(n1074), .ZN(n1254) );
NAND2_X1 U957 ( .A1(n1256), .A2(n1073), .ZN(n1252) );
INV_X1 U958 ( .A(n1255), .ZN(n1073) );
NAND2_X1 U959 ( .A1(n1257), .A2(n1162), .ZN(n1255) );
XOR2_X1 U960 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U961 ( .A(n1245), .B(n1156), .Z(n1259) );
XNOR2_X1 U962 ( .A(n1260), .B(n1261), .ZN(n1156) );
NOR2_X1 U963 ( .A1(G953), .A2(n1105), .ZN(n1261) );
INV_X1 U964 ( .A(G224), .ZN(n1105) );
XNOR2_X1 U965 ( .A(G101), .B(G128), .ZN(n1245) );
XOR2_X1 U966 ( .A(n1157), .B(n1247), .Z(n1258) );
XOR2_X1 U967 ( .A(n1262), .B(n1263), .Z(n1157) );
XNOR2_X1 U968 ( .A(n1264), .B(n1265), .ZN(n1263) );
INV_X1 U969 ( .A(n1137), .ZN(n1265) );
NOR2_X1 U970 ( .A1(KEYINPUT48), .A2(n1266), .ZN(n1264) );
XNOR2_X1 U971 ( .A(G104), .B(n1267), .ZN(n1266) );
NOR2_X1 U972 ( .A1(KEYINPUT23), .A2(n1001), .ZN(n1267) );
XNOR2_X1 U973 ( .A(G110), .B(n1268), .ZN(n1262) );
XOR2_X1 U974 ( .A(KEYINPUT18), .B(G122), .Z(n1268) );
XNOR2_X1 U975 ( .A(KEYINPUT49), .B(n1074), .ZN(n1256) );
NAND2_X1 U976 ( .A1(G210), .A2(n1251), .ZN(n1074) );
NAND2_X1 U977 ( .A1(n1249), .A2(n1162), .ZN(n1251) );
INV_X1 U978 ( .A(G237), .ZN(n1249) );
NOR2_X1 U979 ( .A1(n1027), .A2(n1038), .ZN(n1024) );
INV_X1 U980 ( .A(n1207), .ZN(n1038) );
NAND2_X1 U981 ( .A1(n1269), .A2(n1270), .ZN(n1207) );
NAND3_X1 U982 ( .A1(n1228), .A2(n1068), .A3(n1227), .ZN(n1270) );
INV_X1 U983 ( .A(KEYINPUT55), .ZN(n1227) );
NAND2_X1 U984 ( .A1(KEYINPUT55), .A2(n1201), .ZN(n1269) );
NOR2_X1 U985 ( .A1(n1228), .A2(n1271), .ZN(n1201) );
INV_X1 U986 ( .A(n1068), .ZN(n1271) );
NAND3_X1 U987 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1068) );
OR2_X1 U988 ( .A1(n1275), .A2(n1109), .ZN(n1274) );
NAND3_X1 U989 ( .A1(n1109), .A2(n1275), .A3(n1162), .ZN(n1273) );
NAND2_X1 U990 ( .A1(G217), .A2(n1250), .ZN(n1275) );
AND3_X1 U991 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1109) );
OR2_X1 U992 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND3_X1 U993 ( .A1(n1280), .A2(n1279), .A3(KEYINPUT60), .ZN(n1277) );
XNOR2_X1 U994 ( .A(n1281), .B(G137), .ZN(n1279) );
NAND3_X1 U995 ( .A1(G234), .A2(n1043), .A3(G221), .ZN(n1281) );
AND2_X1 U996 ( .A1(KEYINPUT15), .A2(n1282), .ZN(n1280) );
OR2_X1 U997 ( .A1(n1282), .A2(KEYINPUT60), .ZN(n1276) );
XOR2_X1 U998 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U999 ( .A(G119), .B(n1285), .Z(n1284) );
XNOR2_X1 U1000 ( .A(KEYINPUT28), .B(n1286), .ZN(n1285) );
INV_X1 U1001 ( .A(G128), .ZN(n1286) );
XNOR2_X1 U1002 ( .A(n1287), .B(n1288), .ZN(n1283) );
NAND2_X1 U1003 ( .A1(KEYINPUT53), .A2(n1289), .ZN(n1288) );
INV_X1 U1004 ( .A(G110), .ZN(n1289) );
NAND2_X1 U1005 ( .A1(KEYINPUT38), .A2(n1290), .ZN(n1287) );
XNOR2_X1 U1006 ( .A(n1199), .B(n1094), .ZN(n1290) );
XNOR2_X1 U1007 ( .A(n1260), .B(G140), .ZN(n1094) );
NAND2_X1 U1008 ( .A1(G217), .A2(G902), .ZN(n1272) );
XOR2_X1 U1009 ( .A(n1063), .B(G472), .Z(n1228) );
NAND2_X1 U1010 ( .A1(n1291), .A2(n1162), .ZN(n1063) );
XNOR2_X1 U1011 ( .A(n1137), .B(n1292), .ZN(n1291) );
XOR2_X1 U1012 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR3_X1 U1013 ( .A1(n1132), .A2(KEYINPUT39), .A3(n1130), .ZN(n1294) );
AND3_X1 U1014 ( .A1(G210), .A2(G101), .A3(n1295), .ZN(n1130) );
AND2_X1 U1015 ( .A1(n1296), .A2(n1297), .ZN(n1132) );
INV_X1 U1016 ( .A(G101), .ZN(n1297) );
NAND2_X1 U1017 ( .A1(n1295), .A2(G210), .ZN(n1296) );
NAND3_X1 U1018 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1293) );
NAND2_X1 U1019 ( .A1(n1160), .A2(n1301), .ZN(n1300) );
NAND2_X1 U1020 ( .A1(KEYINPUT4), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U1021 ( .A(KEYINPUT51), .B(n1151), .ZN(n1302) );
INV_X1 U1022 ( .A(n1134), .ZN(n1160) );
NAND3_X1 U1023 ( .A1(KEYINPUT4), .A2(n1134), .A3(n1151), .ZN(n1299) );
XOR2_X1 U1024 ( .A(G128), .B(n1247), .Z(n1134) );
XNOR2_X1 U1025 ( .A(n1303), .B(G146), .ZN(n1247) );
OR2_X1 U1026 ( .A1(n1151), .A2(KEYINPUT4), .ZN(n1298) );
INV_X1 U1027 ( .A(n1136), .ZN(n1151) );
XOR2_X1 U1028 ( .A(n1304), .B(n1305), .Z(n1136) );
INV_X1 U1029 ( .A(n1091), .ZN(n1305) );
XOR2_X1 U1030 ( .A(G131), .B(G137), .Z(n1091) );
NAND2_X1 U1031 ( .A1(KEYINPUT3), .A2(n1306), .ZN(n1304) );
XNOR2_X1 U1032 ( .A(n1307), .B(n1308), .ZN(n1137) );
XOR2_X1 U1033 ( .A(KEYINPUT26), .B(G119), .Z(n1308) );
XNOR2_X1 U1034 ( .A(G116), .B(G113), .ZN(n1307) );
INV_X1 U1035 ( .A(n1011), .ZN(n1027) );
NAND2_X1 U1036 ( .A1(n1309), .A2(n1310), .ZN(n1011) );
OR3_X1 U1037 ( .A1(n1205), .A2(n1069), .A3(KEYINPUT22), .ZN(n1310) );
INV_X1 U1038 ( .A(n1311), .ZN(n1205) );
NAND2_X1 U1039 ( .A1(KEYINPUT22), .A2(n1053), .ZN(n1309) );
NOR2_X1 U1040 ( .A1(n1069), .A2(n1311), .ZN(n1053) );
XOR2_X1 U1041 ( .A(n1066), .B(n1067), .Z(n1311) );
INV_X1 U1042 ( .A(G475), .ZN(n1067) );
NOR2_X1 U1043 ( .A1(n1122), .A2(G902), .ZN(n1066) );
XOR2_X1 U1044 ( .A(n1312), .B(n1313), .Z(n1122) );
XNOR2_X1 U1045 ( .A(G104), .B(n1314), .ZN(n1313) );
NAND2_X1 U1046 ( .A1(n1295), .A2(G214), .ZN(n1314) );
NOR2_X1 U1047 ( .A1(G953), .A2(G237), .ZN(n1295) );
XOR2_X1 U1048 ( .A(n1315), .B(n1316), .Z(n1312) );
XOR2_X1 U1049 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1050 ( .A(G140), .B(G131), .Z(n1318) );
XNOR2_X1 U1051 ( .A(KEYINPUT34), .B(n1199), .ZN(n1317) );
INV_X1 U1052 ( .A(G146), .ZN(n1199) );
XOR2_X1 U1053 ( .A(n1319), .B(n1320), .Z(n1315) );
XOR2_X1 U1054 ( .A(G122), .B(G113), .Z(n1320) );
XNOR2_X1 U1055 ( .A(n1321), .B(n1322), .ZN(n1319) );
NAND2_X1 U1056 ( .A1(KEYINPUT33), .A2(n1260), .ZN(n1322) );
INV_X1 U1057 ( .A(G125), .ZN(n1260) );
NAND2_X1 U1058 ( .A1(KEYINPUT17), .A2(n1303), .ZN(n1321) );
XNOR2_X1 U1059 ( .A(n1323), .B(G478), .ZN(n1069) );
NAND2_X1 U1060 ( .A1(n1162), .A2(n1118), .ZN(n1323) );
NAND2_X1 U1061 ( .A1(n1324), .A2(n1325), .ZN(n1118) );
NAND4_X1 U1062 ( .A1(n1326), .A2(G217), .A3(n1327), .A4(n1043), .ZN(n1325) );
XNOR2_X1 U1063 ( .A(n1328), .B(n1329), .ZN(n1326) );
XOR2_X1 U1064 ( .A(n1330), .B(KEYINPUT2), .Z(n1324) );
NAND2_X1 U1065 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND3_X1 U1066 ( .A1(n1327), .A2(n1043), .A3(G217), .ZN(n1332) );
INV_X1 U1067 ( .A(G953), .ZN(n1043) );
XNOR2_X1 U1068 ( .A(n1250), .B(KEYINPUT35), .ZN(n1327) );
INV_X1 U1069 ( .A(G234), .ZN(n1250) );
XNOR2_X1 U1070 ( .A(n1329), .B(n1333), .ZN(n1331) );
INV_X1 U1071 ( .A(n1328), .ZN(n1333) );
XOR2_X1 U1072 ( .A(G122), .B(n1334), .Z(n1328) );
XNOR2_X1 U1073 ( .A(n1303), .B(G128), .ZN(n1334) );
INV_X1 U1074 ( .A(G143), .ZN(n1303) );
XNOR2_X1 U1075 ( .A(n1335), .B(n1336), .ZN(n1329) );
XNOR2_X1 U1076 ( .A(G116), .B(n1337), .ZN(n1336) );
NAND2_X1 U1077 ( .A1(n1338), .A2(n1001), .ZN(n1337) );
INV_X1 U1078 ( .A(G107), .ZN(n1001) );
XNOR2_X1 U1079 ( .A(KEYINPUT63), .B(KEYINPUT19), .ZN(n1338) );
NAND2_X1 U1080 ( .A1(KEYINPUT0), .A2(n1306), .ZN(n1335) );
INV_X1 U1081 ( .A(G134), .ZN(n1306) );
INV_X1 U1082 ( .A(G902), .ZN(n1162) );
endmodule


