//Key = 0011110011110100100010011011001100111111101110001100111110011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258;

XNOR2_X1 U692 ( .A(G107), .B(n952), .ZN(G9) );
NAND2_X1 U693 ( .A1(KEYINPUT39), .A2(n953), .ZN(n952) );
NAND4_X1 U694 ( .A1(n954), .A2(n955), .A3(n956), .A4(n957), .ZN(G75) );
NAND4_X1 U695 ( .A1(n958), .A2(n959), .A3(n960), .A4(n961), .ZN(n956) );
NOR4_X1 U696 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n961) );
XNOR2_X1 U697 ( .A(G472), .B(n966), .ZN(n964) );
NOR2_X1 U698 ( .A1(n967), .A2(KEYINPUT63), .ZN(n966) );
XNOR2_X1 U699 ( .A(n968), .B(n969), .ZN(n963) );
NAND2_X1 U700 ( .A1(KEYINPUT2), .A2(n970), .ZN(n968) );
XNOR2_X1 U701 ( .A(n971), .B(G475), .ZN(n960) );
NAND2_X1 U702 ( .A1(n972), .A2(n973), .ZN(n955) );
NAND2_X1 U703 ( .A1(n974), .A2(n975), .ZN(n973) );
NAND3_X1 U704 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n975) );
NAND2_X1 U705 ( .A1(n979), .A2(n980), .ZN(n977) );
NAND2_X1 U706 ( .A1(n959), .A2(n981), .ZN(n980) );
OR2_X1 U707 ( .A1(n982), .A2(n983), .ZN(n981) );
NAND2_X1 U708 ( .A1(n984), .A2(n985), .ZN(n979) );
NAND2_X1 U709 ( .A1(n986), .A2(n987), .ZN(n985) );
NAND2_X1 U710 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND3_X1 U711 ( .A1(n984), .A2(n990), .A3(n959), .ZN(n974) );
NAND2_X1 U712 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U713 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U714 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U715 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U716 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U717 ( .A1(n976), .A2(n962), .ZN(n995) );
NAND2_X1 U718 ( .A1(n976), .A2(n1001), .ZN(n991) );
INV_X1 U719 ( .A(n1002), .ZN(n972) );
XOR2_X1 U720 ( .A(n1003), .B(n1004), .Z(G72) );
NOR2_X1 U721 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U722 ( .A1(n1007), .A2(n957), .ZN(n1006) );
NOR2_X1 U723 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR2_X1 U724 ( .A1(G227), .A2(n1010), .ZN(n1008) );
NOR2_X1 U725 ( .A1(n1011), .A2(n1012), .ZN(n1005) );
INV_X1 U726 ( .A(n1010), .ZN(n1012) );
XNOR2_X1 U727 ( .A(n1013), .B(KEYINPUT19), .ZN(n1010) );
NAND2_X1 U728 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U729 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U730 ( .A(n1018), .ZN(n1016) );
XOR2_X1 U731 ( .A(n1019), .B(KEYINPUT14), .Z(n1014) );
NAND2_X1 U732 ( .A1(n1020), .A2(n1018), .ZN(n1019) );
XNOR2_X1 U733 ( .A(n1021), .B(n1022), .ZN(n1018) );
XNOR2_X1 U734 ( .A(KEYINPUT36), .B(n1023), .ZN(n1022) );
XNOR2_X1 U735 ( .A(n1024), .B(n1025), .ZN(n1021) );
NOR2_X1 U736 ( .A1(KEYINPUT18), .A2(n1026), .ZN(n1025) );
NOR2_X1 U737 ( .A1(KEYINPUT33), .A2(n1027), .ZN(n1024) );
XNOR2_X1 U738 ( .A(n1028), .B(KEYINPUT5), .ZN(n1027) );
XOR2_X1 U739 ( .A(KEYINPUT3), .B(n1017), .Z(n1020) );
NOR2_X1 U740 ( .A1(G227), .A2(n957), .ZN(n1011) );
NAND2_X1 U741 ( .A1(n957), .A2(n1029), .ZN(n1003) );
XOR2_X1 U742 ( .A(n1030), .B(n1031), .Z(G69) );
XOR2_X1 U743 ( .A(n1032), .B(n1033), .Z(n1031) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U745 ( .A1(n1036), .A2(n957), .ZN(n1032) );
XNOR2_X1 U746 ( .A(KEYINPUT16), .B(n1037), .ZN(n1036) );
NAND2_X1 U747 ( .A1(G953), .A2(n1038), .ZN(n1030) );
NAND2_X1 U748 ( .A1(G898), .A2(G224), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(G66) );
XOR2_X1 U750 ( .A(n1041), .B(n1042), .Z(n1040) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U752 ( .A1(n1039), .A2(n1045), .ZN(G63) );
XOR2_X1 U753 ( .A(n1046), .B(n1047), .Z(n1045) );
NOR2_X1 U754 ( .A1(n970), .A2(n1048), .ZN(n1047) );
INV_X1 U755 ( .A(G478), .ZN(n970) );
NAND2_X1 U756 ( .A1(KEYINPUT23), .A2(n1049), .ZN(n1046) );
XOR2_X1 U757 ( .A(KEYINPUT27), .B(n1050), .Z(n1049) );
NOR2_X1 U758 ( .A1(n1039), .A2(n1051), .ZN(G60) );
NOR3_X1 U759 ( .A1(n971), .A2(n1052), .A3(n1053), .ZN(n1051) );
NOR4_X1 U760 ( .A1(n1054), .A2(n1048), .A3(KEYINPUT62), .A4(n1055), .ZN(n1053) );
INV_X1 U761 ( .A(n1043), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NOR3_X1 U763 ( .A1(n1055), .A2(KEYINPUT62), .A3(n954), .ZN(n1056) );
XOR2_X1 U764 ( .A(n1058), .B(n1059), .Z(G6) );
XOR2_X1 U765 ( .A(KEYINPUT53), .B(G104), .Z(n1059) );
NAND4_X1 U766 ( .A1(n1060), .A2(n984), .A3(n1061), .A4(n1062), .ZN(n1058) );
XOR2_X1 U767 ( .A(KEYINPUT29), .B(n1001), .Z(n1062) );
NOR2_X1 U768 ( .A1(n1039), .A2(n1063), .ZN(G57) );
XNOR2_X1 U769 ( .A(n1064), .B(n1065), .ZN(n1063) );
NAND2_X1 U770 ( .A1(n1043), .A2(G472), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1039), .A2(n1066), .ZN(G54) );
XOR2_X1 U772 ( .A(n1067), .B(n1068), .Z(n1066) );
XNOR2_X1 U773 ( .A(n1069), .B(n1070), .ZN(n1068) );
NAND2_X1 U774 ( .A1(KEYINPUT24), .A2(n1071), .ZN(n1070) );
XOR2_X1 U775 ( .A(n1072), .B(n1073), .Z(n1071) );
NAND2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U778 ( .A(n1078), .ZN(n1077) );
XNOR2_X1 U779 ( .A(n1026), .B(n1079), .ZN(n1076) );
XNOR2_X1 U780 ( .A(KEYINPUT6), .B(KEYINPUT56), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1026), .A2(n1078), .ZN(n1074) );
XNOR2_X1 U782 ( .A(n1080), .B(KEYINPUT50), .ZN(n1078) );
XOR2_X1 U783 ( .A(n1081), .B(n1082), .Z(n1067) );
XOR2_X1 U784 ( .A(KEYINPUT12), .B(n1083), .Z(n1082) );
NOR2_X1 U785 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U786 ( .A(KEYINPUT45), .B(n1086), .Z(n1085) );
NOR2_X1 U787 ( .A1(G140), .A2(n1087), .ZN(n1086) );
XNOR2_X1 U788 ( .A(KEYINPUT40), .B(n1088), .ZN(n1087) );
NAND2_X1 U789 ( .A1(n1043), .A2(n1089), .ZN(n1081) );
XOR2_X1 U790 ( .A(KEYINPUT22), .B(G469), .Z(n1089) );
NOR2_X1 U791 ( .A1(n957), .A2(G952), .ZN(n1039) );
NOR2_X1 U792 ( .A1(n1090), .A2(n1091), .ZN(G51) );
XOR2_X1 U793 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U794 ( .A(n1035), .B(n1094), .Z(n1093) );
XNOR2_X1 U795 ( .A(n1095), .B(KEYINPUT13), .ZN(n1092) );
NAND3_X1 U796 ( .A1(n1043), .A2(G210), .A3(KEYINPUT48), .ZN(n1095) );
NOR2_X1 U797 ( .A1(n1096), .A2(n954), .ZN(n1043) );
NOR2_X1 U798 ( .A1(n1037), .A2(n1029), .ZN(n954) );
NAND2_X1 U799 ( .A1(n1097), .A2(n1098), .ZN(n1029) );
NOR4_X1 U800 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1098) );
NOR4_X1 U801 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1097) );
INV_X1 U802 ( .A(n1107), .ZN(n1106) );
NAND2_X1 U803 ( .A1(n1108), .A2(n1109), .ZN(n1037) );
NOR4_X1 U804 ( .A1(n1110), .A2(n953), .A3(n1111), .A4(n1112), .ZN(n1109) );
INV_X1 U805 ( .A(n1113), .ZN(n1112) );
INV_X1 U806 ( .A(n1114), .ZN(n1111) );
NOR3_X1 U807 ( .A1(n1115), .A2(n1116), .A3(n1000), .ZN(n953) );
INV_X1 U808 ( .A(n1117), .ZN(n1000) );
NOR4_X1 U809 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1108) );
NOR3_X1 U810 ( .A1(n999), .A2(n1116), .A3(n1115), .ZN(n1121) );
INV_X1 U811 ( .A(n984), .ZN(n1115) );
INV_X1 U812 ( .A(n1060), .ZN(n999) );
NOR2_X1 U813 ( .A1(n1122), .A2(n957), .ZN(n1090) );
XNOR2_X1 U814 ( .A(G952), .B(KEYINPUT34), .ZN(n1122) );
XOR2_X1 U815 ( .A(G146), .B(n1104), .Z(G48) );
AND3_X1 U816 ( .A1(n1060), .A2(n1123), .A3(n1124), .ZN(n1104) );
XNOR2_X1 U817 ( .A(G143), .B(n1107), .ZN(G45) );
NAND4_X1 U818 ( .A1(n1001), .A2(n1123), .A3(n983), .A4(n1125), .ZN(n1107) );
NOR3_X1 U819 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
XNOR2_X1 U820 ( .A(n1129), .B(n1103), .ZN(G42) );
AND3_X1 U821 ( .A1(n1060), .A2(n982), .A3(n1130), .ZN(n1103) );
NAND2_X1 U822 ( .A1(n1131), .A2(n1132), .ZN(G39) );
NAND2_X1 U823 ( .A1(n1105), .A2(n1133), .ZN(n1132) );
INV_X1 U824 ( .A(n1134), .ZN(n1105) );
XOR2_X1 U825 ( .A(n1135), .B(KEYINPUT41), .Z(n1131) );
NAND2_X1 U826 ( .A1(G137), .A2(n1134), .ZN(n1135) );
NAND3_X1 U827 ( .A1(n976), .A2(n959), .A3(n1124), .ZN(n1134) );
XOR2_X1 U828 ( .A(G134), .B(n1102), .Z(G36) );
AND3_X1 U829 ( .A1(n983), .A2(n1117), .A3(n1130), .ZN(n1102) );
XOR2_X1 U830 ( .A(n1136), .B(n1101), .Z(G33) );
AND3_X1 U831 ( .A1(n1060), .A2(n983), .A3(n1130), .ZN(n1101) );
AND3_X1 U832 ( .A1(n1001), .A2(n1137), .A3(n959), .ZN(n1130) );
NOR2_X1 U833 ( .A1(n1138), .A2(n988), .ZN(n959) );
XNOR2_X1 U834 ( .A(G131), .B(KEYINPUT55), .ZN(n1136) );
XNOR2_X1 U835 ( .A(n1139), .B(n1100), .ZN(G30) );
AND3_X1 U836 ( .A1(n1117), .A2(n1123), .A3(n1124), .ZN(n1100) );
AND4_X1 U837 ( .A1(n1140), .A2(n1001), .A3(n965), .A4(n1137), .ZN(n1124) );
XOR2_X1 U838 ( .A(n1110), .B(n1141), .Z(G3) );
NOR2_X1 U839 ( .A1(KEYINPUT0), .A2(n1142), .ZN(n1141) );
AND3_X1 U840 ( .A1(n983), .A2(n1143), .A3(n976), .ZN(n1110) );
XOR2_X1 U841 ( .A(G125), .B(n1099), .Z(G27) );
AND4_X1 U842 ( .A1(n1060), .A2(n978), .A3(n1144), .A4(n982), .ZN(n1099) );
NOR2_X1 U843 ( .A1(n1126), .A2(n986), .ZN(n1144) );
INV_X1 U844 ( .A(n1123), .ZN(n986) );
INV_X1 U845 ( .A(n1137), .ZN(n1126) );
NAND2_X1 U846 ( .A1(n1002), .A2(n1145), .ZN(n1137) );
NAND4_X1 U847 ( .A1(G953), .A2(G902), .A3(n1146), .A4(n1009), .ZN(n1145) );
INV_X1 U848 ( .A(G900), .ZN(n1009) );
XOR2_X1 U849 ( .A(G122), .B(n1120), .Z(G24) );
AND4_X1 U850 ( .A1(n1147), .A2(n984), .A3(n1148), .A4(n1149), .ZN(n1120) );
NOR2_X1 U851 ( .A1(n965), .A2(n1140), .ZN(n984) );
XOR2_X1 U852 ( .A(G119), .B(n1119), .Z(G21) );
AND4_X1 U853 ( .A1(n1147), .A2(n976), .A3(n1140), .A4(n965), .ZN(n1119) );
XNOR2_X1 U854 ( .A(n1150), .B(n1118), .ZN(G18) );
AND3_X1 U855 ( .A1(n983), .A2(n1117), .A3(n1147), .ZN(n1118) );
NOR2_X1 U856 ( .A1(n1148), .A2(n1127), .ZN(n1117) );
INV_X1 U857 ( .A(n1149), .ZN(n1127) );
XNOR2_X1 U858 ( .A(G113), .B(n1113), .ZN(G15) );
NAND3_X1 U859 ( .A1(n1147), .A2(n983), .A3(n1060), .ZN(n1113) );
NOR2_X1 U860 ( .A1(n1149), .A2(n1128), .ZN(n1060) );
INV_X1 U861 ( .A(n1148), .ZN(n1128) );
NOR2_X1 U862 ( .A1(n1151), .A2(n965), .ZN(n983) );
AND2_X1 U863 ( .A1(n978), .A2(n1061), .ZN(n1147) );
AND2_X1 U864 ( .A1(n997), .A2(n993), .ZN(n978) );
INV_X1 U865 ( .A(n1152), .ZN(n997) );
XNOR2_X1 U866 ( .A(G110), .B(n1114), .ZN(G12) );
NAND3_X1 U867 ( .A1(n976), .A2(n1143), .A3(n982), .ZN(n1114) );
AND2_X1 U868 ( .A1(n1153), .A2(n965), .ZN(n982) );
XNOR2_X1 U869 ( .A(n1154), .B(n1044), .ZN(n965) );
AND2_X1 U870 ( .A1(G217), .A2(n1155), .ZN(n1044) );
NAND2_X1 U871 ( .A1(n1156), .A2(n1041), .ZN(n1154) );
NAND2_X1 U872 ( .A1(n1157), .A2(n1158), .ZN(n1041) );
NAND2_X1 U873 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U874 ( .A(KEYINPUT11), .B(n1161), .Z(n1157) );
NOR2_X1 U875 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
XNOR2_X1 U876 ( .A(n1162), .B(G137), .ZN(n1160) );
NAND2_X1 U877 ( .A1(G221), .A2(n1163), .ZN(n1162) );
XOR2_X1 U878 ( .A(n1164), .B(n1165), .Z(n1159) );
NOR2_X1 U879 ( .A1(KEYINPUT57), .A2(n1166), .ZN(n1165) );
XOR2_X1 U880 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U881 ( .A(G119), .B(G110), .ZN(n1168) );
NAND2_X1 U882 ( .A1(KEYINPUT9), .A2(n1139), .ZN(n1167) );
XNOR2_X1 U883 ( .A(G902), .B(KEYINPUT47), .ZN(n1156) );
XNOR2_X1 U884 ( .A(KEYINPUT1), .B(n1140), .ZN(n1153) );
INV_X1 U885 ( .A(n1151), .ZN(n1140) );
XOR2_X1 U886 ( .A(n967), .B(n1169), .Z(n1151) );
NOR2_X1 U887 ( .A1(G472), .A2(KEYINPUT28), .ZN(n1169) );
AND2_X1 U888 ( .A1(n1170), .A2(n1096), .ZN(n967) );
XNOR2_X1 U889 ( .A(KEYINPUT43), .B(n1171), .ZN(n1170) );
INV_X1 U890 ( .A(n1065), .ZN(n1171) );
XNOR2_X1 U891 ( .A(n1172), .B(n1173), .ZN(n1065) );
XOR2_X1 U892 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U893 ( .A(n1176), .B(n1142), .ZN(n1175) );
NAND2_X1 U894 ( .A1(G210), .A2(n1177), .ZN(n1176) );
XNOR2_X1 U895 ( .A(G113), .B(KEYINPUT32), .ZN(n1174) );
XOR2_X1 U896 ( .A(n1178), .B(n1179), .Z(n1172) );
XOR2_X1 U897 ( .A(n1180), .B(n1181), .Z(n1178) );
INV_X1 U898 ( .A(n1116), .ZN(n1143) );
NAND2_X1 U899 ( .A1(n1001), .A2(n1061), .ZN(n1116) );
AND2_X1 U900 ( .A1(n1123), .A2(n1182), .ZN(n1061) );
NAND2_X1 U901 ( .A1(n1002), .A2(n1183), .ZN(n1182) );
NAND3_X1 U902 ( .A1(G902), .A2(n1146), .A3(n1034), .ZN(n1183) );
NOR2_X1 U903 ( .A1(n957), .A2(G898), .ZN(n1034) );
NAND3_X1 U904 ( .A1(n1146), .A2(n957), .A3(G952), .ZN(n1002) );
NAND2_X1 U905 ( .A1(G237), .A2(G234), .ZN(n1146) );
NOR2_X1 U906 ( .A1(n989), .A2(n988), .ZN(n1123) );
AND2_X1 U907 ( .A1(G214), .A2(n1184), .ZN(n988) );
INV_X1 U908 ( .A(n1138), .ZN(n989) );
XNOR2_X1 U909 ( .A(n1185), .B(n1186), .ZN(n1138) );
AND2_X1 U910 ( .A1(n1184), .A2(G210), .ZN(n1186) );
OR2_X1 U911 ( .A1(G902), .A2(G237), .ZN(n1184) );
NAND2_X1 U912 ( .A1(n1187), .A2(n1096), .ZN(n1185) );
XNOR2_X1 U913 ( .A(n1188), .B(n1035), .ZN(n1187) );
XOR2_X1 U914 ( .A(n1189), .B(n1190), .Z(n1035) );
XNOR2_X1 U915 ( .A(n1142), .B(n1191), .ZN(n1190) );
XNOR2_X1 U916 ( .A(G122), .B(n1088), .ZN(n1191) );
XOR2_X1 U917 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR2_X1 U918 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U919 ( .A(n1196), .B(KEYINPUT61), .Z(n1195) );
NAND2_X1 U920 ( .A1(n1197), .A2(G113), .ZN(n1196) );
NOR2_X1 U921 ( .A1(G113), .A2(n1197), .ZN(n1194) );
XNOR2_X1 U922 ( .A(KEYINPUT31), .B(n1181), .ZN(n1197) );
XNOR2_X1 U923 ( .A(n1150), .B(G119), .ZN(n1181) );
INV_X1 U924 ( .A(G116), .ZN(n1150) );
NAND3_X1 U925 ( .A1(n1198), .A2(n1199), .A3(KEYINPUT38), .ZN(n1192) );
NAND2_X1 U926 ( .A1(G104), .A2(n1200), .ZN(n1198) );
NOR2_X1 U927 ( .A1(KEYINPUT17), .A2(n1094), .ZN(n1188) );
XOR2_X1 U928 ( .A(n1180), .B(n1201), .Z(n1094) );
XOR2_X1 U929 ( .A(G125), .B(n1202), .Z(n1201) );
AND2_X1 U930 ( .A1(n957), .A2(G224), .ZN(n1202) );
XNOR2_X1 U931 ( .A(n1203), .B(n1139), .ZN(n1180) );
INV_X1 U932 ( .A(G128), .ZN(n1139) );
NAND2_X1 U933 ( .A1(KEYINPUT44), .A2(n1204), .ZN(n1203) );
XOR2_X1 U934 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U935 ( .A(KEYINPUT51), .B(G146), .Z(n1206) );
NOR2_X1 U936 ( .A1(KEYINPUT21), .A2(n1207), .ZN(n1205) );
XNOR2_X1 U937 ( .A(G143), .B(KEYINPUT4), .ZN(n1207) );
NOR2_X1 U938 ( .A1(n993), .A2(n1152), .ZN(n1001) );
XNOR2_X1 U939 ( .A(n962), .B(KEYINPUT52), .ZN(n1152) );
AND2_X1 U940 ( .A1(G221), .A2(n1155), .ZN(n962) );
NAND2_X1 U941 ( .A1(G234), .A2(n1096), .ZN(n1155) );
XNOR2_X1 U942 ( .A(n958), .B(KEYINPUT37), .ZN(n993) );
XOR2_X1 U943 ( .A(n1208), .B(G469), .Z(n958) );
NAND2_X1 U944 ( .A1(n1209), .A2(n1096), .ZN(n1208) );
INV_X1 U945 ( .A(G902), .ZN(n1096) );
XOR2_X1 U946 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U947 ( .A(n1212), .B(n1213), .Z(n1211) );
NAND2_X1 U948 ( .A1(KEYINPUT35), .A2(n1069), .ZN(n1213) );
AND2_X1 U949 ( .A1(G227), .A2(n957), .ZN(n1069) );
NAND3_X1 U950 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1212) );
NAND2_X1 U951 ( .A1(n1084), .A2(n1080), .ZN(n1216) );
NOR2_X1 U952 ( .A1(n1129), .A2(G110), .ZN(n1084) );
OR3_X1 U953 ( .A1(n1080), .A2(n1088), .A3(n1129), .ZN(n1215) );
INV_X1 U954 ( .A(G110), .ZN(n1088) );
NAND2_X1 U955 ( .A1(n1217), .A2(n1129), .ZN(n1214) );
XNOR2_X1 U956 ( .A(G110), .B(n1080), .ZN(n1217) );
NAND2_X1 U957 ( .A1(n1218), .A2(n1219), .ZN(n1080) );
NAND3_X1 U958 ( .A1(n1220), .A2(n1199), .A3(n1221), .ZN(n1219) );
XOR2_X1 U959 ( .A(KEYINPUT20), .B(n1222), .Z(n1218) );
NOR2_X1 U960 ( .A1(n1223), .A2(n1221), .ZN(n1222) );
XNOR2_X1 U961 ( .A(n1142), .B(KEYINPUT60), .ZN(n1221) );
INV_X1 U962 ( .A(G101), .ZN(n1142) );
AND2_X1 U963 ( .A1(n1199), .A2(n1220), .ZN(n1223) );
XNOR2_X1 U964 ( .A(n1224), .B(KEYINPUT30), .ZN(n1220) );
NAND2_X1 U965 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U966 ( .A(KEYINPUT25), .B(G104), .Z(n1226) );
XNOR2_X1 U967 ( .A(KEYINPUT59), .B(n1200), .ZN(n1225) );
OR2_X1 U968 ( .A1(n1200), .A2(G104), .ZN(n1199) );
XNOR2_X1 U969 ( .A(n1073), .B(n1026), .ZN(n1210) );
XOR2_X1 U970 ( .A(G128), .B(n1227), .Z(n1026) );
NOR2_X1 U971 ( .A1(KEYINPUT15), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U972 ( .A(G146), .B(n1229), .ZN(n1228) );
XOR2_X1 U973 ( .A(n1179), .B(KEYINPUT42), .Z(n1073) );
XOR2_X1 U974 ( .A(G131), .B(n1028), .Z(n1179) );
XNOR2_X1 U975 ( .A(G134), .B(n1133), .ZN(n1028) );
INV_X1 U976 ( .A(G137), .ZN(n1133) );
NOR2_X1 U977 ( .A1(n1149), .A2(n1148), .ZN(n976) );
NAND2_X1 U978 ( .A1(n1230), .A2(n1231), .ZN(n1148) );
NAND2_X1 U979 ( .A1(n1232), .A2(n1055), .ZN(n1231) );
XOR2_X1 U980 ( .A(KEYINPUT8), .B(n1233), .Z(n1230) );
NOR2_X1 U981 ( .A1(n1232), .A2(n1055), .ZN(n1233) );
INV_X1 U982 ( .A(G475), .ZN(n1055) );
XNOR2_X1 U983 ( .A(n971), .B(KEYINPUT49), .ZN(n1232) );
NOR2_X1 U984 ( .A1(n1057), .A2(G902), .ZN(n971) );
INV_X1 U985 ( .A(n1054), .ZN(n1057) );
XNOR2_X1 U986 ( .A(n1234), .B(n1235), .ZN(n1054) );
XOR2_X1 U987 ( .A(G104), .B(n1236), .Z(n1235) );
NOR2_X1 U988 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U989 ( .A(n1239), .B(KEYINPUT26), .Z(n1238) );
NAND2_X1 U990 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U991 ( .A1(n1241), .A2(n1240), .ZN(n1237) );
XOR2_X1 U992 ( .A(KEYINPUT46), .B(G122), .Z(n1240) );
INV_X1 U993 ( .A(G113), .ZN(n1241) );
XOR2_X1 U994 ( .A(n1164), .B(n1242), .Z(n1234) );
NOR2_X1 U995 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U996 ( .A(n1245), .B(KEYINPUT10), .Z(n1244) );
NAND2_X1 U997 ( .A1(n1246), .A2(n1023), .ZN(n1245) );
NOR2_X1 U998 ( .A1(n1246), .A2(n1023), .ZN(n1243) );
INV_X1 U999 ( .A(G131), .ZN(n1023) );
XNOR2_X1 U1000 ( .A(n1247), .B(G143), .ZN(n1246) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1177), .ZN(n1247) );
NOR2_X1 U1002 ( .A1(G953), .A2(G237), .ZN(n1177) );
XNOR2_X1 U1003 ( .A(G146), .B(n1017), .ZN(n1164) );
XNOR2_X1 U1004 ( .A(G125), .B(n1129), .ZN(n1017) );
INV_X1 U1005 ( .A(G140), .ZN(n1129) );
NAND2_X1 U1006 ( .A1(n1248), .A2(n1249), .ZN(n1149) );
NAND2_X1 U1007 ( .A1(G478), .A2(n969), .ZN(n1249) );
XOR2_X1 U1008 ( .A(KEYINPUT54), .B(n1250), .Z(n1248) );
NOR2_X1 U1009 ( .A1(G478), .A2(n969), .ZN(n1250) );
OR2_X1 U1010 ( .A1(n1050), .A2(G902), .ZN(n969) );
XNOR2_X1 U1011 ( .A(n1251), .B(n1252), .ZN(n1050) );
XOR2_X1 U1012 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U1013 ( .A(n1200), .B(n1255), .ZN(n1254) );
NOR2_X1 U1014 ( .A1(KEYINPUT7), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U1015 ( .A(n1229), .B(G128), .ZN(n1256) );
INV_X1 U1016 ( .A(G143), .ZN(n1229) );
INV_X1 U1017 ( .A(G107), .ZN(n1200) );
AND2_X1 U1018 ( .A1(n1163), .A2(G217), .ZN(n1253) );
AND2_X1 U1019 ( .A1(G234), .A2(n957), .ZN(n1163) );
INV_X1 U1020 ( .A(G953), .ZN(n957) );
XOR2_X1 U1021 ( .A(n1257), .B(n1258), .Z(n1251) );
XOR2_X1 U1022 ( .A(KEYINPUT58), .B(G134), .Z(n1258) );
XNOR2_X1 U1023 ( .A(G116), .B(G122), .ZN(n1257) );
endmodule


