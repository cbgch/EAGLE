//Key = 1001110000100001010101011110100001000110110111101111111011011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289;

XOR2_X1 U715 ( .A(n990), .B(n991), .Z(G9) );
XOR2_X1 U716 ( .A(KEYINPUT43), .B(G107), .Z(n991) );
NAND4_X1 U717 ( .A1(KEYINPUT37), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
NOR2_X1 U718 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U719 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n996) );
INV_X1 U720 ( .A(G952), .ZN(n1000) );
NOR2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND4_X1 U722 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n997) );
NAND3_X1 U723 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
XNOR2_X1 U724 ( .A(KEYINPUT6), .B(n1002), .ZN(n1008) );
NAND4_X1 U725 ( .A1(n1010), .A2(n1011), .A3(n994), .A4(n1012), .ZN(n1002) );
NAND3_X1 U726 ( .A1(n1013), .A2(n1014), .A3(n1010), .ZN(n1003) );
INV_X1 U727 ( .A(n1015), .ZN(n1010) );
NAND2_X1 U728 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND3_X1 U729 ( .A1(n1012), .A2(n1018), .A3(n994), .ZN(n1017) );
NAND2_X1 U730 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
INV_X1 U732 ( .A(n1023), .ZN(n1019) );
NAND2_X1 U733 ( .A1(n1011), .A2(n1024), .ZN(n1016) );
NAND2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U735 ( .A1(n994), .A2(n1027), .ZN(n1026) );
NAND2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U737 ( .A1(n1012), .A2(n1030), .ZN(n1025) );
NAND2_X1 U738 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
INV_X1 U740 ( .A(n1035), .ZN(n1031) );
NOR3_X1 U741 ( .A1(n1036), .A2(G953), .A3(n1037), .ZN(n995) );
INV_X1 U742 ( .A(n1005), .ZN(n1037) );
NAND2_X1 U743 ( .A1(n1038), .A2(n1039), .ZN(n1005) );
NOR4_X1 U744 ( .A1(n1009), .A2(n1021), .A3(n1040), .A4(n1041), .ZN(n1039) );
XNOR2_X1 U745 ( .A(G469), .B(n1042), .ZN(n1041) );
NOR2_X1 U746 ( .A1(n1043), .A2(KEYINPUT22), .ZN(n1042) );
XOR2_X1 U747 ( .A(n1044), .B(n1045), .Z(n1040) );
NAND2_X1 U748 ( .A1(KEYINPUT26), .A2(n1046), .ZN(n1044) );
NOR4_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1038) );
XOR2_X1 U750 ( .A(n1051), .B(n1052), .Z(n1047) );
XOR2_X1 U751 ( .A(KEYINPUT46), .B(n1053), .Z(n1052) );
XNOR2_X1 U752 ( .A(G952), .B(KEYINPUT40), .ZN(n1036) );
XOR2_X1 U753 ( .A(n1054), .B(n1055), .Z(G72) );
XOR2_X1 U754 ( .A(n1056), .B(n1057), .Z(n1055) );
NOR2_X1 U755 ( .A1(G953), .A2(n1058), .ZN(n1057) );
NOR2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XNOR2_X1 U757 ( .A(KEYINPUT47), .B(n1061), .ZN(n1060) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
NAND2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U760 ( .A(G900), .ZN(n1065) );
XNOR2_X1 U761 ( .A(G953), .B(KEYINPUT23), .ZN(n1064) );
XOR2_X1 U762 ( .A(n1066), .B(n1067), .Z(n1062) );
XNOR2_X1 U763 ( .A(n1068), .B(n1069), .ZN(n1067) );
XOR2_X1 U764 ( .A(n1070), .B(n1071), .Z(n1066) );
XNOR2_X1 U765 ( .A(KEYINPUT41), .B(KEYINPUT18), .ZN(n1071) );
NAND2_X1 U766 ( .A1(KEYINPUT15), .A2(n1072), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1073), .B(n1074), .Z(n1072) );
XNOR2_X1 U768 ( .A(G137), .B(n1075), .ZN(n1074) );
NOR2_X1 U769 ( .A1(G134), .A2(KEYINPUT35), .ZN(n1073) );
NAND2_X1 U770 ( .A1(G953), .A2(n1076), .ZN(n1054) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1076) );
XOR2_X1 U772 ( .A(n1077), .B(n1078), .Z(G69) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1006), .A2(n1081), .ZN(n1080) );
XOR2_X1 U775 ( .A(KEYINPUT13), .B(n1082), .Z(n1081) );
AND2_X1 U776 ( .A1(G224), .A2(G898), .ZN(n1082) );
NOR2_X1 U777 ( .A1(G953), .A2(n1083), .ZN(n1079) );
NAND4_X1 U778 ( .A1(n1084), .A2(KEYINPUT17), .A3(n1085), .A4(n1086), .ZN(n1077) );
NAND2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U780 ( .A1(G953), .A2(n1089), .ZN(n1085) );
XOR2_X1 U781 ( .A(n1090), .B(KEYINPUT27), .Z(n1084) );
OR2_X1 U782 ( .A1(n1088), .A2(n1087), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1091), .B(n1092), .Z(n1087) );
NAND2_X1 U784 ( .A1(KEYINPUT52), .A2(n1093), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(G66) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U788 ( .A1(KEYINPUT9), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U789 ( .A(n1101), .B(KEYINPUT39), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
XOR2_X1 U791 ( .A(KEYINPUT56), .B(n1053), .Z(n1103) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1096) );
XNOR2_X1 U793 ( .A(KEYINPUT39), .B(n1106), .ZN(n1105) );
INV_X1 U794 ( .A(n1101), .ZN(n1106) );
INV_X1 U795 ( .A(KEYINPUT9), .ZN(n1104) );
NOR2_X1 U796 ( .A1(n1094), .A2(n1107), .ZN(G63) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1110), .B(KEYINPUT51), .Z(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U800 ( .A(n1113), .B(KEYINPUT7), .ZN(n1111) );
NOR2_X1 U801 ( .A1(n1112), .A2(n1114), .ZN(n1108) );
INV_X1 U802 ( .A(n1113), .ZN(n1114) );
AND2_X1 U803 ( .A1(n1115), .A2(G478), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1094), .A2(n1116), .ZN(G60) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U806 ( .A1(n1115), .A2(G475), .ZN(n1118) );
NAND2_X1 U807 ( .A1(KEYINPUT54), .A2(n1119), .ZN(n1117) );
XOR2_X1 U808 ( .A(KEYINPUT55), .B(n1120), .Z(n1119) );
XNOR2_X1 U809 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1094), .A2(n1122), .ZN(G57) );
XOR2_X1 U811 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U812 ( .A1(n1046), .A2(n1102), .ZN(n1124) );
NOR2_X1 U813 ( .A1(n1094), .A2(n1125), .ZN(G54) );
XOR2_X1 U814 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U815 ( .A(n1128), .B(n1129), .ZN(n1127) );
XNOR2_X1 U816 ( .A(n1130), .B(n1131), .ZN(n1126) );
NAND3_X1 U817 ( .A1(n1115), .A2(G469), .A3(KEYINPUT19), .ZN(n1130) );
INV_X1 U818 ( .A(n1102), .ZN(n1115) );
NOR2_X1 U819 ( .A1(n1094), .A2(n1132), .ZN(G51) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U821 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U822 ( .A1(n1137), .A2(n1102), .ZN(n1136) );
NAND2_X1 U823 ( .A1(G902), .A2(n998), .ZN(n1102) );
NAND3_X1 U824 ( .A1(n1083), .A2(n1061), .A3(n1138), .ZN(n998) );
INV_X1 U825 ( .A(n1059), .ZN(n1138) );
NAND4_X1 U826 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1059) );
AND3_X1 U827 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NAND2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NAND2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
OR2_X1 U830 ( .A1(n1028), .A2(KEYINPUT8), .ZN(n1149) );
XNOR2_X1 U831 ( .A(KEYINPUT59), .B(n1029), .ZN(n1148) );
NAND2_X1 U832 ( .A1(n1150), .A2(n1151), .ZN(n1139) );
NAND2_X1 U833 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND3_X1 U834 ( .A1(n1154), .A2(n1001), .A3(KEYINPUT8), .ZN(n1153) );
INV_X1 U835 ( .A(n1155), .ZN(n1001) );
NAND2_X1 U836 ( .A1(n1013), .A2(n1156), .ZN(n1152) );
AND2_X1 U837 ( .A1(n1157), .A2(n1158), .ZN(n1083) );
AND4_X1 U838 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
AND4_X1 U839 ( .A1(n1163), .A2(n1164), .A3(n1121), .A4(n1165), .ZN(n1157) );
NAND3_X1 U840 ( .A1(n992), .A2(n994), .A3(n993), .ZN(n1165) );
NAND3_X1 U841 ( .A1(n992), .A2(n994), .A3(n1150), .ZN(n1121) );
NAND2_X1 U842 ( .A1(KEYINPUT45), .A2(n1166), .ZN(n1135) );
XOR2_X1 U843 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U844 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
AND3_X1 U846 ( .A1(n1171), .A2(n1173), .A3(G125), .ZN(n1169) );
INV_X1 U847 ( .A(KEYINPUT21), .ZN(n1171) );
NAND2_X1 U848 ( .A1(KEYINPUT33), .A2(n1174), .ZN(n1167) );
NOR2_X1 U849 ( .A1(n1006), .A2(G952), .ZN(n1094) );
XOR2_X1 U850 ( .A(n1175), .B(n1176), .Z(G48) );
XNOR2_X1 U851 ( .A(G146), .B(KEYINPUT30), .ZN(n1176) );
NAND2_X1 U852 ( .A1(n1146), .A2(n1150), .ZN(n1175) );
XNOR2_X1 U853 ( .A(G143), .B(n1140), .ZN(G45) );
NAND4_X1 U854 ( .A1(n1156), .A2(n1155), .A3(n1177), .A4(n1049), .ZN(n1140) );
XNOR2_X1 U855 ( .A(G140), .B(n1143), .ZN(G42) );
NAND3_X1 U856 ( .A1(n1178), .A2(n1179), .A3(n1013), .ZN(n1143) );
NAND2_X1 U857 ( .A1(n1180), .A2(n1181), .ZN(G39) );
NAND2_X1 U858 ( .A1(G137), .A2(n1145), .ZN(n1181) );
XOR2_X1 U859 ( .A(KEYINPUT4), .B(n1182), .Z(n1180) );
NOR2_X1 U860 ( .A1(G137), .A2(n1145), .ZN(n1182) );
NAND3_X1 U861 ( .A1(n1013), .A2(n1012), .A3(n1154), .ZN(n1145) );
XNOR2_X1 U862 ( .A(G134), .B(n1144), .ZN(G36) );
NAND3_X1 U863 ( .A1(n1156), .A2(n993), .A3(n1013), .ZN(n1144) );
NAND2_X1 U864 ( .A1(n1183), .A2(n1184), .ZN(G33) );
NAND2_X1 U865 ( .A1(n1185), .A2(n1075), .ZN(n1184) );
XOR2_X1 U866 ( .A(KEYINPUT60), .B(n1186), .Z(n1183) );
NOR2_X1 U867 ( .A1(n1185), .A2(n1075), .ZN(n1186) );
AND3_X1 U868 ( .A1(n1150), .A2(n1187), .A3(n1156), .ZN(n1185) );
AND3_X1 U869 ( .A1(n1023), .A2(n1188), .A3(n1035), .ZN(n1156) );
XOR2_X1 U870 ( .A(KEYINPUT20), .B(n1013), .Z(n1187) );
NOR2_X1 U871 ( .A1(n1189), .A2(n1009), .ZN(n1013) );
XNOR2_X1 U872 ( .A(G128), .B(n1190), .ZN(G30) );
NAND2_X1 U873 ( .A1(n1146), .A2(n993), .ZN(n1190) );
AND2_X1 U874 ( .A1(n1154), .A2(n1155), .ZN(n1146) );
AND4_X1 U875 ( .A1(n1033), .A2(n1023), .A3(n1191), .A4(n1188), .ZN(n1154) );
XNOR2_X1 U876 ( .A(G101), .B(n1164), .ZN(G3) );
NAND3_X1 U877 ( .A1(n992), .A2(n1012), .A3(n1035), .ZN(n1164) );
XOR2_X1 U878 ( .A(G125), .B(n1192), .Z(G27) );
NOR2_X1 U879 ( .A1(KEYINPUT16), .A2(n1061), .ZN(n1192) );
NAND3_X1 U880 ( .A1(n1022), .A2(n1155), .A3(n1178), .ZN(n1061) );
AND3_X1 U881 ( .A1(n1033), .A2(n1150), .A3(n1193), .ZN(n1178) );
AND3_X1 U882 ( .A1(n1034), .A2(n1194), .A3(n1188), .ZN(n1193) );
NAND2_X1 U883 ( .A1(n1015), .A2(n1195), .ZN(n1188) );
NAND4_X1 U884 ( .A1(n1196), .A2(G953), .A3(G902), .A4(n1197), .ZN(n1195) );
XNOR2_X1 U885 ( .A(G900), .B(KEYINPUT58), .ZN(n1196) );
XNOR2_X1 U886 ( .A(G122), .B(n1163), .ZN(G24) );
NAND4_X1 U887 ( .A1(n1198), .A2(n994), .A3(n1177), .A4(n1049), .ZN(n1163) );
NOR2_X1 U888 ( .A1(n1191), .A2(n1033), .ZN(n994) );
XNOR2_X1 U889 ( .A(G119), .B(n1162), .ZN(G21) );
NAND4_X1 U890 ( .A1(n1033), .A2(n1198), .A3(n1012), .A4(n1191), .ZN(n1162) );
XNOR2_X1 U891 ( .A(G116), .B(n1161), .ZN(G18) );
NAND3_X1 U892 ( .A1(n1035), .A2(n993), .A3(n1198), .ZN(n1161) );
INV_X1 U893 ( .A(n1029), .ZN(n993) );
NAND2_X1 U894 ( .A1(n1199), .A2(n1049), .ZN(n1029) );
XNOR2_X1 U895 ( .A(KEYINPUT0), .B(n1200), .ZN(n1199) );
XOR2_X1 U896 ( .A(G113), .B(n1201), .Z(G15) );
NOR2_X1 U897 ( .A1(KEYINPUT63), .A2(n1160), .ZN(n1201) );
NAND3_X1 U898 ( .A1(n1035), .A2(n1150), .A3(n1198), .ZN(n1160) );
AND2_X1 U899 ( .A1(n1011), .A2(n1202), .ZN(n1198) );
NOR2_X1 U900 ( .A1(n1179), .A2(n1021), .ZN(n1011) );
INV_X1 U901 ( .A(n1022), .ZN(n1179) );
NOR2_X1 U902 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
XNOR2_X1 U903 ( .A(G110), .B(n1159), .ZN(G12) );
NAND4_X1 U904 ( .A1(n1033), .A2(n992), .A3(n1034), .A4(n1012), .ZN(n1159) );
NAND2_X1 U905 ( .A1(n1203), .A2(n1204), .ZN(n1012) );
OR2_X1 U906 ( .A1(n1028), .A2(KEYINPUT0), .ZN(n1204) );
INV_X1 U907 ( .A(n1150), .ZN(n1028) );
NOR2_X1 U908 ( .A1(n1049), .A2(n1200), .ZN(n1150) );
NAND3_X1 U909 ( .A1(n1200), .A2(n1205), .A3(KEYINPUT0), .ZN(n1203) );
INV_X1 U910 ( .A(n1049), .ZN(n1205) );
XNOR2_X1 U911 ( .A(n1206), .B(G478), .ZN(n1049) );
NAND2_X1 U912 ( .A1(n1113), .A2(n1207), .ZN(n1206) );
XNOR2_X1 U913 ( .A(n1208), .B(n1209), .ZN(n1113) );
XOR2_X1 U914 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND3_X1 U915 ( .A1(G234), .A2(n1006), .A3(G217), .ZN(n1211) );
NAND2_X1 U916 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
INV_X1 U917 ( .A(G134), .ZN(n1213) );
XNOR2_X1 U918 ( .A(KEYINPUT31), .B(KEYINPUT29), .ZN(n1212) );
XOR2_X1 U919 ( .A(n1214), .B(n1215), .Z(n1208) );
NOR2_X1 U920 ( .A1(KEYINPUT61), .A2(n1216), .ZN(n1215) );
XOR2_X1 U921 ( .A(n1217), .B(G107), .Z(n1216) );
NAND2_X1 U922 ( .A1(n1218), .A2(KEYINPUT24), .ZN(n1217) );
XNOR2_X1 U923 ( .A(G116), .B(G122), .ZN(n1218) );
XNOR2_X1 U924 ( .A(G143), .B(n1219), .ZN(n1214) );
NOR2_X1 U925 ( .A1(KEYINPUT2), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U926 ( .A(KEYINPUT38), .B(n1221), .ZN(n1220) );
INV_X1 U927 ( .A(n1177), .ZN(n1200) );
XOR2_X1 U928 ( .A(n1050), .B(KEYINPUT32), .Z(n1177) );
XNOR2_X1 U929 ( .A(n1222), .B(G475), .ZN(n1050) );
OR2_X1 U930 ( .A1(n1120), .A2(G902), .ZN(n1222) );
XNOR2_X1 U931 ( .A(n1223), .B(n1224), .ZN(n1120) );
XOR2_X1 U932 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U933 ( .A(KEYINPUT57), .B(G143), .Z(n1226) );
NOR2_X1 U934 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
XOR2_X1 U935 ( .A(n1229), .B(KEYINPUT62), .Z(n1228) );
NAND2_X1 U936 ( .A1(n1230), .A2(G104), .ZN(n1229) );
NOR2_X1 U937 ( .A1(G104), .A2(n1230), .ZN(n1227) );
XOR2_X1 U938 ( .A(n1231), .B(G113), .Z(n1230) );
NAND2_X1 U939 ( .A1(KEYINPUT28), .A2(n1232), .ZN(n1231) );
XOR2_X1 U940 ( .A(n1068), .B(n1233), .Z(n1223) );
XOR2_X1 U941 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR2_X1 U942 ( .A1(G131), .A2(KEYINPUT1), .ZN(n1235) );
AND2_X1 U943 ( .A1(G214), .A2(n1236), .ZN(n1234) );
INV_X1 U944 ( .A(n1191), .ZN(n1034) );
XOR2_X1 U945 ( .A(n1045), .B(n1237), .Z(n1191) );
XNOR2_X1 U946 ( .A(KEYINPUT14), .B(n1046), .ZN(n1237) );
INV_X1 U947 ( .A(G472), .ZN(n1046) );
NOR2_X1 U948 ( .A1(n1123), .A2(G902), .ZN(n1045) );
XOR2_X1 U949 ( .A(n1238), .B(n1239), .Z(n1123) );
XOR2_X1 U950 ( .A(n1240), .B(n1241), .Z(n1239) );
NAND2_X1 U951 ( .A1(KEYINPUT48), .A2(n1242), .ZN(n1241) );
INV_X1 U952 ( .A(G119), .ZN(n1242) );
NAND2_X1 U953 ( .A1(n1236), .A2(G210), .ZN(n1240) );
NOR2_X1 U954 ( .A1(G953), .A2(G237), .ZN(n1236) );
XOR2_X1 U955 ( .A(n1128), .B(n1243), .Z(n1238) );
XOR2_X1 U956 ( .A(n1244), .B(n1245), .Z(n1128) );
XNOR2_X1 U957 ( .A(G101), .B(n1173), .ZN(n1244) );
AND2_X1 U958 ( .A1(n1202), .A2(n1023), .ZN(n992) );
NOR2_X1 U959 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
INV_X1 U960 ( .A(n1194), .ZN(n1021) );
NAND2_X1 U961 ( .A1(G221), .A2(n1246), .ZN(n1194) );
XNOR2_X1 U962 ( .A(n1043), .B(G469), .ZN(n1022) );
AND2_X1 U963 ( .A1(n1247), .A2(n1248), .ZN(n1043) );
XNOR2_X1 U964 ( .A(KEYINPUT10), .B(n1207), .ZN(n1248) );
XOR2_X1 U965 ( .A(n1249), .B(n1250), .Z(n1247) );
XOR2_X1 U966 ( .A(n1131), .B(n1251), .Z(n1250) );
NAND2_X1 U967 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1173), .ZN(n1253) );
XOR2_X1 U969 ( .A(KEYINPUT50), .B(n1255), .Z(n1252) );
NOR2_X1 U970 ( .A1(n1254), .A2(n1173), .ZN(n1255) );
XOR2_X1 U971 ( .A(n1256), .B(n1069), .Z(n1173) );
NAND2_X1 U972 ( .A1(n1257), .A2(n1258), .ZN(n1131) );
NAND3_X1 U973 ( .A1(G227), .A2(n1006), .A3(n1259), .ZN(n1258) );
XNOR2_X1 U974 ( .A(G110), .B(G140), .ZN(n1259) );
NAND2_X1 U975 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
NAND2_X1 U976 ( .A1(G227), .A2(n1006), .ZN(n1261) );
XNOR2_X1 U977 ( .A(n1262), .B(G110), .ZN(n1260) );
NAND2_X1 U978 ( .A1(KEYINPUT3), .A2(n1245), .ZN(n1249) );
XNOR2_X1 U979 ( .A(n1075), .B(n1263), .ZN(n1245) );
NOR2_X1 U980 ( .A1(KEYINPUT42), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U981 ( .A(G134), .B(G137), .ZN(n1264) );
INV_X1 U982 ( .A(G131), .ZN(n1075) );
AND2_X1 U983 ( .A1(n1155), .A2(n1265), .ZN(n1202) );
NAND2_X1 U984 ( .A1(n1015), .A2(n1266), .ZN(n1265) );
NAND4_X1 U985 ( .A1(G953), .A2(G902), .A3(n1197), .A4(n1089), .ZN(n1266) );
INV_X1 U986 ( .A(G898), .ZN(n1089) );
NAND3_X1 U987 ( .A1(n1197), .A2(n1006), .A3(G952), .ZN(n1015) );
NAND2_X1 U988 ( .A1(G237), .A2(G234), .ZN(n1197) );
NOR2_X1 U989 ( .A1(n1007), .A2(n1009), .ZN(n1155) );
AND2_X1 U990 ( .A1(G214), .A2(n1267), .ZN(n1009) );
INV_X1 U991 ( .A(n1189), .ZN(n1007) );
XOR2_X1 U992 ( .A(n1048), .B(KEYINPUT11), .Z(n1189) );
XOR2_X1 U993 ( .A(n1268), .B(n1137), .Z(n1048) );
NAND2_X1 U994 ( .A1(G210), .A2(n1267), .ZN(n1137) );
NAND2_X1 U995 ( .A1(n1207), .A2(n1269), .ZN(n1267) );
INV_X1 U996 ( .A(G237), .ZN(n1269) );
NAND2_X1 U997 ( .A1(n1270), .A2(n1207), .ZN(n1268) );
XOR2_X1 U998 ( .A(n1172), .B(n1271), .Z(n1270) );
XNOR2_X1 U999 ( .A(n1133), .B(n1174), .ZN(n1271) );
NAND2_X1 U1000 ( .A1(G224), .A2(n1006), .ZN(n1174) );
INV_X1 U1001 ( .A(G953), .ZN(n1006) );
XNOR2_X1 U1002 ( .A(n1092), .B(n1272), .ZN(n1133) );
XNOR2_X1 U1003 ( .A(n1273), .B(n1274), .ZN(n1272) );
NOR2_X1 U1004 ( .A1(KEYINPUT12), .A2(n1088), .ZN(n1274) );
XNOR2_X1 U1005 ( .A(G110), .B(n1232), .ZN(n1088) );
INV_X1 U1006 ( .A(G122), .ZN(n1232) );
NAND2_X1 U1007 ( .A1(n1275), .A2(KEYINPUT53), .ZN(n1273) );
XNOR2_X1 U1008 ( .A(n1093), .B(KEYINPUT44), .ZN(n1275) );
INV_X1 U1009 ( .A(n1254), .ZN(n1093) );
XNOR2_X1 U1010 ( .A(G101), .B(n1129), .ZN(n1254) );
XOR2_X1 U1011 ( .A(G107), .B(G104), .Z(n1129) );
XOR2_X1 U1012 ( .A(G119), .B(n1243), .Z(n1092) );
XOR2_X1 U1013 ( .A(G116), .B(G113), .Z(n1243) );
XOR2_X1 U1014 ( .A(n1276), .B(n1069), .Z(n1172) );
XOR2_X1 U1015 ( .A(G128), .B(G143), .Z(n1069) );
XOR2_X1 U1016 ( .A(n1277), .B(n1053), .Z(n1033) );
AND2_X1 U1017 ( .A1(G217), .A2(n1246), .ZN(n1053) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1207), .ZN(n1246) );
NAND2_X1 U1019 ( .A1(KEYINPUT25), .A2(n1051), .ZN(n1277) );
NAND2_X1 U1020 ( .A1(n1101), .A2(n1207), .ZN(n1051) );
INV_X1 U1021 ( .A(G902), .ZN(n1207) );
XNOR2_X1 U1022 ( .A(n1278), .B(n1279), .ZN(n1101) );
XOR2_X1 U1023 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U1024 ( .A(G110), .B(G119), .ZN(n1281) );
NAND2_X1 U1025 ( .A1(KEYINPUT5), .A2(n1221), .ZN(n1280) );
INV_X1 U1026 ( .A(G128), .ZN(n1221) );
XOR2_X1 U1027 ( .A(n1068), .B(n1282), .Z(n1278) );
NOR2_X1 U1028 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U1029 ( .A(KEYINPUT34), .B(n1285), .Z(n1284) );
NOR2_X1 U1030 ( .A1(n1286), .A2(G137), .ZN(n1285) );
NOR3_X1 U1031 ( .A1(n1287), .A2(G953), .A3(n1288), .ZN(n1286) );
NOR4_X1 U1032 ( .A1(G953), .A2(n1289), .A3(n1288), .A4(n1287), .ZN(n1283) );
INV_X1 U1033 ( .A(G221), .ZN(n1287) );
INV_X1 U1034 ( .A(G234), .ZN(n1288) );
XNOR2_X1 U1035 ( .A(G137), .B(KEYINPUT36), .ZN(n1289) );
XNOR2_X1 U1036 ( .A(n1276), .B(n1262), .ZN(n1068) );
INV_X1 U1037 ( .A(G140), .ZN(n1262) );
XNOR2_X1 U1038 ( .A(G125), .B(n1256), .ZN(n1276) );
XOR2_X1 U1039 ( .A(G146), .B(KEYINPUT49), .Z(n1256) );
endmodule


