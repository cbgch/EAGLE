//Key = 0100011110110100010100101101101100011011001100111101100000101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344;

XOR2_X1 U727 ( .A(n1011), .B(G107), .Z(G9) );
NAND2_X1 U728 ( .A1(KEYINPUT58), .A2(n1012), .ZN(n1011) );
NOR2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U730 ( .A1(G953), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1014) );
XOR2_X1 U731 ( .A(KEYINPUT28), .B(n1018), .Z(n1017) );
NOR2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR3_X1 U733 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR3_X1 U734 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1022) );
NOR4_X1 U735 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1025) );
NOR2_X1 U736 ( .A1(n1031), .A2(n1032), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR4_X1 U738 ( .A1(n1035), .A2(n1032), .A3(n1029), .A4(n1021), .ZN(n1019) );
NOR2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1036) );
NOR2_X1 U743 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U744 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR3_X1 U745 ( .A1(n1015), .A2(G953), .A3(G952), .ZN(n1013) );
AND4_X1 U746 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1015) );
NOR3_X1 U747 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
XNOR2_X1 U748 ( .A(n1055), .B(n1056), .ZN(n1054) );
XNOR2_X1 U749 ( .A(G478), .B(n1057), .ZN(n1053) );
NOR2_X1 U750 ( .A1(n1058), .A2(KEYINPUT45), .ZN(n1057) );
NAND4_X1 U751 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1052) );
OR2_X1 U752 ( .A1(n1045), .A2(KEYINPUT25), .ZN(n1062) );
NAND2_X1 U753 ( .A1(KEYINPUT25), .A2(n1039), .ZN(n1061) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U755 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NAND2_X1 U756 ( .A1(KEYINPUT16), .A2(n1067), .ZN(n1066) );
OR2_X1 U757 ( .A1(n1068), .A2(KEYINPUT16), .ZN(n1065) );
NAND2_X1 U758 ( .A1(n1068), .A2(G475), .ZN(n1059) );
NOR2_X1 U759 ( .A1(n1069), .A2(KEYINPUT37), .ZN(n1068) );
NOR3_X1 U760 ( .A1(n1070), .A2(n1027), .A3(n1071), .ZN(n1050) );
XOR2_X1 U761 ( .A(n1072), .B(n1073), .Z(G72) );
NOR2_X1 U762 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U763 ( .A(KEYINPUT3), .B(n1076), .Z(n1075) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1076) );
NAND2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1072) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1074), .ZN(n1078) );
XNOR2_X1 U767 ( .A(n1080), .B(n1081), .ZN(n1079) );
NAND3_X1 U768 ( .A1(G900), .A2(n1080), .A3(G953), .ZN(n1077) );
XNOR2_X1 U769 ( .A(n1082), .B(n1083), .ZN(n1080) );
XNOR2_X1 U770 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND2_X1 U771 ( .A1(KEYINPUT48), .A2(n1086), .ZN(n1084) );
XOR2_X1 U772 ( .A(KEYINPUT38), .B(n1087), .Z(n1086) );
XOR2_X1 U773 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U774 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U775 ( .A1(n1092), .A2(G953), .ZN(n1091) );
NOR2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
XOR2_X1 U778 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U779 ( .A1(G898), .A2(n1074), .ZN(n1095) );
NOR2_X1 U780 ( .A1(n1099), .A2(n1074), .ZN(n1088) );
NOR2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U784 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U785 ( .A1(n1102), .A2(n1108), .ZN(G63) );
NOR3_X1 U786 ( .A1(n1058), .A2(n1109), .A3(n1110), .ZN(n1108) );
NOR3_X1 U787 ( .A1(n1111), .A2(n1112), .A3(n1107), .ZN(n1110) );
INV_X1 U788 ( .A(G478), .ZN(n1112) );
NOR2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
AND2_X1 U790 ( .A1(n1016), .A2(G478), .ZN(n1113) );
NOR2_X1 U791 ( .A1(n1102), .A2(n1115), .ZN(G60) );
XOR2_X1 U792 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U793 ( .A1(n1064), .A2(n1107), .ZN(n1117) );
NOR2_X1 U794 ( .A1(KEYINPUT54), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U795 ( .A(n1119), .B(KEYINPUT11), .ZN(n1118) );
XNOR2_X1 U796 ( .A(n1120), .B(n1121), .ZN(G6) );
NOR3_X1 U797 ( .A1(n1122), .A2(KEYINPUT4), .A3(n1123), .ZN(n1121) );
INV_X1 U798 ( .A(n1124), .ZN(n1123) );
NOR2_X1 U799 ( .A1(n1102), .A2(n1125), .ZN(G57) );
XOR2_X1 U800 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U801 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U802 ( .A1(n1055), .A2(n1107), .ZN(n1129) );
XOR2_X1 U803 ( .A(n1130), .B(n1131), .Z(n1126) );
NOR2_X1 U804 ( .A1(G101), .A2(KEYINPUT9), .ZN(n1131) );
NOR2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(G54) );
XOR2_X1 U806 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U807 ( .A(n1136), .B(n1137), .ZN(n1135) );
XOR2_X1 U808 ( .A(n1138), .B(n1139), .Z(n1134) );
NOR2_X1 U809 ( .A1(n1140), .A2(n1107), .ZN(n1139) );
XOR2_X1 U810 ( .A(n1141), .B(KEYINPUT33), .Z(n1138) );
NAND2_X1 U811 ( .A1(KEYINPUT39), .A2(n1142), .ZN(n1141) );
XNOR2_X1 U812 ( .A(n1102), .B(KEYINPUT43), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1102), .A2(n1143), .ZN(G51) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U815 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U816 ( .A1(KEYINPUT10), .A2(n1148), .ZN(n1147) );
XOR2_X1 U817 ( .A(n1149), .B(n1150), .Z(n1144) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1107), .ZN(n1150) );
NAND2_X1 U819 ( .A1(G902), .A2(n1016), .ZN(n1107) );
NAND3_X1 U820 ( .A1(n1081), .A2(n1152), .A3(n1153), .ZN(n1016) );
XOR2_X1 U821 ( .A(n1093), .B(KEYINPUT60), .Z(n1153) );
NAND3_X1 U822 ( .A1(n1154), .A2(n1012), .A3(n1155), .ZN(n1093) );
NAND2_X1 U823 ( .A1(n1124), .A2(n1156), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1157), .A2(n1122), .ZN(n1156) );
NAND2_X1 U825 ( .A1(n1034), .A2(n1158), .ZN(n1122) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1041), .ZN(n1157) );
NAND3_X1 U827 ( .A1(n1124), .A2(n1158), .A3(n1033), .ZN(n1012) );
INV_X1 U828 ( .A(n1094), .ZN(n1152) );
NAND4_X1 U829 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1094) );
NAND2_X1 U830 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
XNOR2_X1 U831 ( .A(KEYINPUT55), .B(n1166), .ZN(n1165) );
INV_X1 U832 ( .A(n1167), .ZN(n1164) );
AND4_X1 U833 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1081) );
NOR4_X1 U834 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
INV_X1 U835 ( .A(n1176), .ZN(n1175) );
NOR2_X1 U836 ( .A1(KEYINPUT15), .A2(n1177), .ZN(n1173) );
NOR2_X1 U837 ( .A1(n1178), .A2(n1167), .ZN(n1172) );
NOR2_X1 U838 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U839 ( .A(n1181), .B(KEYINPUT24), .Z(n1180) );
AND3_X1 U840 ( .A1(n1182), .A2(n1183), .A3(KEYINPUT15), .ZN(n1179) );
NOR3_X1 U841 ( .A1(n1184), .A2(n1045), .A3(n1185), .ZN(n1182) );
NOR2_X1 U842 ( .A1(n1186), .A2(n1187), .ZN(n1170) );
AND3_X1 U843 ( .A1(n1188), .A2(n1034), .A3(n1041), .ZN(n1187) );
INV_X1 U844 ( .A(n1189), .ZN(n1186) );
XNOR2_X1 U845 ( .A(n1190), .B(KEYINPUT20), .ZN(n1151) );
NOR2_X1 U846 ( .A1(n1074), .A2(G952), .ZN(n1102) );
XOR2_X1 U847 ( .A(n1177), .B(n1191), .Z(G48) );
XNOR2_X1 U848 ( .A(G146), .B(KEYINPUT57), .ZN(n1191) );
NAND3_X1 U849 ( .A1(n1183), .A2(n1045), .A3(n1192), .ZN(n1177) );
XNOR2_X1 U850 ( .A(G143), .B(n1189), .ZN(G45) );
NAND4_X1 U851 ( .A1(n1193), .A2(n1045), .A3(n1041), .A4(n1194), .ZN(n1189) );
NOR3_X1 U852 ( .A1(n1167), .A2(n1184), .A3(n1195), .ZN(n1194) );
XNOR2_X1 U853 ( .A(G140), .B(n1168), .ZN(G42) );
NAND3_X1 U854 ( .A1(n1040), .A2(n1034), .A3(n1188), .ZN(n1168) );
XNOR2_X1 U855 ( .A(G137), .B(n1169), .ZN(G39) );
NAND3_X1 U856 ( .A1(n1188), .A2(n1183), .A3(n1159), .ZN(n1169) );
XNOR2_X1 U857 ( .A(G134), .B(n1176), .ZN(G36) );
NAND3_X1 U858 ( .A1(n1041), .A2(n1033), .A3(n1188), .ZN(n1176) );
XOR2_X1 U859 ( .A(G131), .B(n1196), .Z(G33) );
NOR4_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1185), .A4(n1199), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
INV_X1 U862 ( .A(KEYINPUT59), .ZN(n1201) );
NOR3_X1 U863 ( .A1(n1032), .A2(n1045), .A3(n1184), .ZN(n1200) );
NOR2_X1 U864 ( .A1(KEYINPUT59), .A2(n1188), .ZN(n1197) );
NOR3_X1 U865 ( .A1(n1202), .A2(n1184), .A3(n1032), .ZN(n1188) );
OR3_X1 U866 ( .A1(n1070), .A2(n1027), .A3(n1028), .ZN(n1032) );
INV_X1 U867 ( .A(n1030), .ZN(n1070) );
XOR2_X1 U868 ( .A(G128), .B(n1203), .Z(G30) );
NOR2_X1 U869 ( .A1(n1167), .A2(n1181), .ZN(n1203) );
NAND4_X1 U870 ( .A1(n1183), .A2(n1033), .A3(n1045), .A4(n1204), .ZN(n1181) );
XNOR2_X1 U871 ( .A(G101), .B(n1205), .ZN(G3) );
NAND4_X1 U872 ( .A1(n1026), .A2(n1041), .A3(n1045), .A4(n1206), .ZN(n1205) );
XNOR2_X1 U873 ( .A(KEYINPUT49), .B(n1207), .ZN(n1206) );
INV_X1 U874 ( .A(n1202), .ZN(n1045) );
INV_X1 U875 ( .A(n1199), .ZN(n1041) );
NAND2_X1 U876 ( .A1(n1208), .A2(n1209), .ZN(G27) );
NAND2_X1 U877 ( .A1(n1174), .A2(n1210), .ZN(n1209) );
XOR2_X1 U878 ( .A(KEYINPUT31), .B(n1211), .Z(n1208) );
NOR2_X1 U879 ( .A1(n1174), .A2(n1210), .ZN(n1211) );
AND3_X1 U880 ( .A1(n1040), .A2(n1192), .A3(n1212), .ZN(n1174) );
NOR3_X1 U881 ( .A1(n1167), .A2(n1184), .A3(n1185), .ZN(n1192) );
INV_X1 U882 ( .A(n1204), .ZN(n1184) );
NAND2_X1 U883 ( .A1(n1021), .A2(n1213), .ZN(n1204) );
NAND4_X1 U884 ( .A1(G902), .A2(G953), .A3(n1214), .A4(n1215), .ZN(n1213) );
INV_X1 U885 ( .A(G900), .ZN(n1215) );
XOR2_X1 U886 ( .A(G122), .B(n1216), .Z(G24) );
NOR2_X1 U887 ( .A1(n1167), .A2(n1166), .ZN(n1216) );
OR4_X1 U888 ( .A1(n1023), .A2(n1217), .A3(n1195), .A4(n1218), .ZN(n1166) );
NAND2_X1 U889 ( .A1(n1212), .A2(n1158), .ZN(n1023) );
INV_X1 U890 ( .A(n1043), .ZN(n1158) );
NAND2_X1 U891 ( .A1(n1219), .A2(n1220), .ZN(n1043) );
XNOR2_X1 U892 ( .A(G119), .B(n1161), .ZN(G21) );
NAND4_X1 U893 ( .A1(n1026), .A2(n1212), .A3(n1183), .A4(n1207), .ZN(n1161) );
NOR2_X1 U894 ( .A1(n1220), .A2(n1219), .ZN(n1183) );
NOR2_X1 U895 ( .A1(n1029), .A2(n1167), .ZN(n1026) );
XNOR2_X1 U896 ( .A(G116), .B(n1162), .ZN(G18) );
NAND2_X1 U897 ( .A1(n1221), .A2(n1033), .ZN(n1162) );
NOR2_X1 U898 ( .A1(n1195), .A2(n1193), .ZN(n1033) );
XNOR2_X1 U899 ( .A(G113), .B(n1163), .ZN(G15) );
NAND2_X1 U900 ( .A1(n1221), .A2(n1034), .ZN(n1163) );
INV_X1 U901 ( .A(n1185), .ZN(n1034) );
NAND2_X1 U902 ( .A1(n1193), .A2(n1195), .ZN(n1185) );
INV_X1 U903 ( .A(n1217), .ZN(n1193) );
NOR4_X1 U904 ( .A1(n1199), .A2(n1039), .A3(n1167), .A4(n1218), .ZN(n1221) );
INV_X1 U905 ( .A(n1212), .ZN(n1039) );
NOR2_X1 U906 ( .A1(n1046), .A2(n1222), .ZN(n1212) );
INV_X1 U907 ( .A(n1047), .ZN(n1222) );
NAND2_X1 U908 ( .A1(n1219), .A2(n1223), .ZN(n1199) );
XNOR2_X1 U909 ( .A(KEYINPUT46), .B(n1224), .ZN(n1223) );
XNOR2_X1 U910 ( .A(G110), .B(n1154), .ZN(G12) );
NAND3_X1 U911 ( .A1(n1040), .A2(n1124), .A3(n1159), .ZN(n1154) );
INV_X1 U912 ( .A(n1029), .ZN(n1159) );
NAND2_X1 U913 ( .A1(n1195), .A2(n1217), .ZN(n1029) );
NAND2_X1 U914 ( .A1(n1225), .A2(n1226), .ZN(n1217) );
NAND2_X1 U915 ( .A1(n1069), .A2(n1227), .ZN(n1226) );
NAND2_X1 U916 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U917 ( .A1(G475), .A2(n1230), .ZN(n1229) );
NAND2_X1 U918 ( .A1(n1231), .A2(n1064), .ZN(n1225) );
INV_X1 U919 ( .A(G475), .ZN(n1064) );
NAND2_X1 U920 ( .A1(n1230), .A2(n1232), .ZN(n1231) );
NAND2_X1 U921 ( .A1(n1067), .A2(n1228), .ZN(n1232) );
INV_X1 U922 ( .A(KEYINPUT14), .ZN(n1228) );
INV_X1 U923 ( .A(n1069), .ZN(n1067) );
NOR2_X1 U924 ( .A1(n1233), .A2(G902), .ZN(n1069) );
INV_X1 U925 ( .A(n1119), .ZN(n1233) );
XNOR2_X1 U926 ( .A(n1234), .B(n1235), .ZN(n1119) );
XOR2_X1 U927 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U928 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U929 ( .A1(G122), .A2(KEYINPUT18), .ZN(n1238) );
XOR2_X1 U930 ( .A(n1240), .B(n1241), .Z(n1234) );
NOR2_X1 U931 ( .A1(KEYINPUT50), .A2(n1120), .ZN(n1241) );
INV_X1 U932 ( .A(G104), .ZN(n1120) );
XNOR2_X1 U933 ( .A(G113), .B(n1242), .ZN(n1240) );
NOR2_X1 U934 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U935 ( .A(n1245), .B(KEYINPUT19), .Z(n1244) );
NAND2_X1 U936 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR3_X1 U937 ( .A1(n1248), .A2(G953), .A3(n1249), .ZN(n1247) );
INV_X1 U938 ( .A(G143), .ZN(n1246) );
NOR4_X1 U939 ( .A1(G953), .A2(n1250), .A3(n1249), .A4(n1248), .ZN(n1243) );
XOR2_X1 U940 ( .A(G237), .B(KEYINPUT0), .Z(n1248) );
INV_X1 U941 ( .A(G214), .ZN(n1249) );
XNOR2_X1 U942 ( .A(G143), .B(KEYINPUT29), .ZN(n1250) );
INV_X1 U943 ( .A(KEYINPUT26), .ZN(n1230) );
NAND3_X1 U944 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1195) );
NAND2_X1 U945 ( .A1(G478), .A2(n1254), .ZN(n1253) );
OR3_X1 U946 ( .A1(n1254), .A2(G478), .A3(KEYINPUT63), .ZN(n1252) );
OR2_X1 U947 ( .A1(n1058), .A2(KEYINPUT2), .ZN(n1254) );
NAND2_X1 U948 ( .A1(n1058), .A2(KEYINPUT63), .ZN(n1251) );
NOR2_X1 U949 ( .A1(n1114), .A2(G902), .ZN(n1058) );
INV_X1 U950 ( .A(n1111), .ZN(n1114) );
XNOR2_X1 U951 ( .A(n1255), .B(n1256), .ZN(n1111) );
XOR2_X1 U952 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U953 ( .A1(G217), .A2(n1259), .ZN(n1257) );
XNOR2_X1 U954 ( .A(n1260), .B(n1261), .ZN(n1255) );
INV_X1 U955 ( .A(G134), .ZN(n1261) );
NAND2_X1 U956 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND2_X1 U957 ( .A1(G107), .A2(n1264), .ZN(n1263) );
XOR2_X1 U958 ( .A(KEYINPUT30), .B(n1265), .Z(n1262) );
NOR2_X1 U959 ( .A1(G107), .A2(n1264), .ZN(n1265) );
XOR2_X1 U960 ( .A(G122), .B(G116), .Z(n1264) );
NOR3_X1 U961 ( .A1(n1167), .A2(n1218), .A3(n1202), .ZN(n1124) );
NAND2_X1 U962 ( .A1(n1046), .A2(n1047), .ZN(n1202) );
NAND2_X1 U963 ( .A1(G221), .A2(n1266), .ZN(n1047) );
XOR2_X1 U964 ( .A(n1267), .B(n1140), .Z(n1046) );
INV_X1 U965 ( .A(G469), .ZN(n1140) );
NAND2_X1 U966 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U967 ( .A(n1270), .B(n1142), .Z(n1268) );
XNOR2_X1 U968 ( .A(n1082), .B(n1271), .ZN(n1142) );
XOR2_X1 U969 ( .A(n1272), .B(G128), .Z(n1082) );
NAND3_X1 U970 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1272) );
NAND2_X1 U971 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U972 ( .A1(n1278), .A2(n1279), .ZN(n1274) );
INV_X1 U973 ( .A(KEYINPUT17), .ZN(n1279) );
NAND2_X1 U974 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
XNOR2_X1 U975 ( .A(KEYINPUT44), .B(n1277), .ZN(n1280) );
NAND2_X1 U976 ( .A1(KEYINPUT17), .A2(n1282), .ZN(n1273) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
OR3_X1 U978 ( .A1(n1276), .A2(n1277), .A3(KEYINPUT44), .ZN(n1284) );
INV_X1 U979 ( .A(n1281), .ZN(n1276) );
XOR2_X1 U980 ( .A(G146), .B(KEYINPUT42), .Z(n1281) );
NAND2_X1 U981 ( .A1(KEYINPUT44), .A2(n1277), .ZN(n1283) );
XOR2_X1 U982 ( .A(G143), .B(KEYINPUT8), .Z(n1277) );
XNOR2_X1 U983 ( .A(n1285), .B(n1286), .ZN(n1270) );
INV_X1 U984 ( .A(n1136), .ZN(n1286) );
XNOR2_X1 U985 ( .A(n1287), .B(n1288), .ZN(n1136) );
NAND2_X1 U986 ( .A1(n1289), .A2(G227), .ZN(n1287) );
XNOR2_X1 U987 ( .A(G953), .B(KEYINPUT56), .ZN(n1289) );
NAND2_X1 U988 ( .A1(KEYINPUT61), .A2(n1137), .ZN(n1285) );
XOR2_X1 U989 ( .A(G140), .B(G110), .Z(n1137) );
INV_X1 U990 ( .A(n1207), .ZN(n1218) );
NAND2_X1 U991 ( .A1(n1021), .A2(n1290), .ZN(n1207) );
NAND4_X1 U992 ( .A1(G902), .A2(G953), .A3(n1214), .A4(n1101), .ZN(n1290) );
INV_X1 U993 ( .A(G898), .ZN(n1101) );
NAND3_X1 U994 ( .A1(n1214), .A2(n1074), .A3(G952), .ZN(n1021) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1214) );
NAND2_X1 U996 ( .A1(n1030), .A2(n1291), .ZN(n1167) );
OR2_X1 U997 ( .A1(n1028), .A2(n1027), .ZN(n1291) );
NOR2_X1 U998 ( .A1(n1292), .A2(n1190), .ZN(n1027) );
XNOR2_X1 U999 ( .A(n1048), .B(KEYINPUT41), .ZN(n1028) );
NAND2_X1 U1000 ( .A1(n1190), .A2(n1292), .ZN(n1048) );
NAND4_X1 U1001 ( .A1(n1293), .A2(n1269), .A3(n1294), .A4(n1295), .ZN(n1292) );
NAND2_X1 U1002 ( .A1(KEYINPUT34), .A2(n1296), .ZN(n1295) );
NAND2_X1 U1003 ( .A1(n1297), .A2(n1146), .ZN(n1296) );
XNOR2_X1 U1004 ( .A(KEYINPUT62), .B(n1298), .ZN(n1297) );
NAND2_X1 U1005 ( .A1(n1299), .A2(n1300), .ZN(n1294) );
INV_X1 U1006 ( .A(KEYINPUT34), .ZN(n1300) );
NAND2_X1 U1007 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND3_X1 U1008 ( .A1(KEYINPUT62), .A2(n1146), .A3(n1298), .ZN(n1302) );
OR2_X1 U1009 ( .A1(n1298), .A2(KEYINPUT62), .ZN(n1301) );
OR2_X1 U1010 ( .A1(n1146), .A2(n1298), .ZN(n1293) );
XOR2_X1 U1011 ( .A(n1303), .B(n1304), .Z(n1298) );
XOR2_X1 U1012 ( .A(KEYINPUT40), .B(n1149), .Z(n1304) );
NOR2_X1 U1013 ( .A1(n1100), .A2(G953), .ZN(n1149) );
INV_X1 U1014 ( .A(G224), .ZN(n1100) );
NAND2_X1 U1015 ( .A1(KEYINPUT35), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1016 ( .A(KEYINPUT47), .B(n1148), .Z(n1305) );
XNOR2_X1 U1017 ( .A(n1306), .B(n1307), .ZN(n1148) );
XNOR2_X1 U1018 ( .A(G125), .B(KEYINPUT23), .ZN(n1306) );
NAND2_X1 U1019 ( .A1(n1308), .A2(n1309), .ZN(n1146) );
NAND2_X1 U1020 ( .A1(n1310), .A2(n1098), .ZN(n1309) );
XOR2_X1 U1021 ( .A(KEYINPUT1), .B(n1311), .Z(n1308) );
NOR2_X1 U1022 ( .A1(n1098), .A2(n1310), .ZN(n1311) );
XOR2_X1 U1023 ( .A(n1097), .B(KEYINPUT7), .Z(n1310) );
XOR2_X1 U1024 ( .A(n1312), .B(n1313), .Z(n1097) );
XOR2_X1 U1025 ( .A(G119), .B(G116), .Z(n1313) );
XNOR2_X1 U1026 ( .A(G113), .B(n1271), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(n1314), .B(n1315), .ZN(n1271) );
XOR2_X1 U1028 ( .A(KEYINPUT21), .B(G107), .Z(n1315) );
XNOR2_X1 U1029 ( .A(G104), .B(G101), .ZN(n1314) );
XNOR2_X1 U1030 ( .A(G110), .B(G122), .ZN(n1098) );
AND2_X1 U1031 ( .A1(G210), .A2(n1316), .ZN(n1190) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1316), .ZN(n1030) );
NAND2_X1 U1033 ( .A1(n1269), .A2(n1317), .ZN(n1316) );
NOR2_X1 U1034 ( .A1(n1224), .A2(n1219), .ZN(n1040) );
AND2_X1 U1035 ( .A1(n1318), .A2(n1049), .ZN(n1219) );
NAND2_X1 U1036 ( .A1(n1319), .A2(n1320), .ZN(n1049) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1266), .ZN(n1320) );
XOR2_X1 U1038 ( .A(KEYINPUT36), .B(n1071), .Z(n1318) );
NOR3_X1 U1039 ( .A1(n1321), .A2(n1319), .A3(n1106), .ZN(n1071) );
INV_X1 U1040 ( .A(G217), .ZN(n1106) );
NOR2_X1 U1041 ( .A1(n1104), .A2(G902), .ZN(n1319) );
XOR2_X1 U1042 ( .A(n1322), .B(n1323), .Z(n1104) );
XNOR2_X1 U1043 ( .A(n1324), .B(n1236), .ZN(n1323) );
XNOR2_X1 U1044 ( .A(n1325), .B(n1085), .ZN(n1236) );
XNOR2_X1 U1045 ( .A(G140), .B(n1210), .ZN(n1085) );
INV_X1 U1046 ( .A(G125), .ZN(n1210) );
NAND2_X1 U1047 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
NAND2_X1 U1048 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1259), .ZN(n1329) );
INV_X1 U1050 ( .A(G137), .ZN(n1328) );
XOR2_X1 U1051 ( .A(n1330), .B(KEYINPUT12), .Z(n1326) );
NAND3_X1 U1052 ( .A1(G221), .A2(n1259), .A3(G137), .ZN(n1330) );
AND2_X1 U1053 ( .A1(G234), .A2(n1074), .ZN(n1259) );
XNOR2_X1 U1054 ( .A(G110), .B(n1331), .ZN(n1322) );
XOR2_X1 U1055 ( .A(G128), .B(G119), .Z(n1331) );
INV_X1 U1056 ( .A(n1266), .ZN(n1321) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1269), .ZN(n1266) );
INV_X1 U1058 ( .A(n1220), .ZN(n1224) );
XOR2_X1 U1059 ( .A(n1332), .B(n1055), .Z(n1220) );
INV_X1 U1060 ( .A(G472), .ZN(n1055) );
NAND2_X1 U1061 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XOR2_X1 U1062 ( .A(KEYINPUT52), .B(n1056), .Z(n1334) );
AND2_X1 U1063 ( .A1(n1335), .A2(n1336), .ZN(n1056) );
XNOR2_X1 U1064 ( .A(KEYINPUT27), .B(n1269), .ZN(n1336) );
INV_X1 U1065 ( .A(G902), .ZN(n1269) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1335) );
XNOR2_X1 U1067 ( .A(G101), .B(n1130), .ZN(n1338) );
NAND3_X1 U1068 ( .A1(n1317), .A2(n1074), .A3(G210), .ZN(n1130) );
INV_X1 U1069 ( .A(G953), .ZN(n1074) );
INV_X1 U1070 ( .A(G237), .ZN(n1317) );
NOR2_X1 U1071 ( .A1(KEYINPUT53), .A2(n1128), .ZN(n1337) );
XOR2_X1 U1072 ( .A(n1339), .B(n1340), .Z(n1128) );
XOR2_X1 U1073 ( .A(n1341), .B(n1342), .Z(n1340) );
XNOR2_X1 U1074 ( .A(G113), .B(G119), .ZN(n1342) );
NAND2_X1 U1075 ( .A1(KEYINPUT13), .A2(G116), .ZN(n1341) );
XNOR2_X1 U1076 ( .A(n1307), .B(n1288), .ZN(n1339) );
XOR2_X1 U1077 ( .A(n1087), .B(KEYINPUT5), .Z(n1288) );
XNOR2_X1 U1078 ( .A(n1343), .B(n1239), .ZN(n1087) );
XOR2_X1 U1079 ( .A(G131), .B(KEYINPUT51), .Z(n1239) );
XNOR2_X1 U1080 ( .A(G134), .B(G137), .ZN(n1343) );
XNOR2_X1 U1081 ( .A(n1258), .B(n1344), .ZN(n1307) );
NOR2_X1 U1082 ( .A1(KEYINPUT32), .A2(n1325), .ZN(n1344) );
INV_X1 U1083 ( .A(G146), .ZN(n1325) );
XNOR2_X1 U1084 ( .A(G128), .B(G143), .ZN(n1258) );
XNOR2_X1 U1085 ( .A(KEYINPUT6), .B(KEYINPUT22), .ZN(n1333) );
endmodule


