//Key = 1011000000111000011110110001000100011000001000011011001011111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337;

XOR2_X1 U719 ( .A(G107), .B(n1003), .Z(G9) );
NOR2_X1 U720 ( .A1(KEYINPUT38), .A2(n1004), .ZN(n1003) );
NOR2_X1 U721 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR4_X1 U722 ( .A1(G953), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1006) );
NOR2_X1 U723 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U724 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR3_X1 U725 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U726 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U727 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U728 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U729 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U730 ( .A1(n1025), .A2(n1026), .ZN(n1017) );
NOR2_X1 U731 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U732 ( .A1(n1020), .A2(n1029), .A3(n1026), .ZN(n1012) );
NOR2_X1 U733 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U734 ( .A1(n1032), .A2(n1016), .ZN(n1031) );
INV_X1 U735 ( .A(n1033), .ZN(n1016) );
NOR2_X1 U736 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U737 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U738 ( .A1(n1038), .A2(n1014), .ZN(n1030) );
INV_X1 U739 ( .A(n1039), .ZN(n1014) );
NOR2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U741 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
INV_X1 U742 ( .A(n1044), .ZN(n1010) );
NOR3_X1 U743 ( .A1(n1007), .A2(G953), .A3(G952), .ZN(n1005) );
AND4_X1 U744 ( .A1(n1045), .A2(n1039), .A3(n1046), .A4(n1047), .ZN(n1007) );
NOR4_X1 U745 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XOR2_X1 U746 ( .A(n1052), .B(KEYINPUT35), .Z(n1049) );
XNOR2_X1 U747 ( .A(n1053), .B(n1054), .ZN(n1046) );
XOR2_X1 U748 ( .A(n1055), .B(n1056), .Z(G72) );
NOR2_X1 U749 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
AND2_X1 U750 ( .A1(G227), .A2(G900), .ZN(n1057) );
NAND2_X1 U751 ( .A1(n1059), .A2(n1060), .ZN(n1055) );
NAND4_X1 U752 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
XOR2_X1 U753 ( .A(n1065), .B(KEYINPUT1), .Z(n1059) );
NAND2_X1 U754 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U755 ( .A1(n1063), .A2(n1064), .A3(n1062), .ZN(n1067) );
NAND3_X1 U756 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1062) );
XOR2_X1 U757 ( .A(n1071), .B(KEYINPUT18), .Z(n1070) );
INV_X1 U758 ( .A(n1072), .ZN(n1064) );
NAND2_X1 U759 ( .A1(n1071), .A2(n1073), .ZN(n1063) );
NAND2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(n1073) );
NAND2_X1 U761 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
XNOR2_X1 U762 ( .A(KEYINPUT34), .B(n1076), .ZN(n1074) );
XNOR2_X1 U763 ( .A(KEYINPUT22), .B(n1077), .ZN(n1068) );
NAND2_X1 U764 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U765 ( .A(KEYINPUT34), .B(n1076), .Z(n1078) );
NAND2_X1 U766 ( .A1(n1080), .A2(n1081), .ZN(n1071) );
XOR2_X1 U767 ( .A(KEYINPUT47), .B(n1082), .Z(n1080) );
INV_X1 U768 ( .A(n1061), .ZN(n1066) );
NAND2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1061) );
XNOR2_X1 U770 ( .A(KEYINPUT3), .B(n1058), .ZN(n1083) );
XOR2_X1 U771 ( .A(n1085), .B(n1086), .Z(G69) );
XOR2_X1 U772 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U773 ( .A1(G953), .A2(n1089), .ZN(n1088) );
NAND2_X1 U774 ( .A1(G898), .A2(G224), .ZN(n1089) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND2_X1 U777 ( .A1(n1094), .A2(n1058), .ZN(n1085) );
NOR2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(G66) );
NOR3_X1 U779 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NOR2_X1 U780 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U781 ( .A1(n1102), .A2(n1054), .ZN(n1100) );
XOR2_X1 U782 ( .A(KEYINPUT15), .B(n1103), .Z(n1097) );
NOR3_X1 U783 ( .A1(n1104), .A2(n1054), .A3(n1105), .ZN(n1103) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1106), .ZN(G63) );
XNOR2_X1 U785 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U786 ( .A1(n1109), .A2(n1104), .ZN(n1108) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1110), .ZN(G60) );
XOR2_X1 U788 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U789 ( .A1(n1113), .A2(n1104), .ZN(n1111) );
XOR2_X1 U790 ( .A(G104), .B(n1114), .Z(G6) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1115), .ZN(G57) );
XOR2_X1 U792 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U793 ( .A1(KEYINPUT48), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U794 ( .A(n1119), .B(n1120), .ZN(n1118) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U796 ( .A1(n1123), .A2(n1104), .ZN(n1122) );
NAND2_X1 U797 ( .A1(KEYINPUT36), .A2(n1124), .ZN(n1121) );
XOR2_X1 U798 ( .A(KEYINPUT12), .B(n1125), .Z(n1124) );
NOR2_X1 U799 ( .A1(n1095), .A2(n1126), .ZN(G54) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U801 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND4_X1 U802 ( .A1(KEYINPUT56), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
NAND3_X1 U803 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
INV_X1 U804 ( .A(KEYINPUT21), .ZN(n1135) );
OR2_X1 U805 ( .A1(n1136), .A2(n1134), .ZN(n1132) );
NOR2_X1 U806 ( .A1(KEYINPUT41), .A2(n1137), .ZN(n1134) );
NAND2_X1 U807 ( .A1(KEYINPUT21), .A2(n1137), .ZN(n1131) );
XOR2_X1 U808 ( .A(n1138), .B(n1079), .Z(n1137) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1127) );
NOR2_X1 U810 ( .A1(n1141), .A2(n1104), .ZN(n1140) );
NAND2_X1 U811 ( .A1(G902), .A2(n1009), .ZN(n1104) );
NOR2_X1 U812 ( .A1(n1095), .A2(n1142), .ZN(G51) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U814 ( .A(n1090), .B(n1145), .ZN(n1144) );
XNOR2_X1 U815 ( .A(n1146), .B(n1147), .ZN(n1143) );
NAND4_X1 U816 ( .A1(G210), .A2(n1009), .A3(n1148), .A4(n1149), .ZN(n1147) );
NAND2_X1 U817 ( .A1(KEYINPUT46), .A2(G902), .ZN(n1149) );
NAND2_X1 U818 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NAND2_X1 U819 ( .A1(KEYINPUT46), .A2(G237), .ZN(n1150) );
INV_X1 U820 ( .A(n1102), .ZN(n1009) );
NOR2_X1 U821 ( .A1(n1094), .A2(n1084), .ZN(n1102) );
NAND4_X1 U822 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1084) );
NOR4_X1 U823 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
INV_X1 U824 ( .A(n1160), .ZN(n1159) );
NAND2_X1 U825 ( .A1(n1161), .A2(n1035), .ZN(n1154) );
NAND2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1152) );
NAND2_X1 U827 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U828 ( .A(n1027), .B(KEYINPUT5), .ZN(n1164) );
NAND4_X1 U829 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1094) );
NOR4_X1 U830 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1114), .ZN(n1169) );
AND2_X1 U831 ( .A1(n1028), .A2(n1173), .ZN(n1114) );
INV_X1 U832 ( .A(n1004), .ZN(n1170) );
NAND2_X1 U833 ( .A1(n1027), .A2(n1173), .ZN(n1004) );
AND3_X1 U834 ( .A1(n1033), .A2(n1174), .A3(n1022), .ZN(n1173) );
NOR2_X1 U835 ( .A1(n1175), .A2(n1176), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1058), .A2(G952), .ZN(n1095) );
XNOR2_X1 U837 ( .A(n1177), .B(n1178), .ZN(G48) );
NOR2_X1 U838 ( .A1(n1165), .A2(n1179), .ZN(n1178) );
NAND3_X1 U839 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G45) );
OR2_X1 U840 ( .A1(G143), .A2(KEYINPUT23), .ZN(n1182) );
NAND3_X1 U841 ( .A1(KEYINPUT23), .A2(G143), .A3(n1183), .ZN(n1181) );
NAND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1180) );
NAND2_X1 U843 ( .A1(KEYINPUT23), .A2(n1186), .ZN(n1185) );
XOR2_X1 U844 ( .A(KEYINPUT26), .B(G143), .Z(n1186) );
INV_X1 U845 ( .A(n1183), .ZN(n1184) );
NAND2_X1 U846 ( .A1(n1161), .A2(n1187), .ZN(n1183) );
XNOR2_X1 U847 ( .A(KEYINPUT40), .B(n1188), .ZN(n1187) );
AND3_X1 U848 ( .A1(n1041), .A2(n1022), .A3(n1189), .ZN(n1161) );
NOR3_X1 U849 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
XNOR2_X1 U850 ( .A(G140), .B(n1153), .ZN(G42) );
NAND2_X1 U851 ( .A1(n1193), .A2(n1194), .ZN(n1153) );
XNOR2_X1 U852 ( .A(n1195), .B(n1158), .ZN(G39) );
AND2_X1 U853 ( .A1(n1194), .A2(n1196), .ZN(n1158) );
XOR2_X1 U854 ( .A(n1157), .B(n1197), .Z(G36) );
XOR2_X1 U855 ( .A(KEYINPUT14), .B(G134), .Z(n1197) );
AND3_X1 U856 ( .A1(n1041), .A2(n1027), .A3(n1194), .ZN(n1157) );
XNOR2_X1 U857 ( .A(G131), .B(n1198), .ZN(G33) );
NAND2_X1 U858 ( .A1(KEYINPUT19), .A2(n1156), .ZN(n1198) );
AND3_X1 U859 ( .A1(n1028), .A2(n1041), .A3(n1194), .ZN(n1156) );
AND3_X1 U860 ( .A1(n1022), .A2(n1199), .A3(n1039), .ZN(n1194) );
NOR2_X1 U861 ( .A1(n1036), .A2(n1200), .ZN(n1039) );
INV_X1 U862 ( .A(n1037), .ZN(n1200) );
XNOR2_X1 U863 ( .A(n1201), .B(n1202), .ZN(G30) );
AND2_X1 U864 ( .A1(n1027), .A2(n1162), .ZN(n1202) );
INV_X1 U865 ( .A(n1179), .ZN(n1162) );
NAND3_X1 U866 ( .A1(n1203), .A2(n1022), .A3(n1204), .ZN(n1179) );
NOR3_X1 U867 ( .A1(n1188), .A2(n1191), .A3(n1045), .ZN(n1204) );
INV_X1 U868 ( .A(n1199), .ZN(n1191) );
XOR2_X1 U869 ( .A(G101), .B(n1172), .Z(G3) );
AND2_X1 U870 ( .A1(n1205), .A2(n1041), .ZN(n1172) );
XNOR2_X1 U871 ( .A(G125), .B(n1160), .ZN(G27) );
NAND4_X1 U872 ( .A1(n1193), .A2(n1206), .A3(n1035), .A4(n1199), .ZN(n1160) );
NAND2_X1 U873 ( .A1(n1207), .A2(n1208), .ZN(n1199) );
NAND3_X1 U874 ( .A1(n1209), .A2(n1044), .A3(n1072), .ZN(n1208) );
NOR2_X1 U875 ( .A1(n1210), .A2(G900), .ZN(n1072) );
INV_X1 U876 ( .A(n1092), .ZN(n1210) );
XNOR2_X1 U877 ( .A(KEYINPUT61), .B(n1151), .ZN(n1209) );
NOR3_X1 U878 ( .A1(n1042), .A2(n1165), .A3(n1043), .ZN(n1193) );
INV_X1 U879 ( .A(n1028), .ZN(n1165) );
XNOR2_X1 U880 ( .A(G122), .B(n1166), .ZN(G24) );
NAND4_X1 U881 ( .A1(n1211), .A2(n1033), .A3(n1212), .A4(n1051), .ZN(n1166) );
NOR2_X1 U882 ( .A1(n1042), .A2(n1203), .ZN(n1033) );
XNOR2_X1 U883 ( .A(G119), .B(n1167), .ZN(G21) );
NAND2_X1 U884 ( .A1(n1196), .A2(n1211), .ZN(n1167) );
NOR3_X1 U885 ( .A1(n1043), .A2(n1045), .A3(n1020), .ZN(n1196) );
INV_X1 U886 ( .A(n1213), .ZN(n1020) );
XNOR2_X1 U887 ( .A(G116), .B(n1214), .ZN(G18) );
NAND2_X1 U888 ( .A1(KEYINPUT42), .A2(n1176), .ZN(n1214) );
AND3_X1 U889 ( .A1(n1211), .A2(n1027), .A3(n1041), .ZN(n1176) );
NOR2_X1 U890 ( .A1(n1051), .A2(n1190), .ZN(n1027) );
INV_X1 U891 ( .A(n1212), .ZN(n1190) );
XNOR2_X1 U892 ( .A(n1175), .B(n1215), .ZN(G15) );
XOR2_X1 U893 ( .A(KEYINPUT63), .B(G113), .Z(n1215) );
AND3_X1 U894 ( .A1(n1041), .A2(n1211), .A3(n1028), .ZN(n1175) );
NOR2_X1 U895 ( .A1(n1212), .A2(n1192), .ZN(n1028) );
INV_X1 U896 ( .A(n1051), .ZN(n1192) );
AND2_X1 U897 ( .A1(n1206), .A2(n1174), .ZN(n1211) );
INV_X1 U898 ( .A(n1026), .ZN(n1206) );
NAND2_X1 U899 ( .A1(n1052), .A2(n1216), .ZN(n1026) );
INV_X1 U900 ( .A(n1024), .ZN(n1052) );
NOR2_X1 U901 ( .A1(n1045), .A2(n1203), .ZN(n1041) );
NAND2_X1 U902 ( .A1(n1217), .A2(n1218), .ZN(G12) );
NAND2_X1 U903 ( .A1(G110), .A2(n1219), .ZN(n1218) );
XOR2_X1 U904 ( .A(n1220), .B(KEYINPUT7), .Z(n1217) );
NAND2_X1 U905 ( .A1(n1171), .A2(n1221), .ZN(n1220) );
INV_X1 U906 ( .A(n1219), .ZN(n1171) );
NAND3_X1 U907 ( .A1(n1045), .A2(n1203), .A3(n1205), .ZN(n1219) );
AND3_X1 U908 ( .A1(n1022), .A2(n1174), .A3(n1213), .ZN(n1205) );
NOR2_X1 U909 ( .A1(n1212), .A2(n1051), .ZN(n1213) );
XOR2_X1 U910 ( .A(n1222), .B(n1113), .Z(n1051) );
INV_X1 U911 ( .A(G475), .ZN(n1113) );
OR2_X1 U912 ( .A1(n1112), .A2(G902), .ZN(n1222) );
XNOR2_X1 U913 ( .A(n1223), .B(n1224), .ZN(n1112) );
XOR2_X1 U914 ( .A(G104), .B(n1225), .Z(n1224) );
XOR2_X1 U915 ( .A(G122), .B(G113), .Z(n1225) );
XOR2_X1 U916 ( .A(n1226), .B(n1227), .Z(n1223) );
XOR2_X1 U917 ( .A(n1228), .B(n1229), .Z(n1226) );
NOR2_X1 U918 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U919 ( .A(KEYINPUT24), .B(n1082), .Z(n1231) );
INV_X1 U920 ( .A(n1081), .ZN(n1230) );
NAND2_X1 U921 ( .A1(n1232), .A2(KEYINPUT51), .ZN(n1228) );
XOR2_X1 U922 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR4_X1 U923 ( .A1(KEYINPUT52), .A2(G953), .A3(G237), .A4(n1235), .ZN(n1234) );
INV_X1 U924 ( .A(G214), .ZN(n1235) );
XNOR2_X1 U925 ( .A(G131), .B(G143), .ZN(n1233) );
XOR2_X1 U926 ( .A(n1050), .B(KEYINPUT4), .Z(n1212) );
XOR2_X1 U927 ( .A(n1236), .B(n1109), .Z(n1050) );
INV_X1 U928 ( .A(G478), .ZN(n1109) );
NAND2_X1 U929 ( .A1(n1107), .A2(n1151), .ZN(n1236) );
XNOR2_X1 U930 ( .A(n1237), .B(n1238), .ZN(n1107) );
XOR2_X1 U931 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U932 ( .A(G107), .B(n1241), .Z(n1240) );
NOR2_X1 U933 ( .A1(KEYINPUT29), .A2(n1242), .ZN(n1241) );
XOR2_X1 U934 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U935 ( .A(G134), .B(n1201), .ZN(n1244) );
NOR2_X1 U936 ( .A1(G143), .A2(KEYINPUT30), .ZN(n1243) );
AND3_X1 U937 ( .A1(G234), .A2(n1058), .A3(G217), .ZN(n1239) );
XOR2_X1 U938 ( .A(n1245), .B(n1246), .Z(n1237) );
XOR2_X1 U939 ( .A(G122), .B(G116), .Z(n1246) );
XNOR2_X1 U940 ( .A(KEYINPUT27), .B(KEYINPUT17), .ZN(n1245) );
AND2_X1 U941 ( .A1(n1035), .A2(n1247), .ZN(n1174) );
NAND2_X1 U942 ( .A1(n1248), .A2(n1207), .ZN(n1247) );
NAND3_X1 U943 ( .A1(n1044), .A2(n1058), .A3(n1249), .ZN(n1207) );
XNOR2_X1 U944 ( .A(G952), .B(KEYINPUT2), .ZN(n1249) );
NAND4_X1 U945 ( .A1(n1092), .A2(G902), .A3(n1044), .A4(n1093), .ZN(n1248) );
INV_X1 U946 ( .A(G898), .ZN(n1093) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1044) );
XNOR2_X1 U948 ( .A(G953), .B(KEYINPUT20), .ZN(n1092) );
INV_X1 U949 ( .A(n1188), .ZN(n1035) );
NAND2_X1 U950 ( .A1(n1036), .A2(n1037), .ZN(n1188) );
NAND2_X1 U951 ( .A1(G214), .A2(n1250), .ZN(n1037) );
NAND2_X1 U952 ( .A1(n1151), .A2(n1251), .ZN(n1250) );
NAND2_X1 U953 ( .A1(n1252), .A2(n1253), .ZN(n1036) );
NAND2_X1 U954 ( .A1(G210), .A2(n1254), .ZN(n1253) );
NAND2_X1 U955 ( .A1(n1151), .A2(n1255), .ZN(n1254) );
OR2_X1 U956 ( .A1(n1251), .A2(n1256), .ZN(n1255) );
NAND3_X1 U957 ( .A1(n1257), .A2(n1151), .A3(n1256), .ZN(n1252) );
XNOR2_X1 U958 ( .A(n1258), .B(n1259), .ZN(n1256) );
INV_X1 U959 ( .A(n1090), .ZN(n1259) );
XNOR2_X1 U960 ( .A(n1260), .B(n1261), .ZN(n1090) );
XNOR2_X1 U961 ( .A(n1221), .B(n1262), .ZN(n1261) );
XOR2_X1 U962 ( .A(KEYINPUT33), .B(G122), .Z(n1262) );
XNOR2_X1 U963 ( .A(n1119), .B(n1263), .ZN(n1260) );
XOR2_X1 U964 ( .A(n1264), .B(n1265), .Z(n1263) );
NOR2_X1 U965 ( .A1(G104), .A2(KEYINPUT6), .ZN(n1264) );
NAND3_X1 U966 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1258) );
NAND2_X1 U967 ( .A1(n1145), .A2(n1269), .ZN(n1268) );
NAND2_X1 U968 ( .A1(n1270), .A2(KEYINPUT10), .ZN(n1269) );
XNOR2_X1 U969 ( .A(KEYINPUT57), .B(n1146), .ZN(n1270) );
INV_X1 U970 ( .A(n1271), .ZN(n1145) );
NAND3_X1 U971 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1267) );
INV_X1 U972 ( .A(KEYINPUT60), .ZN(n1274) );
NAND2_X1 U973 ( .A1(n1275), .A2(n1276), .ZN(n1272) );
INV_X1 U974 ( .A(KEYINPUT57), .ZN(n1275) );
NAND3_X1 U975 ( .A1(n1146), .A2(n1277), .A3(KEYINPUT60), .ZN(n1266) );
NAND2_X1 U976 ( .A1(KEYINPUT57), .A2(n1276), .ZN(n1277) );
NAND2_X1 U977 ( .A1(KEYINPUT10), .A2(n1271), .ZN(n1276) );
XOR2_X1 U978 ( .A(G125), .B(n1278), .Z(n1271) );
INV_X1 U979 ( .A(n1273), .ZN(n1146) );
NAND2_X1 U980 ( .A1(G224), .A2(n1058), .ZN(n1273) );
NAND2_X1 U981 ( .A1(G237), .A2(G210), .ZN(n1257) );
AND2_X1 U982 ( .A1(n1216), .A2(n1024), .ZN(n1022) );
XOR2_X1 U983 ( .A(n1279), .B(n1141), .Z(n1024) );
INV_X1 U984 ( .A(G469), .ZN(n1141) );
NAND2_X1 U985 ( .A1(n1280), .A2(n1151), .ZN(n1279) );
XOR2_X1 U986 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U987 ( .A(n1136), .B(n1283), .Z(n1282) );
XNOR2_X1 U988 ( .A(KEYINPUT50), .B(n1284), .ZN(n1283) );
NOR2_X1 U989 ( .A1(KEYINPUT37), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U990 ( .A(n1286), .B(n1075), .ZN(n1285) );
INV_X1 U991 ( .A(n1079), .ZN(n1075) );
XNOR2_X1 U992 ( .A(n1287), .B(n1288), .ZN(n1079) );
NOR2_X1 U993 ( .A1(G128), .A2(KEYINPUT9), .ZN(n1288) );
NOR2_X1 U994 ( .A1(KEYINPUT62), .A2(n1138), .ZN(n1286) );
XNOR2_X1 U995 ( .A(n1289), .B(n1265), .ZN(n1138) );
XOR2_X1 U996 ( .A(G101), .B(G107), .Z(n1265) );
XNOR2_X1 U997 ( .A(KEYINPUT54), .B(n1290), .ZN(n1289) );
NOR2_X1 U998 ( .A1(G104), .A2(KEYINPUT55), .ZN(n1290) );
XNOR2_X1 U999 ( .A(n1130), .B(n1291), .ZN(n1281) );
NOR2_X1 U1000 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
AND2_X1 U1001 ( .A1(KEYINPUT16), .A2(n1139), .ZN(n1293) );
NOR2_X1 U1002 ( .A1(KEYINPUT45), .A2(n1139), .ZN(n1292) );
NAND2_X1 U1003 ( .A1(G227), .A2(n1058), .ZN(n1139) );
XNOR2_X1 U1004 ( .A(G140), .B(n1221), .ZN(n1130) );
XNOR2_X1 U1005 ( .A(n1048), .B(KEYINPUT44), .ZN(n1216) );
INV_X1 U1006 ( .A(n1023), .ZN(n1048) );
NAND2_X1 U1007 ( .A1(n1294), .A2(G221), .ZN(n1023) );
XOR2_X1 U1008 ( .A(n1295), .B(KEYINPUT28), .Z(n1294) );
INV_X1 U1009 ( .A(n1043), .ZN(n1203) );
NAND2_X1 U1010 ( .A1(n1296), .A2(n1297), .ZN(n1043) );
NAND2_X1 U1011 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1012 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U1013 ( .A1(n1098), .A2(n1302), .ZN(n1301) );
INV_X1 U1014 ( .A(KEYINPUT13), .ZN(n1300) );
NAND2_X1 U1015 ( .A1(n1303), .A2(n1053), .ZN(n1296) );
INV_X1 U1016 ( .A(n1098), .ZN(n1053) );
NOR2_X1 U1017 ( .A1(n1101), .A2(G902), .ZN(n1098) );
INV_X1 U1018 ( .A(n1105), .ZN(n1101) );
XNOR2_X1 U1019 ( .A(n1304), .B(n1305), .ZN(n1105) );
XNOR2_X1 U1020 ( .A(G137), .B(n1306), .ZN(n1305) );
NAND3_X1 U1021 ( .A1(G234), .A2(n1058), .A3(G221), .ZN(n1306) );
NAND3_X1 U1022 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1304) );
NAND2_X1 U1023 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1024 ( .A1(n1312), .A2(KEYINPUT11), .ZN(n1311) );
XNOR2_X1 U1025 ( .A(KEYINPUT58), .B(n1313), .ZN(n1312) );
XNOR2_X1 U1026 ( .A(G110), .B(n1314), .ZN(n1310) );
NAND3_X1 U1027 ( .A1(KEYINPUT8), .A2(n1315), .A3(n1316), .ZN(n1308) );
INV_X1 U1028 ( .A(n1313), .ZN(n1316) );
NAND2_X1 U1029 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
INV_X1 U1030 ( .A(KEYINPUT58), .ZN(n1317) );
NAND3_X1 U1031 ( .A1(n1319), .A2(n1320), .A3(n1313), .ZN(n1307) );
XNOR2_X1 U1032 ( .A(n1321), .B(n1227), .ZN(n1313) );
XNOR2_X1 U1033 ( .A(n1177), .B(KEYINPUT31), .ZN(n1227) );
INV_X1 U1034 ( .A(G146), .ZN(n1177) );
NAND3_X1 U1035 ( .A1(n1322), .A2(n1323), .A3(n1081), .ZN(n1321) );
NAND2_X1 U1036 ( .A1(G140), .A2(n1324), .ZN(n1081) );
NAND2_X1 U1037 ( .A1(n1082), .A2(n1325), .ZN(n1323) );
INV_X1 U1038 ( .A(KEYINPUT32), .ZN(n1325) );
NOR2_X1 U1039 ( .A1(n1324), .A2(G140), .ZN(n1082) );
INV_X1 U1040 ( .A(G125), .ZN(n1324) );
NAND2_X1 U1041 ( .A1(KEYINPUT32), .A2(G140), .ZN(n1322) );
INV_X1 U1042 ( .A(KEYINPUT8), .ZN(n1320) );
NAND2_X1 U1043 ( .A1(KEYINPUT58), .A2(n1318), .ZN(n1319) );
NAND2_X1 U1044 ( .A1(KEYINPUT11), .A2(n1326), .ZN(n1318) );
XNOR2_X1 U1045 ( .A(n1221), .B(n1314), .ZN(n1326) );
NOR2_X1 U1046 ( .A1(KEYINPUT43), .A2(n1327), .ZN(n1314) );
XNOR2_X1 U1047 ( .A(G119), .B(G128), .ZN(n1327) );
INV_X1 U1048 ( .A(G110), .ZN(n1221) );
NAND2_X1 U1049 ( .A1(n1302), .A2(n1328), .ZN(n1303) );
OR2_X1 U1050 ( .A1(n1298), .A2(KEYINPUT13), .ZN(n1328) );
XNOR2_X1 U1051 ( .A(n1054), .B(KEYINPUT25), .ZN(n1298) );
NAND2_X1 U1052 ( .A1(G217), .A2(n1295), .ZN(n1054) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1151), .ZN(n1295) );
INV_X1 U1054 ( .A(KEYINPUT49), .ZN(n1302) );
INV_X1 U1055 ( .A(n1042), .ZN(n1045) );
XOR2_X1 U1056 ( .A(n1329), .B(n1123), .Z(n1042) );
INV_X1 U1057 ( .A(G472), .ZN(n1123) );
NAND2_X1 U1058 ( .A1(n1330), .A2(n1151), .ZN(n1329) );
INV_X1 U1059 ( .A(G902), .ZN(n1151) );
XOR2_X1 U1060 ( .A(n1117), .B(n1331), .Z(n1330) );
XNOR2_X1 U1061 ( .A(n1125), .B(n1119), .ZN(n1331) );
XOR2_X1 U1062 ( .A(G113), .B(n1332), .Z(n1119) );
XOR2_X1 U1063 ( .A(G119), .B(G116), .Z(n1332) );
XNOR2_X1 U1064 ( .A(n1136), .B(n1278), .ZN(n1125) );
XNOR2_X1 U1065 ( .A(n1201), .B(n1333), .ZN(n1278) );
NOR2_X1 U1066 ( .A1(KEYINPUT53), .A2(n1287), .ZN(n1333) );
XNOR2_X1 U1067 ( .A(G146), .B(G143), .ZN(n1287) );
INV_X1 U1068 ( .A(G128), .ZN(n1201) );
XOR2_X1 U1069 ( .A(n1334), .B(n1076), .Z(n1136) );
XNOR2_X1 U1070 ( .A(n1335), .B(n1336), .ZN(n1076) );
XNOR2_X1 U1071 ( .A(KEYINPUT59), .B(n1195), .ZN(n1336) );
INV_X1 U1072 ( .A(G137), .ZN(n1195) );
XNOR2_X1 U1073 ( .A(G131), .B(G134), .ZN(n1335) );
XNOR2_X1 U1074 ( .A(KEYINPUT39), .B(KEYINPUT0), .ZN(n1334) );
XOR2_X1 U1075 ( .A(n1337), .B(G101), .Z(n1117) );
NAND3_X1 U1076 ( .A1(n1251), .A2(n1058), .A3(G210), .ZN(n1337) );
INV_X1 U1077 ( .A(G953), .ZN(n1058) );
INV_X1 U1078 ( .A(G237), .ZN(n1251) );
endmodule


