//Key = 1110101010011111010001111010011011101011110011011100110100000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356;

XNOR2_X1 U738 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR3_X1 U740 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U742 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1027) );
XOR2_X1 U743 ( .A(n1032), .B(KEYINPUT40), .Z(n1031) );
NAND3_X1 U744 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NOR2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U749 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
AND2_X1 U751 ( .A1(n1049), .A2(KEYINPUT55), .ZN(n1047) );
XOR2_X1 U752 ( .A(n1050), .B(KEYINPUT12), .Z(n1029) );
NAND2_X1 U753 ( .A1(n1033), .A2(n1051), .ZN(n1050) );
NOR2_X1 U754 ( .A1(n1041), .A2(n1046), .ZN(n1033) );
INV_X1 U755 ( .A(n1052), .ZN(n1041) );
NAND3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1024) );
NAND3_X1 U757 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND4_X1 U759 ( .A1(n1061), .A2(n1049), .A3(n1028), .A4(n1062), .ZN(n1060) );
INV_X1 U760 ( .A(KEYINPUT55), .ZN(n1062) );
INV_X1 U761 ( .A(n1044), .ZN(n1061) );
NAND2_X1 U762 ( .A1(n1052), .A2(n1063), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR3_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1044), .ZN(n1052) );
NOR3_X1 U766 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U767 ( .A(n1053), .ZN(n1070) );
NAND4_X1 U768 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1053) );
NOR4_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1069), .A4(n1077), .ZN(n1074) );
XNOR2_X1 U770 ( .A(n1078), .B(n1079), .ZN(n1077) );
XNOR2_X1 U771 ( .A(n1080), .B(KEYINPUT22), .ZN(n1075) );
NOR3_X1 U772 ( .A1(n1081), .A2(n1035), .A3(n1066), .ZN(n1073) );
NOR2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U774 ( .A(KEYINPUT52), .B(n1084), .Z(n1072) );
AND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1084) );
XOR2_X1 U776 ( .A(n1085), .B(KEYINPUT31), .Z(n1083) );
XOR2_X1 U777 ( .A(KEYINPUT49), .B(n1086), .Z(n1071) );
XOR2_X1 U778 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1089) );
NAND3_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1087) );
NAND2_X1 U782 ( .A1(KEYINPUT3), .A2(n1094), .ZN(n1093) );
NAND3_X1 U783 ( .A1(n1095), .A2(n1054), .A3(n1096), .ZN(n1094) );
NAND2_X1 U784 ( .A1(n1097), .A2(n1054), .ZN(n1092) );
NAND2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1095), .ZN(n1099) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
OR2_X1 U788 ( .A1(n1096), .A2(KEYINPUT6), .ZN(n1102) );
INV_X1 U789 ( .A(n1103), .ZN(n1096) );
OR2_X1 U790 ( .A1(n1103), .A2(KEYINPUT3), .ZN(n1101) );
NAND3_X1 U791 ( .A1(KEYINPUT6), .A2(n1103), .A3(n1104), .ZN(n1098) );
NAND4_X1 U792 ( .A1(n1103), .A2(n1105), .A3(KEYINPUT6), .A4(G953), .ZN(n1091) );
XNOR2_X1 U793 ( .A(n1106), .B(n1107), .ZN(n1103) );
XNOR2_X1 U794 ( .A(n1108), .B(n1109), .ZN(n1107) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(G69) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1090), .ZN(n1113) );
XNOR2_X1 U798 ( .A(G953), .B(KEYINPUT19), .ZN(n1090) );
AND2_X1 U799 ( .A1(G224), .A2(G898), .ZN(n1114) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
NAND2_X1 U801 ( .A1(G953), .A2(n1117), .ZN(n1116) );
XNOR2_X1 U802 ( .A(KEYINPUT17), .B(n1118), .ZN(n1115) );
NAND2_X1 U803 ( .A1(n1054), .A2(n1119), .ZN(n1110) );
NAND2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(G66) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U809 ( .A1(KEYINPUT4), .A2(n1130), .ZN(n1126) );
NOR2_X1 U810 ( .A1(KEYINPUT4), .A2(n1130), .ZN(n1124) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1131), .ZN(G63) );
XOR2_X1 U812 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND3_X1 U813 ( .A1(G478), .A2(n1026), .A3(n1134), .ZN(n1133) );
XNOR2_X1 U814 ( .A(G902), .B(KEYINPUT41), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1135), .ZN(G60) );
NOR3_X1 U816 ( .A1(n1082), .A2(n1136), .A3(n1137), .ZN(n1135) );
NOR3_X1 U817 ( .A1(n1138), .A2(n1085), .A3(n1129), .ZN(n1137) );
INV_X1 U818 ( .A(n1139), .ZN(n1138) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1139), .ZN(n1136) );
AND2_X1 U820 ( .A1(n1026), .A2(G475), .ZN(n1140) );
NAND2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(G6) );
NAND2_X1 U822 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U823 ( .A(n1145), .B(KEYINPUT60), .Z(n1141) );
OR2_X1 U824 ( .A1(n1144), .A2(n1143), .ZN(n1145) );
XNOR2_X1 U825 ( .A(G104), .B(KEYINPUT23), .ZN(n1143) );
NOR3_X1 U826 ( .A1(n1122), .A2(n1146), .A3(n1147), .ZN(G57) );
NOR2_X1 U827 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1146) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1153), .ZN(n1159) );
XNOR2_X1 U834 ( .A(n1155), .B(KEYINPUT51), .ZN(n1153) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1152), .ZN(n1158) );
XNOR2_X1 U836 ( .A(n1160), .B(n1161), .ZN(n1155) );
XNOR2_X1 U837 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U838 ( .A1(KEYINPUT5), .A2(n1164), .ZN(n1163) );
XNOR2_X1 U839 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U840 ( .A1(KEYINPUT38), .A2(n1167), .ZN(n1162) );
XNOR2_X1 U841 ( .A(n1168), .B(n1169), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1129), .ZN(n1169) );
NOR3_X1 U843 ( .A1(n1171), .A2(n1122), .A3(n1172), .ZN(G54) );
NOR4_X1 U844 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1129), .ZN(n1172) );
NOR2_X1 U845 ( .A1(KEYINPUT1), .A2(n1176), .ZN(n1174) );
NOR2_X1 U846 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
INV_X1 U847 ( .A(KEYINPUT1), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1179), .ZN(n1171) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1129), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1176), .A2(n1180), .ZN(n1177) );
INV_X1 U851 ( .A(KEYINPUT61), .ZN(n1180) );
XOR2_X1 U852 ( .A(n1181), .B(n1182), .Z(n1176) );
NOR2_X1 U853 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NOR3_X1 U854 ( .A1(n1185), .A2(n1186), .A3(n1108), .ZN(n1184) );
INV_X1 U855 ( .A(KEYINPUT28), .ZN(n1185) );
NOR2_X1 U856 ( .A1(KEYINPUT28), .A2(n1187), .ZN(n1183) );
XNOR2_X1 U857 ( .A(n1188), .B(n1189), .ZN(n1181) );
NOR2_X1 U858 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U859 ( .A(n1192), .B(KEYINPUT15), .Z(n1191) );
NAND2_X1 U860 ( .A1(G110), .A2(n1193), .ZN(n1192) );
NOR2_X1 U861 ( .A1(G110), .A2(n1193), .ZN(n1190) );
NOR2_X1 U862 ( .A1(n1122), .A2(n1194), .ZN(G51) );
XNOR2_X1 U863 ( .A(n1118), .B(n1195), .ZN(n1194) );
XOR2_X1 U864 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U865 ( .A1(n1198), .A2(n1129), .ZN(n1197) );
NAND2_X1 U866 ( .A1(G902), .A2(n1026), .ZN(n1129) );
NAND3_X1 U867 ( .A1(n1104), .A2(n1199), .A3(n1120), .ZN(n1026) );
AND4_X1 U868 ( .A1(n1200), .A2(n1201), .A3(n1144), .A4(n1202), .ZN(n1120) );
AND4_X1 U869 ( .A1(n1021), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1202) );
NAND3_X1 U870 ( .A1(n1206), .A2(n1207), .A3(n1042), .ZN(n1021) );
NAND3_X1 U871 ( .A1(n1206), .A2(n1207), .A3(n1043), .ZN(n1144) );
NAND3_X1 U872 ( .A1(n1056), .A2(n1208), .A3(n1209), .ZN(n1200) );
XNOR2_X1 U873 ( .A(KEYINPUT53), .B(n1121), .ZN(n1199) );
INV_X1 U874 ( .A(n1095), .ZN(n1104) );
NAND4_X1 U875 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1095) );
NOR4_X1 U876 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
AND2_X1 U877 ( .A1(n1218), .A2(n1219), .ZN(n1212) );
NAND4_X1 U878 ( .A1(n1069), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1211) );
NAND2_X1 U879 ( .A1(n1068), .A2(n1223), .ZN(n1222) );
NAND4_X1 U880 ( .A1(n1056), .A2(n1051), .A3(n1028), .A4(n1224), .ZN(n1223) );
NAND2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
OR2_X1 U883 ( .A1(n1224), .A2(n1229), .ZN(n1210) );
INV_X1 U884 ( .A(KEYINPUT21), .ZN(n1224) );
NOR3_X1 U885 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1196) );
NOR2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
INV_X1 U887 ( .A(KEYINPUT11), .ZN(n1233) );
NOR2_X1 U888 ( .A1(KEYINPUT11), .A2(n1235), .ZN(n1231) );
NOR2_X1 U889 ( .A1(n1054), .A2(G952), .ZN(n1122) );
XOR2_X1 U890 ( .A(n1217), .B(n1236), .Z(G48) );
NOR2_X1 U891 ( .A1(KEYINPUT42), .A2(n1237), .ZN(n1236) );
AND3_X1 U892 ( .A1(n1043), .A2(n1051), .A3(n1238), .ZN(n1217) );
XNOR2_X1 U893 ( .A(G143), .B(n1219), .ZN(G45) );
NAND4_X1 U894 ( .A1(n1239), .A2(n1228), .A3(n1048), .A4(n1240), .ZN(n1219) );
NOR3_X1 U895 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
XNOR2_X1 U896 ( .A(G140), .B(n1218), .ZN(G42) );
NAND3_X1 U897 ( .A1(n1244), .A2(n1043), .A3(n1049), .ZN(n1218) );
XNOR2_X1 U898 ( .A(G137), .B(n1229), .ZN(G39) );
NAND3_X1 U899 ( .A1(n1245), .A2(n1068), .A3(n1244), .ZN(n1229) );
XOR2_X1 U900 ( .A(G134), .B(n1216), .Z(G36) );
AND3_X1 U901 ( .A1(n1048), .A2(n1042), .A3(n1244), .ZN(n1216) );
XNOR2_X1 U902 ( .A(G131), .B(n1246), .ZN(G33) );
NAND2_X1 U903 ( .A1(KEYINPUT44), .A2(n1215), .ZN(n1246) );
AND3_X1 U904 ( .A1(n1043), .A2(n1048), .A3(n1244), .ZN(n1215) );
NOR3_X1 U905 ( .A1(n1241), .A2(n1242), .A3(n1028), .ZN(n1244) );
NAND2_X1 U906 ( .A1(n1247), .A2(n1248), .ZN(n1028) );
XOR2_X1 U907 ( .A(n1067), .B(KEYINPUT20), .Z(n1247) );
XNOR2_X1 U908 ( .A(n1080), .B(KEYINPUT35), .ZN(n1067) );
INV_X1 U909 ( .A(n1051), .ZN(n1241) );
XOR2_X1 U910 ( .A(n1208), .B(KEYINPUT43), .Z(n1051) );
XNOR2_X1 U911 ( .A(G128), .B(n1249), .ZN(G30) );
NOR2_X1 U912 ( .A1(n1214), .A2(KEYINPUT63), .ZN(n1249) );
AND3_X1 U913 ( .A1(n1042), .A2(n1208), .A3(n1238), .ZN(n1214) );
NOR4_X1 U914 ( .A1(n1064), .A2(n1225), .A3(n1206), .A4(n1242), .ZN(n1238) );
XOR2_X1 U915 ( .A(n1250), .B(n1251), .Z(G3) );
NAND2_X1 U916 ( .A1(KEYINPUT62), .A2(G101), .ZN(n1251) );
NAND3_X1 U917 ( .A1(n1209), .A2(n1056), .A3(n1252), .ZN(n1250) );
XNOR2_X1 U918 ( .A(n1208), .B(KEYINPUT30), .ZN(n1252) );
XNOR2_X1 U919 ( .A(G125), .B(n1253), .ZN(G27) );
NAND4_X1 U920 ( .A1(n1254), .A2(n1049), .A3(n1255), .A4(n1058), .ZN(n1253) );
NOR2_X1 U921 ( .A1(n1242), .A2(n1064), .ZN(n1255) );
INV_X1 U922 ( .A(n1228), .ZN(n1064) );
INV_X1 U923 ( .A(n1220), .ZN(n1242) );
NAND2_X1 U924 ( .A1(n1044), .A2(n1256), .ZN(n1220) );
NAND4_X1 U925 ( .A1(n1257), .A2(G953), .A3(G902), .A4(n1258), .ZN(n1256) );
INV_X1 U926 ( .A(n1105), .ZN(n1257) );
XOR2_X1 U927 ( .A(G900), .B(KEYINPUT56), .Z(n1105) );
NOR2_X1 U928 ( .A1(n1068), .A2(n1206), .ZN(n1049) );
XNOR2_X1 U929 ( .A(n1043), .B(KEYINPUT2), .ZN(n1254) );
XNOR2_X1 U930 ( .A(G122), .B(n1201), .ZN(G24) );
NAND4_X1 U931 ( .A1(n1206), .A2(n1259), .A3(n1058), .A4(n1260), .ZN(n1201) );
NOR3_X1 U932 ( .A1(n1068), .A2(n1243), .A3(n1261), .ZN(n1260) );
XOR2_X1 U933 ( .A(G119), .B(n1262), .Z(G21) );
NOR2_X1 U934 ( .A1(KEYINPUT9), .A2(n1205), .ZN(n1262) );
NAND4_X1 U935 ( .A1(n1058), .A2(n1245), .A3(n1259), .A4(n1068), .ZN(n1205) );
XNOR2_X1 U936 ( .A(G116), .B(n1204), .ZN(G18) );
NAND3_X1 U937 ( .A1(n1209), .A2(n1042), .A3(n1058), .ZN(n1204) );
INV_X1 U938 ( .A(n1037), .ZN(n1058) );
NOR2_X1 U939 ( .A1(n1263), .A2(n1261), .ZN(n1042) );
XNOR2_X1 U940 ( .A(G113), .B(n1121), .ZN(G15) );
NAND2_X1 U941 ( .A1(n1227), .A2(n1209), .ZN(n1121) );
AND2_X1 U942 ( .A1(n1048), .A2(n1259), .ZN(n1209) );
NOR2_X1 U943 ( .A1(n1069), .A2(n1225), .ZN(n1048) );
NOR2_X1 U944 ( .A1(n1264), .A2(n1037), .ZN(n1227) );
NAND2_X1 U945 ( .A1(n1034), .A2(n1265), .ZN(n1037) );
INV_X1 U946 ( .A(n1043), .ZN(n1264) );
NOR2_X1 U947 ( .A1(n1239), .A2(n1243), .ZN(n1043) );
XNOR2_X1 U948 ( .A(G110), .B(n1203), .ZN(G12) );
NAND2_X1 U949 ( .A1(n1245), .A2(n1207), .ZN(n1203) );
AND3_X1 U950 ( .A1(n1225), .A2(n1259), .A3(n1208), .ZN(n1207) );
NOR2_X1 U951 ( .A1(n1034), .A2(n1035), .ZN(n1208) );
INV_X1 U952 ( .A(n1265), .ZN(n1035) );
NAND2_X1 U953 ( .A1(G221), .A2(n1266), .ZN(n1265) );
XOR2_X1 U954 ( .A(n1076), .B(KEYINPUT32), .Z(n1034) );
XOR2_X1 U955 ( .A(n1267), .B(n1175), .Z(n1076) );
INV_X1 U956 ( .A(G469), .ZN(n1175) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U958 ( .A(n1270), .B(n1271), .ZN(n1268) );
INV_X1 U959 ( .A(n1188), .ZN(n1271) );
XOR2_X1 U960 ( .A(n1167), .B(n1272), .Z(n1188) );
AND2_X1 U961 ( .A1(n1054), .A2(G227), .ZN(n1272) );
XNOR2_X1 U962 ( .A(n1187), .B(n1273), .ZN(n1270) );
NOR2_X1 U963 ( .A1(KEYINPUT10), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U964 ( .A(n1193), .B(n1275), .ZN(n1274) );
NOR2_X1 U965 ( .A1(G110), .A2(KEYINPUT7), .ZN(n1275) );
XNOR2_X1 U966 ( .A(n1108), .B(n1186), .ZN(n1187) );
AND2_X1 U967 ( .A1(n1276), .A2(n1277), .ZN(n1186) );
NAND2_X1 U968 ( .A1(n1278), .A2(n1166), .ZN(n1277) );
XOR2_X1 U969 ( .A(KEYINPUT36), .B(n1279), .Z(n1276) );
NOR2_X1 U970 ( .A1(n1278), .A2(n1166), .ZN(n1279) );
XNOR2_X1 U971 ( .A(G104), .B(G107), .ZN(n1278) );
NAND3_X1 U972 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1108) );
NAND2_X1 U973 ( .A1(n1283), .A2(n1237), .ZN(n1282) );
XNOR2_X1 U974 ( .A(n1284), .B(n1285), .ZN(n1283) );
XNOR2_X1 U975 ( .A(G143), .B(KEYINPUT57), .ZN(n1284) );
NAND3_X1 U976 ( .A1(G146), .A2(n1285), .A3(G143), .ZN(n1281) );
NAND3_X1 U977 ( .A1(G146), .A2(n1286), .A3(n1287), .ZN(n1280) );
AND2_X1 U978 ( .A1(n1228), .A2(n1288), .ZN(n1259) );
NAND2_X1 U979 ( .A1(n1044), .A2(n1289), .ZN(n1288) );
NAND4_X1 U980 ( .A1(G953), .A2(G902), .A3(n1258), .A4(n1117), .ZN(n1289) );
INV_X1 U981 ( .A(G898), .ZN(n1117) );
NAND3_X1 U982 ( .A1(n1258), .A2(n1054), .A3(G952), .ZN(n1044) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1258) );
NOR2_X1 U984 ( .A1(n1290), .A2(n1066), .ZN(n1228) );
INV_X1 U985 ( .A(n1248), .ZN(n1066) );
NAND2_X1 U986 ( .A1(G214), .A2(n1291), .ZN(n1248) );
INV_X1 U987 ( .A(n1080), .ZN(n1290) );
XOR2_X1 U988 ( .A(n1292), .B(n1198), .Z(n1080) );
NAND2_X1 U989 ( .A1(G210), .A2(n1291), .ZN(n1198) );
NAND2_X1 U990 ( .A1(n1293), .A2(n1269), .ZN(n1291) );
NAND3_X1 U991 ( .A1(n1294), .A2(n1269), .A3(n1295), .ZN(n1292) );
XOR2_X1 U992 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U993 ( .A1(n1118), .A2(n1298), .ZN(n1297) );
NAND2_X1 U994 ( .A1(n1234), .A2(n1299), .ZN(n1296) );
INV_X1 U995 ( .A(n1230), .ZN(n1299) );
NOR2_X1 U996 ( .A1(n1235), .A2(n1300), .ZN(n1230) );
NAND2_X1 U997 ( .A1(n1300), .A2(n1235), .ZN(n1234) );
NAND2_X1 U998 ( .A1(G224), .A2(n1054), .ZN(n1235) );
XNOR2_X1 U999 ( .A(G125), .B(n1301), .ZN(n1300) );
INV_X1 U1000 ( .A(n1168), .ZN(n1301) );
NAND2_X1 U1001 ( .A1(n1118), .A2(n1298), .ZN(n1294) );
INV_X1 U1002 ( .A(KEYINPUT8), .ZN(n1298) );
XOR2_X1 U1003 ( .A(n1302), .B(n1303), .Z(n1118) );
XOR2_X1 U1004 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U1005 ( .A(n1306), .B(n1307), .Z(n1302) );
XNOR2_X1 U1006 ( .A(n1308), .B(KEYINPUT46), .ZN(n1307) );
NAND2_X1 U1007 ( .A1(KEYINPUT48), .A2(G104), .ZN(n1308) );
INV_X1 U1008 ( .A(n1068), .ZN(n1225) );
XOR2_X1 U1009 ( .A(n1086), .B(KEYINPUT25), .Z(n1068) );
XOR2_X1 U1010 ( .A(n1309), .B(n1170), .Z(n1086) );
INV_X1 U1011 ( .A(G472), .ZN(n1170) );
NAND2_X1 U1012 ( .A1(n1310), .A2(n1269), .ZN(n1309) );
XOR2_X1 U1013 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U1014 ( .A(n1168), .B(n1313), .ZN(n1312) );
XNOR2_X1 U1015 ( .A(n1165), .B(n1152), .ZN(n1313) );
INV_X1 U1016 ( .A(n1154), .ZN(n1152) );
NOR2_X1 U1017 ( .A1(KEYINPUT54), .A2(n1314), .ZN(n1154) );
XOR2_X1 U1018 ( .A(KEYINPUT37), .B(n1315), .Z(n1314) );
NAND3_X1 U1019 ( .A1(n1293), .A2(n1054), .A3(G210), .ZN(n1165) );
INV_X1 U1020 ( .A(G237), .ZN(n1293) );
XOR2_X1 U1021 ( .A(n1316), .B(n1285), .Z(n1168) );
INV_X1 U1022 ( .A(n1286), .ZN(n1285) );
XOR2_X1 U1023 ( .A(G128), .B(KEYINPUT0), .Z(n1286) );
NAND2_X1 U1024 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1025 ( .A1(G146), .A2(n1287), .ZN(n1318) );
XOR2_X1 U1026 ( .A(KEYINPUT14), .B(n1319), .Z(n1317) );
NOR2_X1 U1027 ( .A1(G146), .A2(n1287), .ZN(n1319) );
XNOR2_X1 U1028 ( .A(n1167), .B(n1304), .ZN(n1311) );
XNOR2_X1 U1029 ( .A(n1166), .B(n1156), .ZN(n1304) );
INV_X1 U1030 ( .A(n1149), .ZN(n1156) );
XNOR2_X1 U1031 ( .A(G113), .B(G116), .ZN(n1149) );
INV_X1 U1032 ( .A(G101), .ZN(n1166) );
XNOR2_X1 U1033 ( .A(n1106), .B(KEYINPUT16), .ZN(n1167) );
XNOR2_X1 U1034 ( .A(G131), .B(n1320), .ZN(n1106) );
XOR2_X1 U1035 ( .A(G137), .B(G134), .Z(n1320) );
NOR2_X1 U1036 ( .A1(n1046), .A2(n1206), .ZN(n1245) );
INV_X1 U1037 ( .A(n1069), .ZN(n1206) );
XOR2_X1 U1038 ( .A(n1321), .B(n1128), .Z(n1069) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1266), .ZN(n1128) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1269), .ZN(n1266) );
OR2_X1 U1041 ( .A1(n1130), .A2(G902), .ZN(n1321) );
XNOR2_X1 U1042 ( .A(n1322), .B(n1323), .ZN(n1130) );
XOR2_X1 U1043 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1044 ( .A(G137), .B(G128), .Z(n1325) );
XNOR2_X1 U1045 ( .A(KEYINPUT26), .B(n1237), .ZN(n1324) );
XOR2_X1 U1046 ( .A(n1306), .B(n1326), .Z(n1322) );
XOR2_X1 U1047 ( .A(n1327), .B(n1109), .Z(n1326) );
XNOR2_X1 U1048 ( .A(G125), .B(n1193), .ZN(n1109) );
INV_X1 U1049 ( .A(G140), .ZN(n1193) );
AND3_X1 U1050 ( .A1(G221), .A2(n1054), .A3(G234), .ZN(n1327) );
XNOR2_X1 U1051 ( .A(G110), .B(n1315), .ZN(n1306) );
XOR2_X1 U1052 ( .A(G119), .B(KEYINPUT18), .Z(n1315) );
INV_X1 U1053 ( .A(n1056), .ZN(n1046) );
NOR2_X1 U1054 ( .A1(n1263), .A2(n1239), .ZN(n1056) );
INV_X1 U1055 ( .A(n1261), .ZN(n1239) );
XNOR2_X1 U1056 ( .A(n1328), .B(n1079), .ZN(n1261) );
AND2_X1 U1057 ( .A1(n1269), .A2(n1132), .ZN(n1079) );
NAND2_X1 U1058 ( .A1(n1329), .A2(n1330), .ZN(n1132) );
NAND2_X1 U1059 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1060 ( .A(KEYINPUT34), .B(n1333), .Z(n1329) );
NOR2_X1 U1061 ( .A1(n1334), .A2(n1332), .ZN(n1333) );
XOR2_X1 U1062 ( .A(n1335), .B(n1336), .Z(n1332) );
XNOR2_X1 U1063 ( .A(n1305), .B(n1337), .ZN(n1336) );
NOR2_X1 U1064 ( .A1(KEYINPUT50), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1065 ( .A(KEYINPUT27), .B(G116), .Z(n1338) );
XOR2_X1 U1066 ( .A(G122), .B(G107), .Z(n1305) );
NAND3_X1 U1067 ( .A1(n1339), .A2(n1340), .A3(KEYINPUT33), .ZN(n1335) );
NAND2_X1 U1068 ( .A1(G134), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1069 ( .A(KEYINPUT24), .B(n1342), .Z(n1339) );
NOR2_X1 U1070 ( .A1(G134), .A2(n1341), .ZN(n1342) );
XNOR2_X1 U1071 ( .A(n1287), .B(G128), .ZN(n1341) );
INV_X1 U1072 ( .A(G143), .ZN(n1287) );
XNOR2_X1 U1073 ( .A(n1331), .B(KEYINPUT47), .ZN(n1334) );
AND3_X1 U1074 ( .A1(G217), .A2(n1054), .A3(G234), .ZN(n1331) );
INV_X1 U1075 ( .A(G953), .ZN(n1054) );
INV_X1 U1076 ( .A(G902), .ZN(n1269) );
NAND2_X1 U1077 ( .A1(KEYINPUT45), .A2(n1078), .ZN(n1328) );
INV_X1 U1078 ( .A(G478), .ZN(n1078) );
INV_X1 U1079 ( .A(n1243), .ZN(n1263) );
XOR2_X1 U1080 ( .A(n1082), .B(n1085), .Z(n1243) );
INV_X1 U1081 ( .A(G475), .ZN(n1085) );
NOR2_X1 U1082 ( .A1(n1139), .A2(G902), .ZN(n1082) );
XNOR2_X1 U1083 ( .A(n1343), .B(n1344), .ZN(n1139) );
XOR2_X1 U1084 ( .A(G113), .B(n1345), .Z(n1344) );
XNOR2_X1 U1085 ( .A(KEYINPUT39), .B(n1346), .ZN(n1345) );
INV_X1 U1086 ( .A(G122), .ZN(n1346) );
XOR2_X1 U1087 ( .A(n1347), .B(G104), .Z(n1343) );
NAND2_X1 U1088 ( .A1(KEYINPUT13), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1089 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1090 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR3_X1 U1091 ( .A1(n1353), .A2(G953), .A3(G237), .ZN(n1352) );
XNOR2_X1 U1092 ( .A(G214), .B(KEYINPUT58), .ZN(n1353) );
NAND2_X1 U1093 ( .A1(n1354), .A2(KEYINPUT29), .ZN(n1351) );
XNOR2_X1 U1094 ( .A(G140), .B(n1355), .ZN(n1354) );
NOR2_X1 U1095 ( .A1(G125), .A2(KEYINPUT59), .ZN(n1355) );
XNOR2_X1 U1096 ( .A(G131), .B(n1356), .ZN(n1349) );
XNOR2_X1 U1097 ( .A(n1237), .B(G143), .ZN(n1356) );
INV_X1 U1098 ( .A(G146), .ZN(n1237) );
endmodule


