//Key = 0111010011110000110110011011010111100111000101000010111001101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;

XNOR2_X1 U781 ( .A(G107), .B(n1082), .ZN(G9) );
NOR2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(G75) );
NOR4_X1 U783 ( .A1(G953), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR3_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1099) );
NOR2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NOR3_X1 U796 ( .A1(n1108), .A2(n1113), .A3(n1102), .ZN(n1095) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR4_X1 U799 ( .A1(n1118), .A2(n1098), .A3(n1102), .A4(n1108), .ZN(n1090) );
INV_X1 U800 ( .A(n1119), .ZN(n1102) );
INV_X1 U801 ( .A(n1120), .ZN(n1098) );
NOR2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
INV_X1 U803 ( .A(n1123), .ZN(n1088) );
NOR3_X1 U804 ( .A1(n1085), .A2(G953), .A3(G952), .ZN(n1083) );
AND4_X1 U805 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1085) );
NOR4_X1 U806 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1127) );
XNOR2_X1 U807 ( .A(G469), .B(n1132), .ZN(n1131) );
XOR2_X1 U808 ( .A(n1133), .B(n1134), .Z(n1130) );
NAND2_X1 U809 ( .A1(KEYINPUT23), .A2(n1135), .ZN(n1134) );
INV_X1 U810 ( .A(n1136), .ZN(n1135) );
NOR3_X1 U811 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1126) );
NAND3_X1 U812 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1125) );
OR2_X1 U813 ( .A1(n1143), .A2(KEYINPUT31), .ZN(n1142) );
NAND3_X1 U814 ( .A1(KEYINPUT31), .A2(n1144), .A3(n1145), .ZN(n1141) );
OR2_X1 U815 ( .A1(n1145), .A2(n1144), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1146), .A2(KEYINPUT59), .ZN(n1144) );
NAND2_X1 U817 ( .A1(G475), .A2(n1147), .ZN(n1124) );
XOR2_X1 U818 ( .A(n1148), .B(n1149), .Z(G72) );
NOR2_X1 U819 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
AND2_X1 U820 ( .A1(G227), .A2(G900), .ZN(n1150) );
NAND2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NAND3_X1 U822 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
INV_X1 U823 ( .A(n1157), .ZN(n1155) );
OR2_X1 U824 ( .A1(n1156), .A2(n1154), .ZN(n1152) );
XNOR2_X1 U825 ( .A(n1158), .B(n1159), .ZN(n1154) );
XNOR2_X1 U826 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U828 ( .A(n1164), .B(KEYINPUT5), .Z(n1163) );
NAND2_X1 U829 ( .A1(G137), .A2(n1165), .ZN(n1164) );
XNOR2_X1 U830 ( .A(KEYINPUT45), .B(n1166), .ZN(n1165) );
NOR2_X1 U831 ( .A1(G137), .A2(n1166), .ZN(n1162) );
XOR2_X1 U832 ( .A(n1167), .B(n1168), .Z(n1158) );
NOR2_X1 U833 ( .A1(KEYINPUT36), .A2(n1169), .ZN(n1168) );
NAND2_X1 U834 ( .A1(n1151), .A2(n1170), .ZN(n1156) );
NAND2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U836 ( .A(n1173), .B(KEYINPUT44), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1174), .B(n1175), .Z(G69) );
XOR2_X1 U838 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR3_X1 U839 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NOR3_X1 U840 ( .A1(n1181), .A2(G953), .A3(G898), .ZN(n1180) );
AND2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
INV_X1 U842 ( .A(KEYINPUT7), .ZN(n1181) );
XOR2_X1 U843 ( .A(n1183), .B(n1184), .Z(n1178) );
XNOR2_X1 U844 ( .A(n1185), .B(n1186), .ZN(n1184) );
XOR2_X1 U845 ( .A(KEYINPUT21), .B(n1187), .Z(n1183) );
NOR2_X1 U846 ( .A1(KEYINPUT12), .A2(n1188), .ZN(n1187) );
NOR2_X1 U847 ( .A1(KEYINPUT22), .A2(n1189), .ZN(n1176) );
NOR2_X1 U848 ( .A1(n1190), .A2(G953), .ZN(n1189) );
NOR3_X1 U849 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
XNOR2_X1 U850 ( .A(n1194), .B(KEYINPUT52), .ZN(n1193) );
NOR2_X1 U851 ( .A1(n1195), .A2(n1182), .ZN(n1174) );
NOR2_X1 U852 ( .A1(G224), .A2(n1151), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1196), .A2(n1197), .ZN(G66) );
XOR2_X1 U854 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U855 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NOR2_X1 U856 ( .A1(n1196), .A2(n1202), .ZN(G63) );
XOR2_X1 U857 ( .A(n1203), .B(n1204), .Z(n1202) );
NAND3_X1 U858 ( .A1(n1205), .A2(n1206), .A3(G478), .ZN(n1203) );
NAND2_X1 U859 ( .A1(KEYINPUT54), .A2(n1201), .ZN(n1206) );
NAND2_X1 U860 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U861 ( .A(KEYINPUT54), .ZN(n1208) );
OR2_X1 U862 ( .A1(n1087), .A2(n1209), .ZN(n1207) );
NOR2_X1 U863 ( .A1(n1196), .A2(n1210), .ZN(G60) );
XNOR2_X1 U864 ( .A(n1211), .B(n1212), .ZN(n1210) );
XOR2_X1 U865 ( .A(KEYINPUT25), .B(n1213), .Z(n1212) );
NOR2_X1 U866 ( .A1(n1214), .A2(n1201), .ZN(n1213) );
XNOR2_X1 U867 ( .A(G104), .B(n1215), .ZN(G6) );
NOR2_X1 U868 ( .A1(n1196), .A2(n1216), .ZN(G57) );
XOR2_X1 U869 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U870 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1217) );
NOR2_X1 U872 ( .A1(KEYINPUT35), .A2(n1223), .ZN(n1222) );
NOR2_X1 U873 ( .A1(n1145), .A2(n1201), .ZN(n1221) );
NOR2_X1 U874 ( .A1(n1196), .A2(n1224), .ZN(G54) );
XOR2_X1 U875 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U876 ( .A(n1227), .B(n1228), .ZN(n1226) );
XNOR2_X1 U877 ( .A(KEYINPUT11), .B(n1229), .ZN(n1228) );
XOR2_X1 U878 ( .A(n1230), .B(n1231), .Z(n1225) );
XOR2_X1 U879 ( .A(n1232), .B(n1233), .Z(n1230) );
NOR2_X1 U880 ( .A1(n1234), .A2(n1201), .ZN(n1233) );
NAND2_X1 U881 ( .A1(KEYINPUT63), .A2(n1235), .ZN(n1232) );
NOR2_X1 U882 ( .A1(n1196), .A2(n1236), .ZN(G51) );
XOR2_X1 U883 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U884 ( .A(n1239), .B(n1240), .Z(n1237) );
NOR2_X1 U885 ( .A1(n1136), .A2(n1201), .ZN(n1240) );
NAND2_X1 U886 ( .A1(G902), .A2(n1087), .ZN(n1201) );
NAND3_X1 U887 ( .A1(n1241), .A2(n1172), .A3(n1242), .ZN(n1087) );
NOR3_X1 U888 ( .A1(n1192), .A2(n1194), .A3(n1173), .ZN(n1242) );
INV_X1 U889 ( .A(n1243), .ZN(n1194) );
AND2_X1 U890 ( .A1(n1244), .A2(n1104), .ZN(n1192) );
XOR2_X1 U891 ( .A(n1245), .B(KEYINPUT33), .Z(n1244) );
AND4_X1 U892 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1172) );
AND4_X1 U893 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
OR2_X1 U894 ( .A1(n1108), .A2(n1254), .ZN(n1251) );
XOR2_X1 U895 ( .A(KEYINPUT2), .B(n1255), .Z(n1254) );
INV_X1 U896 ( .A(n1256), .ZN(n1108) );
NAND2_X1 U897 ( .A1(n1257), .A2(n1258), .ZN(n1248) );
NAND2_X1 U898 ( .A1(n1259), .A2(n1104), .ZN(n1247) );
XOR2_X1 U899 ( .A(n1260), .B(KEYINPUT16), .Z(n1259) );
NAND2_X1 U900 ( .A1(n1261), .A2(n1122), .ZN(n1246) );
INV_X1 U901 ( .A(n1191), .ZN(n1241) );
NAND4_X1 U902 ( .A1(n1215), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1191) );
AND3_X1 U903 ( .A1(n1265), .A2(n1082), .A3(n1266), .ZN(n1264) );
NAND3_X1 U904 ( .A1(n1119), .A2(n1267), .A3(n1121), .ZN(n1082) );
NAND2_X1 U905 ( .A1(n1268), .A2(n1121), .ZN(n1263) );
NAND3_X1 U906 ( .A1(n1119), .A2(n1267), .A3(n1122), .ZN(n1215) );
NAND2_X1 U907 ( .A1(n1269), .A2(n1270), .ZN(n1239) );
INV_X1 U908 ( .A(n1271), .ZN(n1270) );
NAND2_X1 U909 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
NOR2_X1 U910 ( .A1(n1151), .A2(G952), .ZN(n1196) );
XNOR2_X1 U911 ( .A(G146), .B(n1274), .ZN(G48) );
NAND4_X1 U912 ( .A1(n1258), .A2(n1111), .A3(n1275), .A4(n1276), .ZN(n1274) );
NAND2_X1 U913 ( .A1(KEYINPUT32), .A2(n1277), .ZN(n1276) );
NAND2_X1 U914 ( .A1(n1278), .A2(n1279), .ZN(n1275) );
INV_X1 U915 ( .A(KEYINPUT32), .ZN(n1279) );
NAND2_X1 U916 ( .A1(n1280), .A2(n1115), .ZN(n1278) );
INV_X1 U917 ( .A(n1281), .ZN(n1280) );
XNOR2_X1 U918 ( .A(G143), .B(n1250), .ZN(G45) );
NAND4_X1 U919 ( .A1(n1282), .A2(n1110), .A3(n1283), .A4(n1104), .ZN(n1250) );
NOR2_X1 U920 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U921 ( .A(G140), .B(n1286), .ZN(G42) );
NAND3_X1 U922 ( .A1(n1255), .A2(n1256), .A3(KEYINPUT20), .ZN(n1286) );
AND4_X1 U923 ( .A1(n1282), .A2(n1122), .A3(n1287), .A4(n1288), .ZN(n1255) );
XNOR2_X1 U924 ( .A(G137), .B(n1253), .ZN(G39) );
NAND3_X1 U925 ( .A1(n1289), .A2(n1256), .A3(n1257), .ZN(n1253) );
XNOR2_X1 U926 ( .A(n1166), .B(n1173), .ZN(G36) );
AND2_X1 U927 ( .A1(n1261), .A2(n1121), .ZN(n1173) );
XOR2_X1 U928 ( .A(n1290), .B(n1291), .Z(G33) );
XNOR2_X1 U929 ( .A(G131), .B(KEYINPUT18), .ZN(n1291) );
NAND3_X1 U930 ( .A1(n1261), .A2(n1122), .A3(KEYINPUT19), .ZN(n1290) );
AND3_X1 U931 ( .A1(n1282), .A2(n1110), .A3(n1256), .ZN(n1261) );
NOR2_X1 U932 ( .A1(n1105), .A2(n1139), .ZN(n1256) );
INV_X1 U933 ( .A(n1277), .ZN(n1282) );
XNOR2_X1 U934 ( .A(n1292), .B(n1293), .ZN(G30) );
NOR2_X1 U935 ( .A1(n1294), .A2(n1260), .ZN(n1293) );
NAND3_X1 U936 ( .A1(n1121), .A2(n1287), .A3(n1257), .ZN(n1260) );
NOR2_X1 U937 ( .A1(n1277), .A2(n1288), .ZN(n1257) );
NAND2_X1 U938 ( .A1(n1115), .A2(n1281), .ZN(n1277) );
XOR2_X1 U939 ( .A(n1262), .B(n1295), .Z(G3) );
XNOR2_X1 U940 ( .A(G101), .B(KEYINPUT41), .ZN(n1295) );
NAND4_X1 U941 ( .A1(n1110), .A2(n1267), .A3(n1284), .A4(n1296), .ZN(n1262) );
XNOR2_X1 U942 ( .A(G125), .B(n1252), .ZN(G27) );
NAND4_X1 U943 ( .A1(n1258), .A2(n1120), .A3(n1281), .A4(n1288), .ZN(n1252) );
NAND2_X1 U944 ( .A1(n1297), .A2(n1298), .ZN(n1281) );
NAND3_X1 U945 ( .A1(G902), .A2(n1123), .A3(n1157), .ZN(n1298) );
NOR2_X1 U946 ( .A1(n1151), .A2(G900), .ZN(n1157) );
AND3_X1 U947 ( .A1(n1104), .A2(n1287), .A3(n1122), .ZN(n1258) );
XNOR2_X1 U948 ( .A(G122), .B(n1265), .ZN(G24) );
NAND4_X1 U949 ( .A1(n1299), .A2(n1119), .A3(n1129), .A4(n1092), .ZN(n1265) );
NOR2_X1 U950 ( .A1(n1287), .A2(n1111), .ZN(n1119) );
XOR2_X1 U951 ( .A(G119), .B(n1300), .Z(G21) );
NOR2_X1 U952 ( .A1(n1294), .A2(n1245), .ZN(n1300) );
NAND4_X1 U953 ( .A1(n1289), .A2(n1111), .A3(n1120), .A4(n1301), .ZN(n1245) );
INV_X1 U954 ( .A(n1288), .ZN(n1111) );
INV_X1 U955 ( .A(n1104), .ZN(n1294) );
XOR2_X1 U956 ( .A(G116), .B(n1302), .Z(G18) );
NOR3_X1 U957 ( .A1(n1303), .A2(KEYINPUT15), .A3(n1304), .ZN(n1302) );
INV_X1 U958 ( .A(n1121), .ZN(n1304) );
NOR2_X1 U959 ( .A1(n1092), .A2(n1285), .ZN(n1121) );
INV_X1 U960 ( .A(n1129), .ZN(n1285) );
XNOR2_X1 U961 ( .A(n1305), .B(n1243), .ZN(G15) );
NAND2_X1 U962 ( .A1(n1122), .A2(n1268), .ZN(n1243) );
INV_X1 U963 ( .A(n1303), .ZN(n1268) );
NAND2_X1 U964 ( .A1(n1110), .A2(n1299), .ZN(n1303) );
AND3_X1 U965 ( .A1(n1120), .A2(n1301), .A3(n1104), .ZN(n1299) );
NAND2_X1 U966 ( .A1(n1306), .A2(n1307), .ZN(n1120) );
OR3_X1 U967 ( .A1(n1308), .A2(n1117), .A3(KEYINPUT46), .ZN(n1307) );
NAND2_X1 U968 ( .A1(KEYINPUT46), .A2(n1115), .ZN(n1306) );
NOR2_X1 U969 ( .A1(n1288), .A2(n1287), .ZN(n1110) );
NOR2_X1 U970 ( .A1(n1129), .A2(n1284), .ZN(n1122) );
NAND2_X1 U971 ( .A1(KEYINPUT26), .A2(n1309), .ZN(n1305) );
NAND2_X1 U972 ( .A1(n1310), .A2(n1311), .ZN(G12) );
NAND2_X1 U973 ( .A1(n1312), .A2(n1227), .ZN(n1311) );
NAND2_X1 U974 ( .A1(n1313), .A2(G110), .ZN(n1310) );
NAND2_X1 U975 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
OR2_X1 U976 ( .A1(n1266), .A2(KEYINPUT34), .ZN(n1315) );
NAND2_X1 U977 ( .A1(KEYINPUT34), .A2(n1316), .ZN(n1314) );
INV_X1 U978 ( .A(n1312), .ZN(n1316) );
NOR2_X1 U979 ( .A1(KEYINPUT40), .A2(n1266), .ZN(n1312) );
NAND3_X1 U980 ( .A1(n1267), .A2(n1288), .A3(n1289), .ZN(n1266) );
NOR3_X1 U981 ( .A1(n1094), .A2(n1112), .A3(n1092), .ZN(n1289) );
INV_X1 U982 ( .A(n1284), .ZN(n1092) );
NOR2_X1 U983 ( .A1(n1317), .A2(n1138), .ZN(n1284) );
NOR2_X1 U984 ( .A1(n1147), .A2(G475), .ZN(n1138) );
AND2_X1 U985 ( .A1(n1318), .A2(n1147), .ZN(n1317) );
NAND2_X1 U986 ( .A1(n1319), .A2(n1211), .ZN(n1147) );
XNOR2_X1 U987 ( .A(n1320), .B(n1321), .ZN(n1211) );
XNOR2_X1 U988 ( .A(n1322), .B(n1323), .ZN(n1321) );
XOR2_X1 U989 ( .A(n1324), .B(n1325), .Z(n1323) );
AND2_X1 U990 ( .A1(n1326), .A2(G214), .ZN(n1325) );
NAND3_X1 U991 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1324) );
NAND2_X1 U992 ( .A1(KEYINPUT28), .A2(G125), .ZN(n1329) );
NAND3_X1 U993 ( .A1(n1330), .A2(n1331), .A3(n1229), .ZN(n1328) );
INV_X1 U994 ( .A(KEYINPUT28), .ZN(n1331) );
OR2_X1 U995 ( .A1(n1229), .A2(n1330), .ZN(n1327) );
NOR2_X1 U996 ( .A1(G125), .A2(KEYINPUT49), .ZN(n1330) );
XOR2_X1 U997 ( .A(n1332), .B(n1333), .Z(n1320) );
XNOR2_X1 U998 ( .A(KEYINPUT60), .B(n1160), .ZN(n1333) );
INV_X1 U999 ( .A(G131), .ZN(n1160) );
XOR2_X1 U1000 ( .A(n1334), .B(G104), .Z(n1332) );
NAND3_X1 U1001 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1002 ( .A1(KEYINPUT55), .A2(G113), .ZN(n1337) );
NAND3_X1 U1003 ( .A1(n1309), .A2(n1338), .A3(G122), .ZN(n1336) );
NAND2_X1 U1004 ( .A1(n1339), .A2(n1340), .ZN(n1335) );
INV_X1 U1005 ( .A(G122), .ZN(n1340) );
NAND2_X1 U1006 ( .A1(n1341), .A2(n1338), .ZN(n1339) );
INV_X1 U1007 ( .A(KEYINPUT55), .ZN(n1338) );
XNOR2_X1 U1008 ( .A(KEYINPUT39), .B(n1309), .ZN(n1341) );
INV_X1 U1009 ( .A(G113), .ZN(n1309) );
XNOR2_X1 U1010 ( .A(KEYINPUT37), .B(n1209), .ZN(n1319) );
XNOR2_X1 U1011 ( .A(KEYINPUT4), .B(n1214), .ZN(n1318) );
INV_X1 U1012 ( .A(G475), .ZN(n1214) );
INV_X1 U1013 ( .A(n1287), .ZN(n1112) );
XOR2_X1 U1014 ( .A(n1128), .B(KEYINPUT13), .Z(n1287) );
XOR2_X1 U1015 ( .A(n1342), .B(n1200), .Z(n1128) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1343), .ZN(n1200) );
OR2_X1 U1017 ( .A1(n1199), .A2(G902), .ZN(n1342) );
XNOR2_X1 U1018 ( .A(n1344), .B(n1345), .ZN(n1199) );
XOR2_X1 U1019 ( .A(n1346), .B(n1347), .Z(n1345) );
NAND2_X1 U1020 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1021 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
XOR2_X1 U1022 ( .A(n1167), .B(KEYINPUT51), .Z(n1350) );
NAND2_X1 U1023 ( .A1(G146), .A2(n1352), .ZN(n1348) );
XOR2_X1 U1024 ( .A(n1167), .B(KEYINPUT9), .Z(n1352) );
XNOR2_X1 U1025 ( .A(G125), .B(G140), .ZN(n1167) );
NAND2_X1 U1026 ( .A1(G221), .A2(n1353), .ZN(n1346) );
XOR2_X1 U1027 ( .A(n1354), .B(n1355), .Z(n1344) );
XNOR2_X1 U1028 ( .A(G137), .B(n1227), .ZN(n1355) );
NAND3_X1 U1029 ( .A1(n1356), .A2(n1357), .A3(n1358), .ZN(n1354) );
OR2_X1 U1030 ( .A1(n1359), .A2(G119), .ZN(n1358) );
NAND3_X1 U1031 ( .A1(G119), .A2(n1359), .A3(n1292), .ZN(n1357) );
NAND2_X1 U1032 ( .A1(G128), .A2(n1360), .ZN(n1356) );
NAND2_X1 U1033 ( .A1(n1361), .A2(n1359), .ZN(n1360) );
INV_X1 U1034 ( .A(KEYINPUT14), .ZN(n1359) );
XNOR2_X1 U1035 ( .A(G119), .B(KEYINPUT8), .ZN(n1361) );
INV_X1 U1036 ( .A(n1296), .ZN(n1094) );
XOR2_X1 U1037 ( .A(n1129), .B(KEYINPUT62), .Z(n1296) );
XNOR2_X1 U1038 ( .A(n1362), .B(G478), .ZN(n1129) );
NAND2_X1 U1039 ( .A1(n1204), .A2(n1209), .ZN(n1362) );
XNOR2_X1 U1040 ( .A(n1363), .B(n1364), .ZN(n1204) );
XNOR2_X1 U1041 ( .A(n1365), .B(n1366), .ZN(n1364) );
NAND2_X1 U1042 ( .A1(G217), .A2(n1353), .ZN(n1365) );
AND2_X1 U1043 ( .A1(G234), .A2(n1151), .ZN(n1353) );
XNOR2_X1 U1044 ( .A(n1367), .B(n1166), .ZN(n1363) );
INV_X1 U1045 ( .A(G134), .ZN(n1166) );
NAND2_X1 U1046 ( .A1(n1368), .A2(KEYINPUT57), .ZN(n1367) );
XOR2_X1 U1047 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1048 ( .A(G107), .B(G122), .ZN(n1369) );
NAND2_X1 U1049 ( .A1(n1371), .A2(n1372), .ZN(n1288) );
NAND2_X1 U1050 ( .A1(n1373), .A2(n1143), .ZN(n1372) );
NAND2_X1 U1051 ( .A1(KEYINPUT29), .A2(n1374), .ZN(n1373) );
NAND2_X1 U1052 ( .A1(KEYINPUT3), .A2(n1145), .ZN(n1374) );
INV_X1 U1053 ( .A(G472), .ZN(n1145) );
NAND2_X1 U1054 ( .A1(G472), .A2(n1375), .ZN(n1371) );
NAND2_X1 U1055 ( .A1(KEYINPUT3), .A2(n1376), .ZN(n1375) );
NAND2_X1 U1056 ( .A1(n1146), .A2(KEYINPUT29), .ZN(n1376) );
INV_X1 U1057 ( .A(n1143), .ZN(n1146) );
NAND3_X1 U1058 ( .A1(n1377), .A2(n1378), .A3(n1209), .ZN(n1143) );
NAND2_X1 U1059 ( .A1(KEYINPUT43), .A2(n1379), .ZN(n1378) );
NAND2_X1 U1060 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
NAND2_X1 U1061 ( .A1(n1219), .A2(n1382), .ZN(n1381) );
NAND2_X1 U1062 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NAND2_X1 U1063 ( .A1(KEYINPUT61), .A2(n1385), .ZN(n1384) );
NAND2_X1 U1064 ( .A1(n1386), .A2(n1387), .ZN(n1380) );
NAND2_X1 U1065 ( .A1(KEYINPUT61), .A2(n1383), .ZN(n1387) );
NAND4_X1 U1066 ( .A1(n1388), .A2(n1389), .A3(n1383), .A4(n1390), .ZN(n1377) );
INV_X1 U1067 ( .A(KEYINPUT43), .ZN(n1390) );
XNOR2_X1 U1068 ( .A(n1219), .B(KEYINPUT24), .ZN(n1383) );
NAND2_X1 U1069 ( .A1(n1385), .A2(n1391), .ZN(n1389) );
NAND2_X1 U1070 ( .A1(n1219), .A2(n1392), .ZN(n1391) );
XNOR2_X1 U1071 ( .A(n1393), .B(G101), .ZN(n1219) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1326), .ZN(n1393) );
NOR2_X1 U1073 ( .A1(G953), .A2(G237), .ZN(n1326) );
NAND2_X1 U1074 ( .A1(n1386), .A2(n1392), .ZN(n1388) );
INV_X1 U1075 ( .A(KEYINPUT61), .ZN(n1392) );
INV_X1 U1076 ( .A(n1385), .ZN(n1386) );
XOR2_X1 U1077 ( .A(n1223), .B(n1220), .Z(n1385) );
XNOR2_X1 U1078 ( .A(n1394), .B(n1395), .ZN(n1220) );
AND3_X1 U1079 ( .A1(n1115), .A2(n1301), .A3(n1104), .ZN(n1267) );
NOR2_X1 U1080 ( .A1(n1396), .A2(n1139), .ZN(n1104) );
INV_X1 U1081 ( .A(n1106), .ZN(n1139) );
NAND2_X1 U1082 ( .A1(G214), .A2(n1397), .ZN(n1106) );
INV_X1 U1083 ( .A(n1105), .ZN(n1396) );
XOR2_X1 U1084 ( .A(n1133), .B(n1136), .Z(n1105) );
NAND2_X1 U1085 ( .A1(G210), .A2(n1397), .ZN(n1136) );
NAND2_X1 U1086 ( .A1(n1398), .A2(n1209), .ZN(n1397) );
INV_X1 U1087 ( .A(G237), .ZN(n1398) );
NAND2_X1 U1088 ( .A1(n1399), .A2(n1209), .ZN(n1133) );
XNOR2_X1 U1089 ( .A(n1400), .B(n1238), .ZN(n1399) );
XNOR2_X1 U1090 ( .A(n1401), .B(n1185), .ZN(n1238) );
XNOR2_X1 U1091 ( .A(n1402), .B(n1403), .ZN(n1185) );
NAND2_X1 U1092 ( .A1(KEYINPUT17), .A2(n1404), .ZN(n1402) );
XNOR2_X1 U1093 ( .A(n1188), .B(n1405), .ZN(n1401) );
NOR2_X1 U1094 ( .A1(KEYINPUT47), .A2(n1186), .ZN(n1405) );
XNOR2_X1 U1095 ( .A(n1395), .B(KEYINPUT58), .ZN(n1186) );
XNOR2_X1 U1096 ( .A(n1406), .B(n1370), .ZN(n1395) );
XOR2_X1 U1097 ( .A(G116), .B(KEYINPUT1), .Z(n1370) );
XNOR2_X1 U1098 ( .A(G113), .B(G119), .ZN(n1406) );
XNOR2_X1 U1099 ( .A(G122), .B(n1227), .ZN(n1188) );
NAND2_X1 U1100 ( .A1(n1407), .A2(n1408), .ZN(n1400) );
NAND2_X1 U1101 ( .A1(n1273), .A2(n1409), .ZN(n1408) );
NAND2_X1 U1102 ( .A1(KEYINPUT53), .A2(n1410), .ZN(n1409) );
NAND2_X1 U1103 ( .A1(n1271), .A2(KEYINPUT53), .ZN(n1407) );
NOR2_X1 U1104 ( .A1(n1273), .A2(n1272), .ZN(n1271) );
INV_X1 U1105 ( .A(n1410), .ZN(n1272) );
NAND2_X1 U1106 ( .A1(G224), .A2(n1151), .ZN(n1410) );
XNOR2_X1 U1107 ( .A(n1223), .B(G125), .ZN(n1273) );
AND2_X1 U1108 ( .A1(n1411), .A2(n1412), .ZN(n1223) );
NAND2_X1 U1109 ( .A1(n1366), .A2(G146), .ZN(n1412) );
NAND2_X1 U1110 ( .A1(n1413), .A2(n1351), .ZN(n1411) );
XNOR2_X1 U1111 ( .A(n1366), .B(KEYINPUT42), .ZN(n1413) );
XNOR2_X1 U1112 ( .A(G143), .B(n1292), .ZN(n1366) );
INV_X1 U1113 ( .A(G128), .ZN(n1292) );
NAND2_X1 U1114 ( .A1(n1297), .A2(n1414), .ZN(n1301) );
NAND3_X1 U1115 ( .A1(G902), .A2(n1123), .A3(n1182), .ZN(n1414) );
NOR2_X1 U1116 ( .A1(n1151), .A2(G898), .ZN(n1182) );
NAND3_X1 U1117 ( .A1(n1123), .A2(n1151), .A3(G952), .ZN(n1297) );
NAND2_X1 U1118 ( .A1(G237), .A2(n1415), .ZN(n1123) );
NOR2_X1 U1119 ( .A1(n1308), .A2(n1416), .ZN(n1115) );
INV_X1 U1120 ( .A(n1117), .ZN(n1416) );
XOR2_X1 U1121 ( .A(n1417), .B(n1234), .Z(n1117) );
INV_X1 U1122 ( .A(G469), .ZN(n1234) );
NAND2_X1 U1123 ( .A1(KEYINPUT38), .A2(n1418), .ZN(n1417) );
INV_X1 U1124 ( .A(n1132), .ZN(n1418) );
NAND2_X1 U1125 ( .A1(n1419), .A2(n1209), .ZN(n1132) );
XNOR2_X1 U1126 ( .A(n1231), .B(n1420), .ZN(n1419) );
XOR2_X1 U1127 ( .A(n1421), .B(n1235), .Z(n1420) );
XOR2_X1 U1128 ( .A(n1394), .B(KEYINPUT48), .Z(n1235) );
XOR2_X1 U1129 ( .A(n1422), .B(n1423), .Z(n1394) );
XOR2_X1 U1130 ( .A(KEYINPUT10), .B(G137), .Z(n1423) );
XNOR2_X1 U1131 ( .A(G131), .B(G134), .ZN(n1422) );
NAND3_X1 U1132 ( .A1(KEYINPUT27), .A2(n1424), .A3(n1425), .ZN(n1421) );
XOR2_X1 U1133 ( .A(n1426), .B(KEYINPUT56), .Z(n1425) );
NAND2_X1 U1134 ( .A1(G110), .A2(n1229), .ZN(n1426) );
INV_X1 U1135 ( .A(G140), .ZN(n1229) );
NAND2_X1 U1136 ( .A1(G140), .A2(n1227), .ZN(n1424) );
INV_X1 U1137 ( .A(G110), .ZN(n1227) );
XNOR2_X1 U1138 ( .A(n1427), .B(n1428), .ZN(n1231) );
XOR2_X1 U1139 ( .A(n1403), .B(n1429), .Z(n1428) );
XOR2_X1 U1140 ( .A(KEYINPUT50), .B(n1430), .Z(n1429) );
AND2_X1 U1141 ( .A1(n1151), .A2(G227), .ZN(n1430) );
INV_X1 U1142 ( .A(G953), .ZN(n1151) );
XOR2_X1 U1143 ( .A(G101), .B(G107), .Z(n1403) );
XNOR2_X1 U1144 ( .A(n1169), .B(n1404), .ZN(n1427) );
XNOR2_X1 U1145 ( .A(G104), .B(KEYINPUT6), .ZN(n1404) );
XNOR2_X1 U1146 ( .A(G128), .B(n1322), .ZN(n1169) );
XNOR2_X1 U1147 ( .A(G143), .B(n1351), .ZN(n1322) );
INV_X1 U1148 ( .A(G146), .ZN(n1351) );
XOR2_X1 U1149 ( .A(n1137), .B(KEYINPUT30), .Z(n1308) );
INV_X1 U1150 ( .A(n1116), .ZN(n1137) );
NAND2_X1 U1151 ( .A1(G221), .A2(n1343), .ZN(n1116) );
NAND2_X1 U1152 ( .A1(n1415), .A2(n1209), .ZN(n1343) );
INV_X1 U1153 ( .A(G902), .ZN(n1209) );
XOR2_X1 U1154 ( .A(G234), .B(KEYINPUT0), .Z(n1415) );
endmodule


