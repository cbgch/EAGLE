//Key = 1100100100101010011100010000000011110110001110100010100000011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;

XNOR2_X1 U758 ( .A(G107), .B(n1045), .ZN(G9) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XNOR2_X1 U761 ( .A(n1052), .B(KEYINPUT39), .ZN(n1051) );
NOR4_X1 U762 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1050) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1053) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1057) );
XNOR2_X1 U766 ( .A(n1064), .B(KEYINPUT57), .ZN(n1063) );
NAND4_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1048) );
NAND4_X1 U768 ( .A1(n1064), .A2(n1062), .A3(n1069), .A4(n1070), .ZN(n1065) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
OR4_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(KEYINPUT52), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1075) );
OR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1084), .ZN(n1071) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1073), .A2(n1087), .ZN(n1086) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U779 ( .A1(n1090), .A2(n1091), .A3(KEYINPUT52), .ZN(n1089) );
NAND2_X1 U780 ( .A1(n1080), .A2(n1092), .ZN(n1085) );
NAND3_X1 U781 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NAND2_X1 U782 ( .A1(KEYINPUT55), .A2(n1096), .ZN(n1094) );
OR3_X1 U783 ( .A1(n1097), .A2(KEYINPUT55), .A3(n1096), .ZN(n1093) );
INV_X1 U784 ( .A(n1060), .ZN(n1064) );
NOR3_X1 U785 ( .A1(n1098), .A2(G953), .A3(G952), .ZN(n1046) );
INV_X1 U786 ( .A(n1067), .ZN(n1098) );
NAND4_X1 U787 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1067) );
NOR3_X1 U788 ( .A1(n1103), .A2(n1054), .A3(n1055), .ZN(n1102) );
XNOR2_X1 U789 ( .A(G478), .B(n1104), .ZN(n1103) );
XNOR2_X1 U790 ( .A(n1105), .B(n1106), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1107), .A2(KEYINPUT54), .ZN(n1106) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1099) );
XOR2_X1 U793 ( .A(n1110), .B(G472), .Z(n1109) );
XNOR2_X1 U794 ( .A(KEYINPUT56), .B(KEYINPUT33), .ZN(n1108) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(G72) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1068), .ZN(n1112) );
AND2_X1 U797 ( .A1(G227), .A2(G900), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1068), .ZN(n1115) );
XNOR2_X1 U800 ( .A(n1052), .B(n1117), .ZN(n1116) );
NAND3_X1 U801 ( .A1(G900), .A2(n1117), .A3(G953), .ZN(n1114) );
XOR2_X1 U802 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U803 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U804 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR2_X1 U805 ( .A1(KEYINPUT48), .A2(n1124), .ZN(n1123) );
NAND2_X1 U806 ( .A1(KEYINPUT18), .A2(n1125), .ZN(n1122) );
XOR2_X1 U807 ( .A(KEYINPUT32), .B(G131), .Z(n1125) );
XNOR2_X1 U808 ( .A(G125), .B(n1126), .ZN(n1118) );
XNOR2_X1 U809 ( .A(KEYINPUT42), .B(n1127), .ZN(n1126) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(G69) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND3_X1 U812 ( .A1(n1132), .A2(n1068), .A3(KEYINPUT50), .ZN(n1131) );
NAND2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U814 ( .A(n1066), .B(KEYINPUT30), .Z(n1133) );
NAND2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1136) );
XNOR2_X1 U817 ( .A(KEYINPUT58), .B(n1068), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1128) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U820 ( .A(n1141), .B(KEYINPUT60), .ZN(n1140) );
NAND2_X1 U821 ( .A1(KEYINPUT0), .A2(n1142), .ZN(n1141) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1139) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(G66) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U826 ( .A1(KEYINPUT49), .A2(n1151), .ZN(n1150) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
AND2_X1 U828 ( .A1(n1151), .A2(KEYINPUT49), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1154), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR3_X1 U831 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
XNOR2_X1 U832 ( .A(KEYINPUT8), .B(n1160), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1145), .A2(n1161), .ZN(G60) );
XOR2_X1 U834 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U835 ( .A1(n1152), .A2(G475), .ZN(n1163) );
XOR2_X1 U836 ( .A(G104), .B(n1164), .Z(G6) );
NOR2_X1 U837 ( .A1(n1088), .A2(n1165), .ZN(n1164) );
NOR2_X1 U838 ( .A1(n1145), .A2(n1166), .ZN(G57) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U840 ( .A(KEYINPUT5), .B(n1169), .Z(n1168) );
NOR2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
AND2_X1 U842 ( .A1(n1171), .A2(n1170), .ZN(n1167) );
XNOR2_X1 U843 ( .A(n1172), .B(n1173), .ZN(n1171) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U845 ( .A(n1176), .B(KEYINPUT17), .Z(n1172) );
NAND2_X1 U846 ( .A1(n1152), .A2(G472), .ZN(n1176) );
NOR3_X1 U847 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(G54) );
NOR3_X1 U848 ( .A1(n1180), .A2(G953), .A3(G952), .ZN(n1179) );
AND2_X1 U849 ( .A1(n1180), .A2(n1145), .ZN(n1178) );
INV_X1 U850 ( .A(KEYINPUT22), .ZN(n1180) );
XOR2_X1 U851 ( .A(n1181), .B(n1182), .Z(n1177) );
XOR2_X1 U852 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U853 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U854 ( .A1(KEYINPUT36), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U855 ( .A(n1188), .B(n1127), .ZN(n1187) );
NAND2_X1 U856 ( .A1(KEYINPUT7), .A2(n1189), .ZN(n1188) );
NAND2_X1 U857 ( .A1(n1152), .A2(G469), .ZN(n1183) );
XNOR2_X1 U858 ( .A(n1190), .B(n1191), .ZN(n1181) );
NOR2_X1 U859 ( .A1(n1145), .A2(n1192), .ZN(G51) );
XOR2_X1 U860 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND2_X1 U861 ( .A1(n1152), .A2(n1195), .ZN(n1193) );
AND2_X1 U862 ( .A1(G902), .A2(n1160), .ZN(n1152) );
NAND3_X1 U863 ( .A1(n1052), .A2(n1066), .A3(n1134), .ZN(n1160) );
INV_X1 U864 ( .A(n1049), .ZN(n1134) );
NAND4_X1 U865 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1049) );
AND3_X1 U866 ( .A1(n1200), .A2(n1045), .A3(n1201), .ZN(n1199) );
NAND4_X1 U867 ( .A1(n1083), .A2(n1062), .A3(n1202), .A4(n1203), .ZN(n1045) );
OR2_X1 U868 ( .A1(n1204), .A2(KEYINPUT40), .ZN(n1198) );
NAND3_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1069), .ZN(n1197) );
NAND2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U871 ( .A1(n1062), .A2(n1209), .ZN(n1205) );
NAND4_X1 U872 ( .A1(n1210), .A2(n1088), .A3(n1211), .A4(n1212), .ZN(n1209) );
AND3_X1 U873 ( .A1(KEYINPUT40), .A2(n1073), .A3(n1213), .ZN(n1212) );
NAND2_X1 U874 ( .A1(n1214), .A2(n1215), .ZN(n1196) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U876 ( .A(KEYINPUT10), .B(n1165), .ZN(n1217) );
NAND4_X1 U877 ( .A1(n1082), .A2(n1062), .A3(n1203), .A4(n1210), .ZN(n1165) );
XOR2_X1 U878 ( .A(n1218), .B(KEYINPUT24), .Z(n1216) );
NAND2_X1 U879 ( .A1(n1219), .A2(n1220), .ZN(n1066) );
XNOR2_X1 U880 ( .A(KEYINPUT16), .B(n1059), .ZN(n1220) );
INV_X1 U881 ( .A(n1207), .ZN(n1219) );
AND4_X1 U882 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1052) );
NOR4_X1 U883 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
INV_X1 U884 ( .A(n1229), .ZN(n1228) );
NOR2_X1 U885 ( .A1(n1230), .A2(n1231), .ZN(n1223) );
INV_X1 U886 ( .A(n1232), .ZN(n1231) );
NAND3_X1 U887 ( .A1(n1082), .A2(n1214), .A3(n1233), .ZN(n1222) );
NAND2_X1 U888 ( .A1(n1080), .A2(n1234), .ZN(n1221) );
XOR2_X1 U889 ( .A(KEYINPUT20), .B(n1235), .Z(n1234) );
NOR2_X1 U890 ( .A1(n1068), .A2(G952), .ZN(n1145) );
XOR2_X1 U891 ( .A(G146), .B(n1236), .Z(G48) );
NOR3_X1 U892 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
XNOR2_X1 U893 ( .A(n1214), .B(KEYINPUT28), .ZN(n1238) );
XNOR2_X1 U894 ( .A(G143), .B(n1240), .ZN(G45) );
NAND2_X1 U895 ( .A1(KEYINPUT1), .A2(n1227), .ZN(n1240) );
AND4_X1 U896 ( .A1(n1241), .A2(n1214), .A3(n1213), .A4(n1211), .ZN(n1227) );
XNOR2_X1 U897 ( .A(G140), .B(n1232), .ZN(G42) );
NAND3_X1 U898 ( .A1(n1069), .A2(n1208), .A3(n1242), .ZN(n1232) );
XOR2_X1 U899 ( .A(G137), .B(n1226), .Z(G39) );
NOR3_X1 U900 ( .A1(n1056), .A2(n1054), .A3(n1237), .ZN(n1226) );
INV_X1 U901 ( .A(n1079), .ZN(n1056) );
XNOR2_X1 U902 ( .A(G134), .B(n1243), .ZN(G36) );
NAND2_X1 U903 ( .A1(n1235), .A2(n1080), .ZN(n1243) );
AND2_X1 U904 ( .A1(n1241), .A2(n1083), .ZN(n1235) );
NOR3_X1 U905 ( .A1(n1095), .A2(n1244), .A3(n1059), .ZN(n1241) );
XOR2_X1 U906 ( .A(G131), .B(n1230), .Z(G33) );
AND2_X1 U907 ( .A1(n1242), .A2(n1245), .ZN(n1230) );
NOR4_X1 U908 ( .A1(n1239), .A2(n1054), .A3(n1095), .A4(n1244), .ZN(n1242) );
INV_X1 U909 ( .A(n1080), .ZN(n1054) );
NOR2_X1 U910 ( .A1(n1077), .A2(n1091), .ZN(n1080) );
INV_X1 U911 ( .A(n1082), .ZN(n1239) );
XOR2_X1 U912 ( .A(G128), .B(n1225), .Z(G30) );
AND3_X1 U913 ( .A1(n1083), .A2(n1214), .A3(n1233), .ZN(n1225) );
INV_X1 U914 ( .A(n1237), .ZN(n1233) );
NAND4_X1 U915 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1208), .ZN(n1237) );
XOR2_X1 U916 ( .A(G101), .B(n1249), .Z(G3) );
NOR2_X1 U917 ( .A1(n1059), .A2(n1207), .ZN(n1249) );
NAND3_X1 U918 ( .A1(n1202), .A2(n1246), .A3(n1079), .ZN(n1207) );
INV_X1 U919 ( .A(n1095), .ZN(n1246) );
INV_X1 U920 ( .A(n1245), .ZN(n1059) );
XNOR2_X1 U921 ( .A(G125), .B(n1229), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1073), .A2(n1069), .A3(n1082), .A4(n1250), .ZN(n1229) );
NOR3_X1 U923 ( .A1(n1088), .A2(n1062), .A3(n1244), .ZN(n1250) );
INV_X1 U924 ( .A(n1248), .ZN(n1244) );
NAND2_X1 U925 ( .A1(n1060), .A2(n1251), .ZN(n1248) );
NAND4_X1 U926 ( .A1(G953), .A2(G902), .A3(n1252), .A4(n1253), .ZN(n1251) );
INV_X1 U927 ( .A(G900), .ZN(n1253) );
XNOR2_X1 U928 ( .A(G122), .B(n1204), .ZN(G24) );
NAND3_X1 U929 ( .A1(n1254), .A2(n1062), .A3(n1255), .ZN(n1204) );
NOR3_X1 U930 ( .A1(n1061), .A2(n1101), .A3(n1256), .ZN(n1255) );
XNOR2_X1 U931 ( .A(G119), .B(n1200), .ZN(G21) );
NAND4_X1 U932 ( .A1(n1254), .A2(n1079), .A3(n1247), .A4(n1208), .ZN(n1200) );
XNOR2_X1 U933 ( .A(n1061), .B(KEYINPUT59), .ZN(n1247) );
NAND2_X1 U934 ( .A1(n1257), .A2(n1258), .ZN(G18) );
NAND2_X1 U935 ( .A1(G116), .A2(n1201), .ZN(n1258) );
XOR2_X1 U936 ( .A(KEYINPUT38), .B(n1259), .Z(n1257) );
NOR2_X1 U937 ( .A1(G116), .A2(n1201), .ZN(n1259) );
NAND3_X1 U938 ( .A1(n1245), .A2(n1083), .A3(n1254), .ZN(n1201) );
AND2_X1 U939 ( .A1(n1073), .A2(n1202), .ZN(n1254) );
NOR2_X1 U940 ( .A1(n1088), .A2(n1260), .ZN(n1202) );
NOR2_X1 U941 ( .A1(n1211), .A2(n1256), .ZN(n1083) );
XNOR2_X1 U942 ( .A(n1261), .B(n1262), .ZN(G15) );
NOR2_X1 U943 ( .A1(n1088), .A2(n1218), .ZN(n1262) );
NAND4_X1 U944 ( .A1(n1082), .A2(n1245), .A3(n1073), .A4(n1210), .ZN(n1218) );
INV_X1 U945 ( .A(n1055), .ZN(n1073) );
NAND2_X1 U946 ( .A1(n1263), .A2(n1096), .ZN(n1055) );
INV_X1 U947 ( .A(n1097), .ZN(n1263) );
NOR2_X1 U948 ( .A1(n1208), .A2(n1069), .ZN(n1245) );
INV_X1 U949 ( .A(n1061), .ZN(n1069) );
NOR2_X1 U950 ( .A1(n1213), .A2(n1101), .ZN(n1082) );
INV_X1 U951 ( .A(n1211), .ZN(n1101) );
INV_X1 U952 ( .A(n1214), .ZN(n1088) );
XNOR2_X1 U953 ( .A(G110), .B(n1264), .ZN(G12) );
NAND3_X1 U954 ( .A1(n1079), .A2(n1203), .A3(n1265), .ZN(n1264) );
NOR3_X1 U955 ( .A1(n1266), .A2(n1062), .A3(n1260), .ZN(n1265) );
INV_X1 U956 ( .A(n1210), .ZN(n1260) );
NAND2_X1 U957 ( .A1(n1060), .A2(n1267), .ZN(n1210) );
NAND3_X1 U958 ( .A1(G902), .A2(n1252), .A3(n1137), .ZN(n1267) );
NOR2_X1 U959 ( .A1(n1068), .A2(G898), .ZN(n1137) );
NAND3_X1 U960 ( .A1(n1252), .A2(n1068), .A3(G952), .ZN(n1060) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1252) );
INV_X1 U962 ( .A(n1208), .ZN(n1062) );
NAND2_X1 U963 ( .A1(n1268), .A2(n1269), .ZN(n1208) );
OR2_X1 U964 ( .A1(n1270), .A2(n1107), .ZN(n1269) );
XOR2_X1 U965 ( .A(n1271), .B(KEYINPUT25), .Z(n1268) );
NAND2_X1 U966 ( .A1(n1107), .A2(n1270), .ZN(n1271) );
XOR2_X1 U967 ( .A(n1153), .B(KEYINPUT23), .Z(n1270) );
INV_X1 U968 ( .A(n1105), .ZN(n1153) );
NAND2_X1 U969 ( .A1(G217), .A2(n1272), .ZN(n1105) );
AND2_X1 U970 ( .A1(n1273), .A2(n1151), .ZN(n1107) );
XNOR2_X1 U971 ( .A(n1274), .B(n1275), .ZN(n1151) );
XOR2_X1 U972 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U973 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U974 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR2_X1 U975 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NOR2_X1 U976 ( .A1(KEYINPUT27), .A2(n1284), .ZN(n1282) );
NOR2_X1 U977 ( .A1(KEYINPUT29), .A2(n1127), .ZN(n1284) );
NOR2_X1 U978 ( .A1(G140), .A2(n1285), .ZN(n1280) );
NOR2_X1 U979 ( .A1(n1286), .A2(KEYINPUT29), .ZN(n1285) );
NOR2_X1 U980 ( .A1(KEYINPUT27), .A2(G125), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1287), .A2(n1288), .ZN(n1278) );
NAND2_X1 U982 ( .A1(G110), .A2(n1289), .ZN(n1288) );
XOR2_X1 U983 ( .A(KEYINPUT37), .B(n1290), .Z(n1287) );
NOR2_X1 U984 ( .A1(G110), .A2(n1289), .ZN(n1290) );
XNOR2_X1 U985 ( .A(G128), .B(n1291), .ZN(n1289) );
NOR2_X1 U986 ( .A1(G119), .A2(KEYINPUT2), .ZN(n1291) );
NAND2_X1 U987 ( .A1(G221), .A2(n1292), .ZN(n1276) );
XNOR2_X1 U988 ( .A(G137), .B(n1293), .ZN(n1274) );
XOR2_X1 U989 ( .A(KEYINPUT53), .B(G146), .Z(n1293) );
XNOR2_X1 U990 ( .A(n1214), .B(KEYINPUT13), .ZN(n1266) );
NOR2_X1 U991 ( .A1(n1090), .A2(n1091), .ZN(n1214) );
INV_X1 U992 ( .A(n1078), .ZN(n1091) );
NAND2_X1 U993 ( .A1(G214), .A2(n1294), .ZN(n1078) );
INV_X1 U994 ( .A(n1077), .ZN(n1090) );
XNOR2_X1 U995 ( .A(n1295), .B(n1195), .ZN(n1077) );
AND2_X1 U996 ( .A1(G210), .A2(n1294), .ZN(n1195) );
NAND2_X1 U997 ( .A1(n1296), .A2(n1158), .ZN(n1294) );
INV_X1 U998 ( .A(G237), .ZN(n1296) );
NAND2_X1 U999 ( .A1(n1273), .A2(n1194), .ZN(n1295) );
XNOR2_X1 U1000 ( .A(n1297), .B(n1298), .ZN(n1194) );
XOR2_X1 U1001 ( .A(n1143), .B(n1142), .Z(n1298) );
XOR2_X1 U1002 ( .A(n1299), .B(n1300), .Z(n1142) );
XOR2_X1 U1003 ( .A(G119), .B(n1301), .Z(n1300) );
NOR2_X1 U1004 ( .A1(KEYINPUT47), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U1005 ( .A(G116), .B(KEYINPUT62), .ZN(n1302) );
NAND2_X1 U1006 ( .A1(KEYINPUT61), .A2(n1261), .ZN(n1299) );
XNOR2_X1 U1007 ( .A(G110), .B(n1303), .ZN(n1143) );
XNOR2_X1 U1008 ( .A(KEYINPUT4), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1009 ( .A(n1190), .B(n1305), .ZN(n1297) );
XNOR2_X1 U1010 ( .A(n1283), .B(n1306), .ZN(n1305) );
AND2_X1 U1011 ( .A1(n1068), .A2(G224), .ZN(n1306) );
NOR2_X1 U1012 ( .A1(n1061), .A2(n1095), .ZN(n1203) );
NAND2_X1 U1013 ( .A1(n1097), .A2(n1096), .ZN(n1095) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1272), .ZN(n1096) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1158), .ZN(n1272) );
INV_X1 U1016 ( .A(G902), .ZN(n1158) );
XNOR2_X1 U1017 ( .A(n1307), .B(G469), .ZN(n1097) );
NAND2_X1 U1018 ( .A1(n1308), .A2(n1273), .ZN(n1307) );
XOR2_X1 U1019 ( .A(n1309), .B(n1191), .Z(n1308) );
XNOR2_X1 U1020 ( .A(n1310), .B(n1311), .ZN(n1309) );
NAND2_X1 U1021 ( .A1(KEYINPUT44), .A2(n1190), .ZN(n1311) );
XOR2_X1 U1022 ( .A(n1144), .B(n1124), .Z(n1190) );
XOR2_X1 U1023 ( .A(G101), .B(n1312), .Z(n1144) );
XNOR2_X1 U1024 ( .A(n1313), .B(G104), .ZN(n1312) );
INV_X1 U1025 ( .A(G107), .ZN(n1313) );
NAND3_X1 U1026 ( .A1(n1314), .A2(n1315), .A3(KEYINPUT34), .ZN(n1310) );
NAND2_X1 U1027 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
INV_X1 U1028 ( .A(KEYINPUT31), .ZN(n1317) );
XOR2_X1 U1029 ( .A(n1185), .B(n1318), .Z(n1316) );
NAND3_X1 U1030 ( .A1(n1318), .A2(n1185), .A3(KEYINPUT31), .ZN(n1314) );
NAND2_X1 U1031 ( .A1(G227), .A2(n1068), .ZN(n1185) );
XNOR2_X1 U1032 ( .A(n1189), .B(G140), .ZN(n1318) );
INV_X1 U1033 ( .A(G110), .ZN(n1189) );
NAND2_X1 U1034 ( .A1(n1319), .A2(n1320), .ZN(n1061) );
NAND2_X1 U1035 ( .A1(G472), .A2(n1110), .ZN(n1320) );
XOR2_X1 U1036 ( .A(KEYINPUT35), .B(n1321), .Z(n1319) );
NOR2_X1 U1037 ( .A1(G472), .A2(n1110), .ZN(n1321) );
NAND2_X1 U1038 ( .A1(n1273), .A2(n1322), .ZN(n1110) );
XOR2_X1 U1039 ( .A(n1323), .B(n1170), .Z(n1322) );
XOR2_X1 U1040 ( .A(n1324), .B(G101), .Z(n1170) );
NAND2_X1 U1041 ( .A1(G210), .A2(n1325), .ZN(n1324) );
NAND3_X1 U1042 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1323) );
NAND2_X1 U1043 ( .A1(n1329), .A2(n1174), .ZN(n1328) );
NAND2_X1 U1044 ( .A1(KEYINPUT11), .A2(n1330), .ZN(n1327) );
NAND2_X1 U1045 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XNOR2_X1 U1046 ( .A(KEYINPUT9), .B(n1174), .ZN(n1331) );
NAND2_X1 U1047 ( .A1(n1333), .A2(n1334), .ZN(n1326) );
INV_X1 U1048 ( .A(KEYINPUT11), .ZN(n1334) );
NAND2_X1 U1049 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
OR3_X1 U1050 ( .A1(n1329), .A2(n1174), .A3(KEYINPUT9), .ZN(n1336) );
INV_X1 U1051 ( .A(n1332), .ZN(n1329) );
XOR2_X1 U1052 ( .A(n1175), .B(n1337), .Z(n1332) );
XOR2_X1 U1053 ( .A(KEYINPUT41), .B(KEYINPUT26), .Z(n1337) );
XOR2_X1 U1054 ( .A(n1191), .B(n1124), .Z(n1175) );
XNOR2_X1 U1055 ( .A(n1338), .B(n1339), .ZN(n1124) );
XOR2_X1 U1056 ( .A(KEYINPUT19), .B(G128), .Z(n1339) );
XOR2_X1 U1057 ( .A(G131), .B(n1120), .Z(n1191) );
XOR2_X1 U1058 ( .A(G134), .B(G137), .Z(n1120) );
NAND2_X1 U1059 ( .A1(KEYINPUT9), .A2(n1174), .ZN(n1335) );
XOR2_X1 U1060 ( .A(n1340), .B(n1261), .Z(n1174) );
NAND2_X1 U1061 ( .A1(KEYINPUT43), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1062 ( .A(G119), .B(G116), .Z(n1341) );
NOR2_X1 U1063 ( .A1(n1211), .A2(n1213), .ZN(n1079) );
INV_X1 U1064 ( .A(n1256), .ZN(n1213) );
XOR2_X1 U1065 ( .A(n1342), .B(n1104), .Z(n1256) );
NAND2_X1 U1066 ( .A1(n1156), .A2(n1273), .ZN(n1104) );
XOR2_X1 U1067 ( .A(n1343), .B(n1344), .Z(n1156) );
XOR2_X1 U1068 ( .A(G134), .B(n1345), .Z(n1344) );
NOR2_X1 U1069 ( .A1(KEYINPUT15), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1070 ( .A(G128), .B(n1347), .ZN(n1346) );
XOR2_X1 U1071 ( .A(n1348), .B(n1349), .Z(n1343) );
AND2_X1 U1072 ( .A1(n1292), .A2(G217), .ZN(n1349) );
AND2_X1 U1073 ( .A1(G234), .A2(n1068), .ZN(n1292) );
INV_X1 U1074 ( .A(G953), .ZN(n1068) );
NAND2_X1 U1075 ( .A1(KEYINPUT63), .A2(n1350), .ZN(n1348) );
XNOR2_X1 U1076 ( .A(G107), .B(n1351), .ZN(n1350) );
NAND2_X1 U1077 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1078 ( .A1(G116), .A2(n1304), .ZN(n1353) );
XOR2_X1 U1079 ( .A(n1354), .B(KEYINPUT6), .Z(n1352) );
OR2_X1 U1080 ( .A1(n1304), .A2(G116), .ZN(n1354) );
INV_X1 U1081 ( .A(G122), .ZN(n1304) );
NAND2_X1 U1082 ( .A1(KEYINPUT12), .A2(n1159), .ZN(n1342) );
INV_X1 U1083 ( .A(G478), .ZN(n1159) );
XOR2_X1 U1084 ( .A(G475), .B(n1355), .Z(n1211) );
AND2_X1 U1085 ( .A1(n1162), .A2(n1273), .ZN(n1355) );
XNOR2_X1 U1086 ( .A(G902), .B(KEYINPUT21), .ZN(n1273) );
NAND2_X1 U1087 ( .A1(n1356), .A2(n1357), .ZN(n1162) );
NAND2_X1 U1088 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1089 ( .A(KEYINPUT14), .B(n1360), .Z(n1356) );
NOR2_X1 U1090 ( .A1(n1358), .A2(n1359), .ZN(n1360) );
XNOR2_X1 U1091 ( .A(n1361), .B(n1362), .ZN(n1359) );
XNOR2_X1 U1092 ( .A(G131), .B(n1363), .ZN(n1362) );
NAND2_X1 U1093 ( .A1(G214), .A2(n1325), .ZN(n1363) );
NOR2_X1 U1094 ( .A1(G953), .A2(G237), .ZN(n1325) );
XNOR2_X1 U1095 ( .A(n1364), .B(n1338), .ZN(n1361) );
XNOR2_X1 U1096 ( .A(G146), .B(n1347), .ZN(n1338) );
XOR2_X1 U1097 ( .A(G143), .B(KEYINPUT45), .Z(n1347) );
NAND3_X1 U1098 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1364) );
NAND2_X1 U1099 ( .A1(KEYINPUT3), .A2(G125), .ZN(n1367) );
NAND3_X1 U1100 ( .A1(n1283), .A2(n1368), .A3(G140), .ZN(n1366) );
NAND2_X1 U1101 ( .A1(n1369), .A2(n1127), .ZN(n1365) );
INV_X1 U1102 ( .A(G140), .ZN(n1127) );
NAND2_X1 U1103 ( .A1(n1370), .A2(n1368), .ZN(n1369) );
INV_X1 U1104 ( .A(KEYINPUT3), .ZN(n1368) );
XNOR2_X1 U1105 ( .A(KEYINPUT46), .B(n1283), .ZN(n1370) );
INV_X1 U1106 ( .A(G125), .ZN(n1283) );
XOR2_X1 U1107 ( .A(n1371), .B(n1372), .Z(n1358) );
XNOR2_X1 U1108 ( .A(n1261), .B(G122), .ZN(n1372) );
INV_X1 U1109 ( .A(G113), .ZN(n1261) );
OR2_X1 U1110 ( .A1(G104), .A2(KEYINPUT51), .ZN(n1371) );
endmodule


