//Key = 1010100111110000100100011010101111111000010010100011010001000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372;

NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(G9) );
OR2_X1 U758 ( .A1(n1050), .A2(G107), .ZN(n1049) );
XOR2_X1 U759 ( .A(n1051), .B(KEYINPUT55), .Z(n1048) );
NAND2_X1 U760 ( .A1(G107), .A2(n1050), .ZN(n1051) );
NOR2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
XNOR2_X1 U763 ( .A(n1058), .B(KEYINPUT1), .ZN(n1057) );
NOR3_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1056) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR3_X1 U771 ( .A1(n1069), .A2(n1074), .A3(n1071), .ZN(n1062) );
INV_X1 U772 ( .A(n1075), .ZN(n1071) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
XOR2_X1 U776 ( .A(KEYINPUT25), .B(n1082), .Z(n1081) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1076) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
AND2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
INV_X1 U781 ( .A(n1091), .ZN(n1069) );
INV_X1 U782 ( .A(KEYINPUT50), .ZN(n1059) );
NAND3_X1 U783 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1054) );
NAND3_X1 U784 ( .A1(n1095), .A2(n1091), .A3(n1096), .ZN(n1094) );
NOR3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1100), .B(KEYINPUT22), .Z(n1098) );
NAND2_X1 U787 ( .A1(KEYINPUT50), .A2(n1101), .ZN(n1100) );
AND2_X1 U788 ( .A1(n1092), .A2(n1102), .ZN(n1052) );
NAND4_X1 U789 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1092) );
NOR4_X1 U790 ( .A1(n1107), .A2(n1108), .A3(n1084), .A4(n1109), .ZN(n1106) );
XNOR2_X1 U791 ( .A(G478), .B(n1110), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1107) );
NOR2_X1 U793 ( .A1(KEYINPUT12), .A2(n1113), .ZN(n1112) );
XNOR2_X1 U794 ( .A(G472), .B(KEYINPUT10), .ZN(n1113) );
AND2_X1 U795 ( .A1(n1114), .A2(n1099), .ZN(n1105) );
XNOR2_X1 U796 ( .A(G469), .B(n1115), .ZN(n1104) );
NAND2_X1 U797 ( .A1(KEYINPUT4), .A2(n1116), .ZN(n1115) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1103) );
XNOR2_X1 U799 ( .A(n1119), .B(KEYINPUT0), .ZN(n1118) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(G72) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1093), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
NAND2_X1 U804 ( .A1(n1127), .A2(n1093), .ZN(n1126) );
XOR2_X1 U805 ( .A(n1055), .B(n1128), .Z(n1127) );
NAND3_X1 U806 ( .A1(G900), .A2(n1128), .A3(G953), .ZN(n1125) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U808 ( .A(KEYINPUT20), .B(G140), .Z(n1130) );
XOR2_X1 U809 ( .A(n1131), .B(n1132), .Z(n1129) );
NOR2_X1 U810 ( .A1(KEYINPUT13), .A2(n1133), .ZN(n1132) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(G69) );
NOR2_X1 U812 ( .A1(KEYINPUT17), .A2(n1136), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U814 ( .A1(n1058), .A2(G953), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U817 ( .A1(G898), .A2(n1093), .ZN(n1139) );
NAND2_X1 U818 ( .A1(G953), .A2(n1143), .ZN(n1134) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1143) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U821 ( .A(n1146), .B(n1147), .Z(n1144) );
NOR2_X1 U822 ( .A1(KEYINPUT62), .A2(n1148), .ZN(n1147) );
NAND2_X1 U823 ( .A1(n1149), .A2(G217), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(G63) );
XOR2_X1 U825 ( .A(n1145), .B(KEYINPUT59), .Z(n1151) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1150) );
NOR2_X1 U827 ( .A1(KEYINPUT27), .A2(n1154), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
INV_X1 U829 ( .A(n1157), .ZN(n1156) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1155) );
NAND2_X1 U831 ( .A1(n1149), .A2(G478), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1160), .A2(n1145), .ZN(G60) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U834 ( .A1(n1149), .A2(G475), .ZN(n1161) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(G6) );
NAND3_X1 U836 ( .A1(n1165), .A2(n1166), .A3(n1073), .ZN(n1164) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1145), .ZN(G57) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(KEYINPUT11), .Z(n1169) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
XNOR2_X1 U842 ( .A(n1173), .B(n1174), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U844 ( .A1(KEYINPUT61), .A2(n1177), .ZN(n1176) );
NAND2_X1 U845 ( .A1(n1149), .A2(G472), .ZN(n1175) );
XNOR2_X1 U846 ( .A(n1178), .B(n1179), .ZN(n1173) );
NOR2_X1 U847 ( .A1(n1180), .A2(n1145), .ZN(G54) );
XOR2_X1 U848 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U849 ( .A1(KEYINPUT56), .A2(n1183), .ZN(n1182) );
XOR2_X1 U850 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U851 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U852 ( .A(n1188), .B(n1189), .ZN(n1187) );
NOR2_X1 U853 ( .A1(G110), .A2(KEYINPUT60), .ZN(n1189) );
NAND2_X1 U854 ( .A1(KEYINPUT26), .A2(n1190), .ZN(n1188) );
XOR2_X1 U855 ( .A(KEYINPUT3), .B(n1177), .Z(n1190) );
XOR2_X1 U856 ( .A(n1191), .B(n1192), .Z(n1184) );
XOR2_X1 U857 ( .A(KEYINPUT38), .B(G140), .Z(n1192) );
NAND2_X1 U858 ( .A1(n1149), .A2(G469), .ZN(n1181) );
NOR2_X1 U859 ( .A1(n1145), .A2(n1193), .ZN(G51) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U862 ( .A1(n1149), .A2(n1119), .ZN(n1197) );
AND2_X1 U863 ( .A1(G902), .A2(n1198), .ZN(n1149) );
NAND2_X1 U864 ( .A1(n1199), .A2(n1058), .ZN(n1198) );
AND4_X1 U865 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1058) );
AND3_X1 U866 ( .A1(n1204), .A2(n1205), .A3(n1050), .ZN(n1203) );
NAND3_X1 U867 ( .A1(n1072), .A2(n1166), .A3(n1165), .ZN(n1050) );
NAND2_X1 U868 ( .A1(n1206), .A2(n1207), .ZN(n1202) );
NAND2_X1 U869 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND3_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1073), .ZN(n1200) );
NAND2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND3_X1 U872 ( .A1(n1214), .A2(n1215), .A3(n1083), .ZN(n1213) );
NAND2_X1 U873 ( .A1(KEYINPUT36), .A2(n1216), .ZN(n1215) );
NAND2_X1 U874 ( .A1(n1217), .A2(n1218), .ZN(n1214) );
INV_X1 U875 ( .A(KEYINPUT36), .ZN(n1218) );
NAND3_X1 U876 ( .A1(n1219), .A2(n1068), .A3(n1088), .ZN(n1217) );
NAND2_X1 U877 ( .A1(n1220), .A2(n1206), .ZN(n1212) );
INV_X1 U878 ( .A(n1055), .ZN(n1199) );
NAND4_X1 U879 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1055) );
NOR4_X1 U880 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NOR2_X1 U881 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
NOR2_X1 U882 ( .A1(n1068), .A2(n1231), .ZN(n1230) );
XOR2_X1 U883 ( .A(KEYINPUT24), .B(n1232), .Z(n1231) );
XNOR2_X1 U884 ( .A(n1233), .B(n1234), .ZN(n1194) );
NAND2_X1 U885 ( .A1(n1235), .A2(n1236), .ZN(n1145) );
OR3_X1 U886 ( .A1(n1093), .A2(G952), .A3(KEYINPUT58), .ZN(n1236) );
NAND2_X1 U887 ( .A1(KEYINPUT58), .A2(n1102), .ZN(n1235) );
XOR2_X1 U888 ( .A(G146), .B(n1229), .Z(G48) );
AND3_X1 U889 ( .A1(n1206), .A2(n1237), .A3(n1073), .ZN(n1229) );
XOR2_X1 U890 ( .A(n1238), .B(n1239), .Z(G45) );
NAND2_X1 U891 ( .A1(n1232), .A2(n1206), .ZN(n1239) );
AND3_X1 U892 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1232) );
XNOR2_X1 U893 ( .A(G140), .B(n1221), .ZN(G42) );
NAND3_X1 U894 ( .A1(n1075), .A2(n1088), .A3(n1243), .ZN(n1221) );
XOR2_X1 U895 ( .A(G137), .B(n1228), .Z(G39) );
AND3_X1 U896 ( .A1(n1075), .A2(n1237), .A3(n1091), .ZN(n1228) );
XOR2_X1 U897 ( .A(G134), .B(n1227), .Z(G36) );
AND3_X1 U898 ( .A1(n1241), .A2(n1072), .A3(n1075), .ZN(n1227) );
XOR2_X1 U899 ( .A(G131), .B(n1226), .Z(G33) );
AND3_X1 U900 ( .A1(n1075), .A2(n1241), .A3(n1073), .ZN(n1226) );
NOR2_X1 U901 ( .A1(n1244), .A2(n1097), .ZN(n1075) );
XNOR2_X1 U902 ( .A(KEYINPUT18), .B(n1099), .ZN(n1244) );
XNOR2_X1 U903 ( .A(n1225), .B(n1245), .ZN(G30) );
NAND2_X1 U904 ( .A1(KEYINPUT57), .A2(G128), .ZN(n1245) );
AND3_X1 U905 ( .A1(n1206), .A2(n1237), .A3(n1072), .ZN(n1225) );
NAND2_X1 U906 ( .A1(n1246), .A2(n1247), .ZN(n1237) );
NAND4_X1 U907 ( .A1(n1088), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1247) );
INV_X1 U908 ( .A(KEYINPUT29), .ZN(n1250) );
NOR2_X1 U909 ( .A1(n1210), .A2(n1083), .ZN(n1249) );
NAND2_X1 U910 ( .A1(KEYINPUT29), .A2(n1241), .ZN(n1246) );
AND4_X1 U911 ( .A1(n1210), .A2(n1088), .A3(n1248), .A4(n1251), .ZN(n1241) );
XNOR2_X1 U912 ( .A(G101), .B(n1201), .ZN(G3) );
NAND4_X1 U913 ( .A1(n1091), .A2(n1165), .A3(n1210), .A4(n1251), .ZN(n1201) );
XOR2_X1 U914 ( .A(n1133), .B(n1252), .Z(G27) );
NAND2_X1 U915 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U916 ( .A1(KEYINPUT9), .A2(n1222), .ZN(n1254) );
NAND2_X1 U917 ( .A1(KEYINPUT40), .A2(n1255), .ZN(n1253) );
INV_X1 U918 ( .A(n1222), .ZN(n1255) );
NAND3_X1 U919 ( .A1(n1243), .A2(n1206), .A3(n1256), .ZN(n1222) );
AND3_X1 U920 ( .A1(n1073), .A2(n1248), .A3(n1082), .ZN(n1243) );
NAND2_X1 U921 ( .A1(n1257), .A2(n1258), .ZN(n1248) );
NAND3_X1 U922 ( .A1(G952), .A2(n1101), .A3(n1093), .ZN(n1258) );
NAND4_X1 U923 ( .A1(n1259), .A2(n1124), .A3(G902), .A4(G953), .ZN(n1257) );
INV_X1 U924 ( .A(G900), .ZN(n1124) );
XOR2_X1 U925 ( .A(n1101), .B(KEYINPUT42), .Z(n1259) );
XOR2_X1 U926 ( .A(n1260), .B(n1261), .Z(G24) );
NAND2_X1 U927 ( .A1(n1262), .A2(n1206), .ZN(n1261) );
XOR2_X1 U928 ( .A(n1209), .B(KEYINPUT30), .Z(n1262) );
NAND4_X1 U929 ( .A1(n1242), .A2(n1095), .A3(n1240), .A4(n1219), .ZN(n1209) );
INV_X1 U930 ( .A(n1065), .ZN(n1095) );
NAND2_X1 U931 ( .A1(n1256), .A2(n1166), .ZN(n1065) );
INV_X1 U932 ( .A(n1086), .ZN(n1166) );
NAND2_X1 U933 ( .A1(n1210), .A2(n1083), .ZN(n1086) );
XOR2_X1 U934 ( .A(n1263), .B(n1204), .Z(G21) );
NAND4_X1 U935 ( .A1(n1264), .A2(n1220), .A3(n1091), .A4(n1206), .ZN(n1204) );
XOR2_X1 U936 ( .A(n1084), .B(KEYINPUT29), .Z(n1264) );
XOR2_X1 U937 ( .A(n1265), .B(n1266), .Z(G18) );
NOR2_X1 U938 ( .A1(n1068), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U939 ( .A(KEYINPUT44), .B(n1208), .ZN(n1267) );
NAND3_X1 U940 ( .A1(n1072), .A2(n1210), .A3(n1220), .ZN(n1208) );
AND2_X1 U941 ( .A1(n1240), .A2(n1268), .ZN(n1072) );
NAND2_X1 U942 ( .A1(KEYINPUT31), .A2(n1269), .ZN(n1265) );
XNOR2_X1 U943 ( .A(G113), .B(n1270), .ZN(G15) );
NAND3_X1 U944 ( .A1(n1220), .A2(n1073), .A3(n1271), .ZN(n1270) );
NOR3_X1 U945 ( .A1(n1084), .A2(KEYINPUT47), .A3(n1068), .ZN(n1271) );
NOR2_X1 U946 ( .A1(n1268), .A2(n1240), .ZN(n1073) );
INV_X1 U947 ( .A(n1242), .ZN(n1268) );
AND3_X1 U948 ( .A1(n1219), .A2(n1251), .A3(n1256), .ZN(n1220) );
INV_X1 U949 ( .A(n1079), .ZN(n1256) );
NAND2_X1 U950 ( .A1(n1089), .A2(n1114), .ZN(n1079) );
XNOR2_X1 U951 ( .A(G110), .B(n1205), .ZN(G12) );
NAND3_X1 U952 ( .A1(n1091), .A2(n1165), .A3(n1082), .ZN(n1205) );
NOR2_X1 U953 ( .A1(n1251), .A2(n1210), .ZN(n1082) );
INV_X1 U954 ( .A(n1084), .ZN(n1210) );
NAND3_X1 U955 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1084) );
NAND2_X1 U956 ( .A1(n1275), .A2(n1148), .ZN(n1274) );
OR3_X1 U957 ( .A1(n1148), .A2(n1275), .A3(G902), .ZN(n1273) );
NOR2_X1 U958 ( .A1(n1276), .A2(G234), .ZN(n1275) );
INV_X1 U959 ( .A(G217), .ZN(n1276) );
XNOR2_X1 U960 ( .A(n1277), .B(n1278), .ZN(n1148) );
XOR2_X1 U961 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U962 ( .A(G146), .B(G137), .Z(n1280) );
NOR2_X1 U963 ( .A1(KEYINPUT52), .A2(n1281), .ZN(n1279) );
XOR2_X1 U964 ( .A(n1282), .B(n1283), .Z(n1277) );
AND3_X1 U965 ( .A1(G221), .A2(n1093), .A3(G234), .ZN(n1283) );
NAND3_X1 U966 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1282) );
NAND2_X1 U967 ( .A1(G110), .A2(n1287), .ZN(n1286) );
OR3_X1 U968 ( .A1(n1287), .A2(G110), .A3(KEYINPUT54), .ZN(n1285) );
OR2_X1 U969 ( .A1(KEYINPUT14), .A2(n1288), .ZN(n1287) );
NAND2_X1 U970 ( .A1(KEYINPUT54), .A2(n1288), .ZN(n1284) );
XOR2_X1 U971 ( .A(n1263), .B(G128), .Z(n1288) );
NAND2_X1 U972 ( .A1(G217), .A2(G902), .ZN(n1272) );
INV_X1 U973 ( .A(n1083), .ZN(n1251) );
XOR2_X1 U974 ( .A(n1111), .B(G472), .Z(n1083) );
NAND3_X1 U975 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1111) );
OR3_X1 U976 ( .A1(n1172), .A2(n1292), .A3(KEYINPUT34), .ZN(n1290) );
INV_X1 U977 ( .A(n1293), .ZN(n1172) );
NAND2_X1 U978 ( .A1(n1294), .A2(KEYINPUT34), .ZN(n1289) );
XOR2_X1 U979 ( .A(n1295), .B(n1292), .Z(n1294) );
XNOR2_X1 U980 ( .A(n1296), .B(n1178), .ZN(n1292) );
XOR2_X1 U981 ( .A(n1297), .B(G119), .Z(n1178) );
NAND3_X1 U982 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1296) );
NAND2_X1 U983 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U984 ( .A1(KEYINPUT8), .A2(n1303), .ZN(n1302) );
XOR2_X1 U985 ( .A(KEYINPUT15), .B(n1179), .Z(n1303) );
NAND3_X1 U986 ( .A1(KEYINPUT8), .A2(n1177), .A3(n1179), .ZN(n1299) );
INV_X1 U987 ( .A(n1301), .ZN(n1177) );
XNOR2_X1 U988 ( .A(n1304), .B(KEYINPUT5), .ZN(n1301) );
OR2_X1 U989 ( .A1(n1179), .A2(KEYINPUT8), .ZN(n1298) );
NOR2_X1 U990 ( .A1(n1293), .A2(n1305), .ZN(n1295) );
XNOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT23), .ZN(n1305) );
XOR2_X1 U992 ( .A(n1306), .B(G101), .Z(n1293) );
NAND2_X1 U993 ( .A1(n1307), .A2(G210), .ZN(n1306) );
INV_X1 U994 ( .A(n1216), .ZN(n1165) );
NAND3_X1 U995 ( .A1(n1219), .A2(n1206), .A3(n1088), .ZN(n1216) );
NOR2_X1 U996 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
INV_X1 U997 ( .A(n1114), .ZN(n1090) );
NAND2_X1 U998 ( .A1(G221), .A2(n1308), .ZN(n1114) );
NAND2_X1 U999 ( .A1(G234), .A2(n1291), .ZN(n1308) );
XOR2_X1 U1000 ( .A(n1116), .B(G469), .Z(n1089) );
NAND2_X1 U1001 ( .A1(n1309), .A2(n1291), .ZN(n1116) );
XOR2_X1 U1002 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1003 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1004 ( .A(KEYINPUT2), .B(G140), .Z(n1313) );
XOR2_X1 U1005 ( .A(KEYINPUT5), .B(KEYINPUT3), .Z(n1312) );
XOR2_X1 U1006 ( .A(n1314), .B(n1315), .Z(n1310) );
INV_X1 U1007 ( .A(n1186), .ZN(n1315) );
XOR2_X1 U1008 ( .A(n1316), .B(n1317), .Z(n1186) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1123), .ZN(n1317) );
INV_X1 U1010 ( .A(G227), .ZN(n1123) );
XOR2_X1 U1011 ( .A(n1131), .B(G110), .Z(n1314) );
XOR2_X1 U1012 ( .A(n1191), .B(n1304), .Z(n1131) );
XOR2_X1 U1013 ( .A(G131), .B(n1318), .Z(n1304) );
XOR2_X1 U1014 ( .A(G137), .B(G134), .Z(n1318) );
NAND2_X1 U1015 ( .A1(n1319), .A2(n1320), .ZN(n1191) );
NAND2_X1 U1016 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n1323), .Z(n1319) );
NOR2_X1 U1018 ( .A1(n1321), .A2(n1322), .ZN(n1323) );
INV_X1 U1019 ( .A(G128), .ZN(n1322) );
XOR2_X1 U1020 ( .A(G143), .B(n1324), .Z(n1321) );
XOR2_X1 U1021 ( .A(KEYINPUT19), .B(G146), .Z(n1324) );
INV_X1 U1022 ( .A(n1068), .ZN(n1206) );
NAND2_X1 U1023 ( .A1(n1325), .A2(n1097), .ZN(n1068) );
XOR2_X1 U1024 ( .A(n1119), .B(n1326), .Z(n1097) );
NOR2_X1 U1025 ( .A1(KEYINPUT43), .A2(n1117), .ZN(n1326) );
NAND2_X1 U1026 ( .A1(n1327), .A2(n1291), .ZN(n1117) );
XNOR2_X1 U1027 ( .A(n1328), .B(n1234), .ZN(n1327) );
XNOR2_X1 U1028 ( .A(n1329), .B(n1142), .ZN(n1234) );
XOR2_X1 U1029 ( .A(G110), .B(n1330), .Z(n1142) );
NOR2_X1 U1030 ( .A1(KEYINPUT21), .A2(n1260), .ZN(n1330) );
INV_X1 U1031 ( .A(G122), .ZN(n1260) );
NAND2_X1 U1032 ( .A1(n1331), .A2(n1332), .ZN(n1329) );
NAND2_X1 U1033 ( .A1(n1141), .A2(n1333), .ZN(n1332) );
INV_X1 U1034 ( .A(KEYINPUT39), .ZN(n1333) );
XOR2_X1 U1035 ( .A(n1334), .B(n1335), .Z(n1141) );
NAND3_X1 U1036 ( .A1(n1334), .A2(n1335), .A3(KEYINPUT39), .ZN(n1331) );
INV_X1 U1037 ( .A(n1316), .ZN(n1335) );
XNOR2_X1 U1038 ( .A(G101), .B(n1336), .ZN(n1316) );
XOR2_X1 U1039 ( .A(G107), .B(G104), .Z(n1336) );
NAND2_X1 U1040 ( .A1(n1337), .A2(n1338), .ZN(n1334) );
NAND2_X1 U1041 ( .A1(n1297), .A2(G119), .ZN(n1338) );
NAND2_X1 U1042 ( .A1(n1339), .A2(n1263), .ZN(n1337) );
INV_X1 U1043 ( .A(G119), .ZN(n1263) );
XNOR2_X1 U1044 ( .A(n1297), .B(KEYINPUT37), .ZN(n1339) );
XNOR2_X1 U1045 ( .A(n1269), .B(n1340), .ZN(n1297) );
NAND2_X1 U1046 ( .A1(n1341), .A2(KEYINPUT53), .ZN(n1328) );
XOR2_X1 U1047 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1048 ( .A(KEYINPUT46), .B(n1196), .ZN(n1343) );
NAND2_X1 U1049 ( .A1(G224), .A2(n1093), .ZN(n1196) );
NAND2_X1 U1050 ( .A1(KEYINPUT28), .A2(n1233), .ZN(n1342) );
XNOR2_X1 U1051 ( .A(n1344), .B(n1179), .ZN(n1233) );
XNOR2_X1 U1052 ( .A(n1345), .B(n1346), .ZN(n1179) );
INV_X1 U1053 ( .A(G146), .ZN(n1345) );
XOR2_X1 U1054 ( .A(n1133), .B(KEYINPUT41), .Z(n1344) );
AND2_X1 U1055 ( .A1(G210), .A2(n1347), .ZN(n1119) );
XOR2_X1 U1056 ( .A(KEYINPUT18), .B(n1099), .Z(n1325) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1347), .ZN(n1099) );
NAND2_X1 U1058 ( .A1(n1348), .A2(n1291), .ZN(n1347) );
INV_X1 U1059 ( .A(G237), .ZN(n1348) );
NOR3_X1 U1060 ( .A1(n1349), .A2(n1060), .A3(n1102), .ZN(n1219) );
NOR2_X1 U1061 ( .A1(G953), .A2(G952), .ZN(n1102) );
INV_X1 U1062 ( .A(n1101), .ZN(n1060) );
NAND2_X1 U1063 ( .A1(G237), .A2(G234), .ZN(n1101) );
AND2_X1 U1064 ( .A1(G953), .A2(n1350), .ZN(n1349) );
OR2_X1 U1065 ( .A1(n1291), .A2(G898), .ZN(n1350) );
NOR2_X1 U1066 ( .A1(n1242), .A2(n1240), .ZN(n1091) );
XOR2_X1 U1067 ( .A(n1351), .B(G478), .Z(n1240) );
NAND2_X1 U1068 ( .A1(KEYINPUT32), .A2(n1110), .ZN(n1351) );
NAND2_X1 U1069 ( .A1(n1291), .A2(n1352), .ZN(n1110) );
NAND2_X1 U1070 ( .A1(n1353), .A2(n1157), .ZN(n1352) );
NAND2_X1 U1071 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
OR2_X1 U1072 ( .A1(n1159), .A2(n1158), .ZN(n1353) );
NAND3_X1 U1073 ( .A1(G234), .A2(n1093), .A3(G217), .ZN(n1158) );
INV_X1 U1074 ( .A(G953), .ZN(n1093) );
NAND2_X1 U1075 ( .A1(n1354), .A2(n1355), .ZN(n1159) );
NAND2_X1 U1076 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1077 ( .A(KEYINPUT7), .B(n1358), .Z(n1354) );
NOR2_X1 U1078 ( .A1(n1356), .A2(n1357), .ZN(n1358) );
XNOR2_X1 U1079 ( .A(n1359), .B(n1360), .ZN(n1357) );
XOR2_X1 U1080 ( .A(KEYINPUT49), .B(G122), .Z(n1360) );
XOR2_X1 U1081 ( .A(n1269), .B(G107), .Z(n1359) );
INV_X1 U1082 ( .A(G116), .ZN(n1269) );
XNOR2_X1 U1083 ( .A(G134), .B(n1346), .ZN(n1356) );
XOR2_X1 U1084 ( .A(G128), .B(G143), .Z(n1346) );
XOR2_X1 U1085 ( .A(n1361), .B(n1108), .Z(n1242) );
XNOR2_X1 U1086 ( .A(n1362), .B(G475), .ZN(n1108) );
NAND2_X1 U1087 ( .A1(n1162), .A2(n1291), .ZN(n1362) );
INV_X1 U1088 ( .A(G902), .ZN(n1291) );
XNOR2_X1 U1089 ( .A(n1363), .B(n1364), .ZN(n1162) );
XOR2_X1 U1090 ( .A(n1365), .B(n1366), .Z(n1364) );
XOR2_X1 U1091 ( .A(n1367), .B(G122), .Z(n1366) );
NAND2_X1 U1092 ( .A1(n1307), .A2(G214), .ZN(n1367) );
NOR2_X1 U1093 ( .A1(G953), .A2(G237), .ZN(n1307) );
XOR2_X1 U1094 ( .A(n1238), .B(G146), .Z(n1365) );
INV_X1 U1095 ( .A(G143), .ZN(n1238) );
XOR2_X1 U1096 ( .A(n1368), .B(n1369), .Z(n1363) );
XNOR2_X1 U1097 ( .A(n1370), .B(n1371), .ZN(n1369) );
NOR2_X1 U1098 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1371) );
NAND2_X1 U1099 ( .A1(KEYINPUT33), .A2(n1163), .ZN(n1370) );
INV_X1 U1100 ( .A(G104), .ZN(n1163) );
XNOR2_X1 U1101 ( .A(n1281), .B(n1340), .ZN(n1368) );
XOR2_X1 U1102 ( .A(G113), .B(KEYINPUT35), .Z(n1340) );
XNOR2_X1 U1103 ( .A(n1133), .B(n1372), .ZN(n1281) );
XOR2_X1 U1104 ( .A(KEYINPUT63), .B(G140), .Z(n1372) );
INV_X1 U1105 ( .A(G125), .ZN(n1133) );
XNOR2_X1 U1106 ( .A(KEYINPUT45), .B(KEYINPUT16), .ZN(n1361) );
endmodule


