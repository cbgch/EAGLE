//Key = 01101110001100011011000101111111111111100100110001100000011011000000111100011000001111
module c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, 
        G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, 
        G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, 
        G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, 
        G1698, G2897, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, 
        KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, 
        KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, 
        KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, 
        KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, 
        KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, 
        KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, 
        KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, 
        KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, 
        KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, 
        KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, 
        KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, 
        KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, 
        KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, 
        KEYINPUT83, KEYINPUT84, KEYINPUT85, G353, G355, G361, G358, G351, 
        G372_enc, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378,
                 G375, G381, G407_enc, G409, G405, G402 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3,
         KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9,
         KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
         KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
         KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
         KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
         KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
         KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39,
         KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
         KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
         KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
         KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
         KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
         KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
         KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
         KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79,
         KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84,
         KEYINPUT85;

  output G353, G355, G361, G358, G351, G372_enc, G369, G399, G364, G396, G384,
           G367, G387, G393, G390, G378, G375, G381, G407_enc, G409, G405, G402;
   wire   n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193;


  NOR3_X2 U1621 ( .A1(n2859), .A2(n2867), .A3(n2856), .ZN(n2480) );
  NOR3_X2 U1622 ( .A1(G1698), .A2(G33), .A3(n3146), .ZN(n2977) );
  NOR3_X2 U1623 ( .A1(n2855), .A2(G200), .A3(n2856), .ZN(n2479) );
  OR4_X1 U1624 ( .A1(n2382), .A2(n2383), .A3(KEYINPUT43), .A4(n2384), .ZN(G409) );
  NOR2_X1 U1625 ( .A1(G343), .A2(n2385), .ZN(n2382) );
  NOR3_X1 U1626 ( .A1(n2386), .A2(KEYINPUT42), .A3(n2384), .ZN(G407_enc) );
  NOR4_X1 U1627 ( .A1(G384), .A2(G396), .A3(n2385), .A4(n2387), .ZN(n2384) );
  OR4_X1 U1628 ( .A1(G393), .A2(G390), .A3(G387), .A4(G381), .ZN(n2387) );
  INV_X1 U1629 ( .A(KEYINPUT41), .ZN(n2386) );
  XOR2_X1 U1630 ( .A(n2388), .B(n2389), .Z(G405) );
  NAND2_X1 U1631 ( .A1(n2390), .A2(n2391), .ZN(n2388) );
  NAND2_X1 U1632 ( .A1(G2897), .A2(n2392), .ZN(n2391) );
  XOR2_X1 U1633 ( .A(n2393), .B(n2394), .Z(n2390) );
  NOR2_X1 U1634 ( .A1(n2395), .A2(n2392), .ZN(n2394) );
  OR2_X1 U1635 ( .A1(n2396), .A2(n2392), .ZN(n2393) );
  NOR2_X1 U1636 ( .A1(n2383), .A2(G343), .ZN(n2392) );
  INV_X1 U1637 ( .A(G213), .ZN(n2383) );
  NAND3_X1 U1638 ( .A1(n2397), .A2(n2398), .A3(n2399), .ZN(G402) );
  NAND2_X1 U1639 ( .A1(n2389), .A2(n2400), .ZN(n2399) );
  INV_X1 U1640 ( .A(n2385), .ZN(n2400) );
  NAND2_X1 U1641 ( .A1(n2396), .A2(n2395), .ZN(n2385) );
  INV_X1 U1642 ( .A(G378), .ZN(n2395) );
  OR3_X1 U1643 ( .A1(n2389), .A2(n2396), .A3(G378), .ZN(n2398) );
  INV_X1 U1644 ( .A(G375), .ZN(n2396) );
  NAND2_X1 U1645 ( .A1(n2401), .A2(G378), .ZN(n2397) );
  XNOR2_X1 U1646 ( .A(n2389), .B(G375), .ZN(n2401) );
  XOR2_X1 U1647 ( .A(n2402), .B(n2403), .Z(n2389) );
  XNOR2_X1 U1648 ( .A(G387), .B(n2404), .ZN(n2403) );
  XOR2_X1 U1649 ( .A(G393), .B(G390), .Z(n2404) );
  XNOR2_X1 U1650 ( .A(n2405), .B(G384), .ZN(n2402) );
  XNOR2_X1 U1651 ( .A(G381), .B(G396), .ZN(n2405) );
  NAND2_X1 U1652 ( .A1(n2406), .A2(n2407), .ZN(G396) );
  NAND2_X1 U1653 ( .A1(n2408), .A2(n2409), .ZN(n2407) );
  XNOR2_X1 U1654 ( .A(n2410), .B(n2411), .ZN(n2408) );
  NAND4_X1 U1655 ( .A1(n2412), .A2(n2413), .A3(n2414), .A4(n2415), .ZN(n2406) );
  NOR2_X1 U1656 ( .A1(n2416), .A2(n2417), .ZN(n2414) );
  NOR2_X1 U1657 ( .A1(n2418), .A2(n2419), .ZN(n2417) );
  NOR3_X1 U1658 ( .A1(n2420), .A2(n2421), .A3(n2422), .ZN(n2418) );
  NOR2_X1 U1659 ( .A1(n2423), .A2(n2424), .ZN(n2422) );
  NOR2_X1 U1660 ( .A1(n2425), .A2(n2426), .ZN(n2424) );
  AND2_X1 U1661 ( .A1(G45), .A2(n2427), .ZN(n2426) );
  NOR2_X1 U1662 ( .A1(G45), .A2(n2428), .ZN(n2425) );
  NOR3_X1 U1663 ( .A1(n2429), .A2(G116), .A3(n2430), .ZN(n2421) );
  AND2_X1 U1664 ( .A1(G355), .A2(n2430), .ZN(n2420) );
  NOR4_X1 U1665 ( .A1(n2431), .A2(n2432), .A3(n2433), .A4(n2434), .ZN(n2416) );
  NOR2_X1 U1666 ( .A1(n2435), .A2(n2436), .ZN(n2434) );
  NOR2_X1 U1667 ( .A1(n2437), .A2(n2438), .ZN(n2433) );
  NAND3_X1 U1668 ( .A1(n2439), .A2(n2440), .A3(n2441), .ZN(n2432) );
  NAND2_X1 U1669 ( .A1(n2442), .A2(G97), .ZN(n2441) );
  NAND2_X1 U1670 ( .A1(n2443), .A2(G68), .ZN(n2440) );
  NAND2_X1 U1671 ( .A1(n2444), .A2(G87), .ZN(n2439) );
  NAND4_X1 U1672 ( .A1(n2445), .A2(n2446), .A3(n2447), .A4(n2448), .ZN(n2431) );
  NAND2_X1 U1673 ( .A1(n2449), .A2(G50), .ZN(n2448) );
  NAND2_X1 U1674 ( .A1(n2450), .A2(G159), .ZN(n2447) );
  NAND2_X1 U1675 ( .A1(n2451), .A2(G58), .ZN(n2446) );
  NAND4_X1 U1676 ( .A1(KEYINPUT25), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2413) );
  OR2_X1 U1677 ( .A1(n2455), .A2(n2456), .ZN(n2454) );
  NAND3_X1 U1678 ( .A1(KEYINPUT45), .A2(n2455), .A3(n2456), .ZN(n2453) );
  NOR2_X1 U1679 ( .A1(KEYINPUT47), .A2(n2457), .ZN(n2455) );
  NAND4_X1 U1680 ( .A1(n2458), .A2(n2459), .A3(n2460), .A4(n2461), .ZN(n2412) );
  NOR4_X1 U1681 ( .A1(n2462), .A2(n2463), .A3(n2464), .A4(n2465), .ZN(n2461) );
  NOR2_X1 U1682 ( .A1(n2466), .A2(n2467), .ZN(n2464) );
  AND2_X1 U1683 ( .A1(G329), .A2(n2450), .ZN(n2463) );
  NOR2_X1 U1684 ( .A1(n2468), .A2(n2469), .ZN(n2462) );
  NOR3_X1 U1685 ( .A1(n2470), .A2(n2471), .A3(n2472), .ZN(n2460) );
  NOR2_X1 U1686 ( .A1(n2473), .A2(n2474), .ZN(n2472) );
  NOR2_X1 U1687 ( .A1(n2475), .A2(n2476), .ZN(n2471) );
  NOR2_X1 U1688 ( .A1(n2477), .A2(n2478), .ZN(n2470) );
  NAND2_X1 U1689 ( .A1(G311), .A2(n2479), .ZN(n2459) );
  NAND2_X1 U1690 ( .A1(n2480), .A2(G283), .ZN(n2458) );
  NAND3_X1 U1691 ( .A1(n2481), .A2(n2482), .A3(n2483), .ZN(G393) );
  NAND4_X1 U1692 ( .A1(n2484), .A2(n2485), .A3(n2486), .A4(n2487), .ZN(n2483) );
  NOR2_X1 U1693 ( .A1(n2488), .A2(n2409), .ZN(n2487) );
  NOR2_X1 U1694 ( .A1(n2489), .A2(n2419), .ZN(n2488) );
  NOR3_X1 U1695 ( .A1(n2490), .A2(n2491), .A3(n2492), .ZN(n2489) );
  NOR4_X1 U1696 ( .A1(n2423), .A2(KEYINPUT24), .A3(n2493), .A4(n2494), .ZN(n2492) );
  NOR2_X1 U1697 ( .A1(n2495), .A2(n2496), .ZN(n2494) );
  NOR2_X1 U1698 ( .A1(G45), .A2(n2497), .ZN(n2493) );
  NOR2_X1 U1699 ( .A1(n2498), .A2(KEYINPUT80), .ZN(n2497) );
  NOR4_X1 U1700 ( .A1(G50), .A2(n2499), .A3(n2500), .A4(n2501), .ZN(n2498) );
  NOR3_X1 U1701 ( .A1(n2429), .A2(G107), .A3(n2430), .ZN(n2491) );
  AND2_X1 U1702 ( .A1(n2501), .A2(n2430), .ZN(n2490) );
  NAND4_X1 U1703 ( .A1(n2502), .A2(n2503), .A3(n2504), .A4(n2505), .ZN(n2486) );
  NOR4_X1 U1704 ( .A1(n2506), .A2(n2507), .A3(n2508), .A4(n2509), .ZN(n2505) );
  NOR2_X1 U1705 ( .A1(n2510), .A2(n2466), .ZN(n2508) );
  NOR2_X1 U1706 ( .A1(n2511), .A2(n2512), .ZN(n2507) );
  NOR2_X1 U1707 ( .A1(n2513), .A2(n2468), .ZN(n2506) );
  NOR3_X1 U1708 ( .A1(n2514), .A2(n2515), .A3(n2516), .ZN(n2504) );
  NOR2_X1 U1709 ( .A1(n2500), .A2(n2475), .ZN(n2515) );
  NAND2_X1 U1710 ( .A1(n2479), .A2(G68), .ZN(n2503) );
  NAND4_X1 U1711 ( .A1(KEYINPUT29), .A2(n2452), .A3(n2517), .A4(n2518), .ZN(n2485) );
  OR2_X1 U1712 ( .A1(n2519), .A2(n2520), .ZN(n2518) );
  NAND3_X1 U1713 ( .A1(KEYINPUT57), .A2(n2519), .A3(n2520), .ZN(n2517) );
  NOR2_X1 U1714 ( .A1(KEYINPUT56), .A2(n2521), .ZN(n2519) );
  NAND4_X1 U1715 ( .A1(n2522), .A2(n2523), .A3(n2524), .A4(n2525), .ZN(n2484) );
  NOR4_X1 U1716 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2465), .ZN(n2525) );
  NOR2_X1 U1717 ( .A1(n2466), .A2(n2476), .ZN(n2528) );
  NOR2_X1 U1718 ( .A1(n2512), .A2(n2469), .ZN(n2527) );
  INV_X1 U1719 ( .A(G326), .ZN(n2469) );
  NOR2_X1 U1720 ( .A1(n2468), .A2(n2467), .ZN(n2526) );
  NOR3_X1 U1721 ( .A1(n2529), .A2(n2530), .A3(n2531), .ZN(n2524) );
  NOR2_X1 U1722 ( .A1(n2477), .A2(n2474), .ZN(n2531) );
  NOR2_X1 U1723 ( .A1(n2475), .A2(n2532), .ZN(n2530) );
  NOR2_X1 U1724 ( .A1(n2533), .A2(n2478), .ZN(n2529) );
  NAND2_X1 U1725 ( .A1(n2479), .A2(G303), .ZN(n2523) );
  NAND2_X1 U1726 ( .A1(n2480), .A2(G116), .ZN(n2522) );
  NAND2_X1 U1727 ( .A1(n2534), .A2(n2535), .ZN(n2482) );
  NAND3_X1 U1728 ( .A1(n2536), .A2(n2537), .A3(n2538), .ZN(n2481) );
  NAND3_X1 U1729 ( .A1(n2539), .A2(n2540), .A3(n2541), .ZN(G390) );
  NAND2_X1 U1730 ( .A1(n2542), .A2(n2535), .ZN(n2541) );
  NAND4_X1 U1731 ( .A1(n2543), .A2(n2544), .A3(n2545), .A4(n2546), .ZN(n2540) );
  NOR2_X1 U1732 ( .A1(n2547), .A2(n2409), .ZN(n2546) );
  NOR2_X1 U1733 ( .A1(n2548), .A2(n2419), .ZN(n2547) );
  NOR3_X1 U1734 ( .A1(n2430), .A2(n2549), .A3(n2550), .ZN(n2548) );
  NOR2_X1 U1735 ( .A1(n2423), .A2(n2551), .ZN(n2550) );
  NOR2_X1 U1736 ( .A1(G97), .A2(n2429), .ZN(n2549) );
  NAND4_X1 U1737 ( .A1(n2552), .A2(n2553), .A3(n2554), .A4(n2555), .ZN(n2545) );
  NOR4_X1 U1738 ( .A1(n2556), .A2(n2557), .A3(n2558), .A4(n2509), .ZN(n2555) );
  NOR2_X1 U1739 ( .A1(n2513), .A2(n2466), .ZN(n2558) );
  NOR2_X1 U1740 ( .A1(n2559), .A2(n2512), .ZN(n2557) );
  NOR2_X1 U1741 ( .A1(n2511), .A2(n2468), .ZN(n2556) );
  NOR3_X1 U1742 ( .A1(n2560), .A2(n2561), .A3(n2562), .ZN(n2554) );
  NOR2_X1 U1743 ( .A1(n2563), .A2(n2474), .ZN(n2562) );
  NOR2_X1 U1744 ( .A1(n2510), .A2(n2475), .ZN(n2561) );
  NAND2_X1 U1745 ( .A1(n2479), .A2(G58), .ZN(n2553) );
  NAND4_X1 U1746 ( .A1(KEYINPUT27), .A2(n2452), .A3(n2564), .A4(n2565), .ZN(n2544) );
  OR2_X1 U1747 ( .A1(n2566), .A2(n2567), .ZN(n2565) );
  NAND3_X1 U1748 ( .A1(KEYINPUT49), .A2(n2566), .A3(n2567), .ZN(n2564) );
  NOR2_X1 U1749 ( .A1(KEYINPUT53), .A2(n2568), .ZN(n2566) );
  INV_X1 U1750 ( .A(n2569), .ZN(n2568) );
  NAND4_X1 U1751 ( .A1(n2570), .A2(n2571), .A3(n2572), .A4(n2573), .ZN(n2543) );
  NOR4_X1 U1752 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2465), .ZN(n2573) );
  NOR2_X1 U1753 ( .A1(n2466), .A2(n2532), .ZN(n2576) );
  NOR2_X1 U1754 ( .A1(n2512), .A2(n2467), .ZN(n2575) );
  INV_X1 U1755 ( .A(G322), .ZN(n2467) );
  NOR2_X1 U1756 ( .A1(n2468), .A2(n2476), .ZN(n2574) );
  INV_X1 U1757 ( .A(G317), .ZN(n2476) );
  NOR3_X1 U1758 ( .A1(n2577), .A2(n2578), .A3(n2579), .ZN(n2572) );
  NOR2_X1 U1759 ( .A1(n2533), .A2(n2474), .ZN(n2579) );
  NOR2_X1 U1760 ( .A1(n2473), .A2(n2475), .ZN(n2578) );
  NOR2_X1 U1761 ( .A1(n2580), .A2(n2478), .ZN(n2577) );
  NAND2_X1 U1762 ( .A1(n2479), .A2(G294), .ZN(n2571) );
  NAND2_X1 U1763 ( .A1(n2480), .A2(G107), .ZN(n2570) );
  NAND3_X1 U1764 ( .A1(n2581), .A2(n2582), .A3(n2537), .ZN(n2539) );
  NAND2_X1 U1765 ( .A1(n2538), .A2(n2583), .ZN(n2582) );
  NAND2_X1 U1766 ( .A1(n2534), .A2(n2584), .ZN(n2581) );
  NAND2_X1 U1767 ( .A1(n2583), .A2(n2536), .ZN(n2584) );
  INV_X1 U1768 ( .A(n2542), .ZN(n2583) );
  OR3_X1 U1769 ( .A1(KEYINPUT81), .A2(n2585), .A3(n2586), .ZN(G387) );
  NOR2_X1 U1770 ( .A1(n2587), .A2(n2588), .ZN(n2586) );
  XOR2_X1 U1771 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR2_X1 U1772 ( .A(n2591), .B(n2592), .Z(n2590) );
  NOR2_X1 U1773 ( .A1(n2593), .A2(n2594), .ZN(n2592) );
  NOR2_X1 U1774 ( .A1(n2595), .A2(n2596), .ZN(n2591) );
  NOR2_X1 U1775 ( .A1(n2597), .A2(n2598), .ZN(n2596) );
  NAND3_X1 U1776 ( .A1(n2599), .A2(n2600), .A3(KEYINPUT32), .ZN(n2589) );
  OR2_X1 U1777 ( .A1(n2601), .A2(n2602), .ZN(n2600) );
  NAND3_X1 U1778 ( .A1(KEYINPUT61), .A2(n2601), .A3(n2602), .ZN(n2599) );
  NOR2_X1 U1779 ( .A1(KEYINPUT63), .A2(n2603), .ZN(n2601) );
  NOR2_X1 U1780 ( .A1(n2604), .A2(n2535), .ZN(n2587) );
  NAND2_X1 U1781 ( .A1(n2605), .A2(n2606), .ZN(n2535) );
  NAND2_X1 U1782 ( .A1(n2537), .A2(n2607), .ZN(n2606) );
  AND3_X1 U1783 ( .A1(n2534), .A2(n2542), .A3(n2537), .ZN(n2604) );
  NAND3_X1 U1784 ( .A1(n2608), .A2(n2609), .A3(n2610), .ZN(n2542) );
  OR2_X1 U1785 ( .A1(n2593), .A2(G399), .ZN(n2610) );
  NAND2_X1 U1786 ( .A1(n2611), .A2(n2594), .ZN(G399) );
  OR3_X1 U1787 ( .A1(n2611), .A2(n2612), .A3(n2613), .ZN(n2609) );
  NAND2_X1 U1788 ( .A1(n2613), .A2(n2614), .ZN(n2608) );
  NAND2_X1 U1789 ( .A1(n2615), .A2(n2616), .ZN(n2614) );
  NAND2_X1 U1790 ( .A1(n2593), .A2(n2611), .ZN(n2616) );
  INV_X1 U1791 ( .A(n2595), .ZN(n2615) );
  NOR2_X1 U1792 ( .A1(n2611), .A2(n2593), .ZN(n2595) );
  INV_X1 U1793 ( .A(n2612), .ZN(n2593) );
  NAND3_X1 U1794 ( .A1(n2617), .A2(n2618), .A3(KEYINPUT28), .ZN(n2612) );
  NAND2_X1 U1795 ( .A1(n2619), .A2(n2620), .ZN(n2618) );
  NAND2_X1 U1796 ( .A1(n2569), .A2(n2621), .ZN(n2619) );
  NAND4_X1 U1797 ( .A1(n2569), .A2(n2621), .A3(KEYINPUT50), .A4(n2567), .ZN(n2617) );
  INV_X1 U1798 ( .A(KEYINPUT52), .ZN(n2621) );
  NOR2_X1 U1799 ( .A1(n2622), .A2(KEYINPUT51), .ZN(n2569) );
  NOR2_X1 U1800 ( .A1(n2623), .A2(n2624), .ZN(n2622) );
  NAND2_X1 U1801 ( .A1(n2624), .A2(n2625), .ZN(n2611) );
  NAND2_X1 U1802 ( .A1(n2626), .A2(n2627), .ZN(n2625) );
  NAND2_X1 U1803 ( .A1(n2628), .A2(n2629), .ZN(n2626) );
  INV_X1 U1804 ( .A(n2594), .ZN(n2613) );
  NAND2_X1 U1805 ( .A1(n2630), .A2(n2629), .ZN(n2594) );
  INV_X1 U1806 ( .A(n2538), .ZN(n2534) );
  XOR2_X1 U1807 ( .A(n2630), .B(n2631), .Z(n2538) );
  XOR2_X1 U1808 ( .A(n2629), .B(n2632), .Z(n2631) );
  NAND2_X1 U1809 ( .A1(n2628), .A2(n2624), .ZN(n2632) );
  NAND3_X1 U1810 ( .A1(n2633), .A2(n2634), .A3(KEYINPUT30), .ZN(n2629) );
  OR2_X1 U1811 ( .A1(n2635), .A2(n2520), .ZN(n2634) );
  NAND3_X1 U1812 ( .A1(KEYINPUT58), .A2(n2635), .A3(n2520), .ZN(n2633) );
  NOR2_X1 U1813 ( .A1(KEYINPUT55), .A2(n2521), .ZN(n2635) );
  OR2_X1 U1814 ( .A1(n2636), .A2(KEYINPUT54), .ZN(n2521) );
  NOR2_X1 U1815 ( .A1(n2637), .A2(n2624), .ZN(n2636) );
  AND2_X1 U1816 ( .A1(G330), .A2(n2410), .ZN(n2630) );
  NAND3_X1 U1817 ( .A1(n2638), .A2(n2639), .A3(KEYINPUT26), .ZN(n2410) );
  OR2_X1 U1818 ( .A1(n2640), .A2(n2456), .ZN(n2639) );
  NAND3_X1 U1819 ( .A1(KEYINPUT44), .A2(n2640), .A3(n2456), .ZN(n2638) );
  NOR2_X1 U1820 ( .A1(KEYINPUT46), .A2(n2457), .ZN(n2640) );
  OR2_X1 U1821 ( .A1(n2641), .A2(KEYINPUT48), .ZN(n2457) );
  NOR2_X1 U1822 ( .A1(n2642), .A2(n2624), .ZN(n2641) );
  NOR4_X1 U1823 ( .A1(n2643), .A2(n2644), .A3(n2645), .A4(n2646), .ZN(n2585) );
  NOR4_X1 U1824 ( .A1(n2647), .A2(n2648), .A3(n2649), .A4(n2650), .ZN(n2646) );
  NOR2_X1 U1825 ( .A1(n2580), .A2(n2474), .ZN(n2650) );
  NOR2_X1 U1826 ( .A1(n2473), .A2(n2466), .ZN(n2649) );
  NAND3_X1 U1827 ( .A1(n2651), .A2(n2652), .A3(n2653), .ZN(n2648) );
  NAND2_X1 U1828 ( .A1(G317), .A2(n2450), .ZN(n2653) );
  NAND2_X1 U1829 ( .A1(G311), .A2(n2449), .ZN(n2652) );
  NAND2_X1 U1830 ( .A1(n2442), .A2(G107), .ZN(n2651) );
  NAND4_X1 U1831 ( .A1(n2654), .A2(n2655), .A3(n2502), .A4(n2656), .ZN(n2647) );
  NAND2_X1 U1832 ( .A1(n2479), .A2(G283), .ZN(n2656) );
  NAND2_X1 U1833 ( .A1(n2480), .A2(G97), .ZN(n2502) );
  NAND2_X1 U1834 ( .A1(n2443), .A2(G294), .ZN(n2655) );
  NOR2_X1 U1835 ( .A1(n2657), .A2(n2419), .ZN(n2645) );
  OR2_X1 U1836 ( .A1(n2658), .A2(n2452), .ZN(n2419) );
  NOR3_X1 U1837 ( .A1(n2430), .A2(n2659), .A3(n2660), .ZN(n2657) );
  NOR2_X1 U1838 ( .A1(n2423), .A2(n2661), .ZN(n2660) );
  INV_X1 U1839 ( .A(n2429), .ZN(n2423) );
  NOR2_X1 U1840 ( .A1(G87), .A2(n2429), .ZN(n2659) );
  NOR2_X1 U1841 ( .A1(n2662), .A2(n2663), .ZN(n2429) );
  NOR2_X1 U1842 ( .A1(n2663), .A2(G33), .ZN(n2430) );
  NOR4_X1 U1843 ( .A1(n2664), .A2(n2665), .A3(n2666), .A4(n2667), .ZN(n2644) );
  NOR2_X1 U1844 ( .A1(n2513), .A2(n2475), .ZN(n2667) );
  NOR2_X1 U1845 ( .A1(n2511), .A2(n2466), .ZN(n2666) );
  NAND3_X1 U1846 ( .A1(n2668), .A2(n2669), .A3(n2670), .ZN(n2665) );
  NAND2_X1 U1847 ( .A1(n2450), .A2(G137), .ZN(n2670) );
  NAND4_X1 U1848 ( .A1(n2445), .A2(n2671), .A3(n2672), .A4(n2673), .ZN(n2664) );
  NAND2_X1 U1849 ( .A1(n2444), .A2(G58), .ZN(n2673) );
  NAND2_X1 U1850 ( .A1(n2479), .A2(G50), .ZN(n2672) );
  NAND2_X1 U1851 ( .A1(n2449), .A2(G143), .ZN(n2671) );
  NAND2_X1 U1852 ( .A1(n2415), .A2(n2674), .ZN(n2643) );
  NAND4_X1 U1853 ( .A1(KEYINPUT31), .A2(n2452), .A3(n2675), .A4(n2676), .ZN(n2674) );
  OR2_X1 U1854 ( .A1(n2677), .A2(n2602), .ZN(n2676) );
  NAND3_X1 U1855 ( .A1(KEYINPUT60), .A2(n2677), .A3(n2602), .ZN(n2675) );
  NOR2_X1 U1856 ( .A1(KEYINPUT64), .A2(n2603), .ZN(n2677) );
  OR2_X1 U1857 ( .A1(n2678), .A2(KEYINPUT62), .ZN(n2603) );
  NOR2_X1 U1858 ( .A1(n2679), .A2(n2624), .ZN(n2678) );
  NOR2_X1 U1859 ( .A1(n2680), .A2(G20), .ZN(n2452) );
  NAND2_X1 U1860 ( .A1(n2681), .A2(n2682), .ZN(G384) );
  NAND4_X1 U1861 ( .A1(n2683), .A2(n2684), .A3(n2685), .A4(n2409), .ZN(n2682) );
  NAND2_X1 U1862 ( .A1(n2686), .A2(n2536), .ZN(n2685) );
  NAND3_X1 U1863 ( .A1(n2687), .A2(n2688), .A3(n2689), .ZN(n2684) );
  NAND2_X1 U1864 ( .A1(n2690), .A2(n2691), .ZN(n2683) );
  XNOR2_X1 U1865 ( .A(n2687), .B(n2686), .ZN(n2690) );
  NAND4_X1 U1866 ( .A1(n2692), .A2(n2693), .A3(n2694), .A4(n2415), .ZN(n2681) );
  NOR2_X1 U1867 ( .A1(n2695), .A2(n2696), .ZN(n2694) );
  NOR2_X1 U1868 ( .A1(G77), .A2(n2697), .ZN(n2696) );
  NOR4_X1 U1869 ( .A1(n2698), .A2(n2699), .A3(n2700), .A4(n2701), .ZN(n2695) );
  NOR2_X1 U1870 ( .A1(n2563), .A2(n2436), .ZN(n2701) );
  NOR2_X1 U1871 ( .A1(n2513), .A2(n2438), .ZN(n2700) );
  NAND3_X1 U1872 ( .A1(n2702), .A2(n2703), .A3(n2704), .ZN(n2699) );
  NAND2_X1 U1873 ( .A1(n2442), .A2(G58), .ZN(n2704) );
  NAND2_X1 U1874 ( .A1(n2443), .A2(G150), .ZN(n2703) );
  NAND2_X1 U1875 ( .A1(n2444), .A2(G50), .ZN(n2702) );
  INV_X1 U1876 ( .A(n2474), .ZN(n2444) );
  NAND4_X1 U1877 ( .A1(n2445), .A2(n2705), .A3(n2706), .A4(n2707), .ZN(n2698) );
  NAND2_X1 U1878 ( .A1(n2449), .A2(G137), .ZN(n2707) );
  NAND2_X1 U1879 ( .A1(G132), .A2(n2450), .ZN(n2706) );
  NAND2_X1 U1880 ( .A1(n2451), .A2(G143), .ZN(n2705) );
  NAND4_X1 U1881 ( .A1(KEYINPUT33), .A2(n2708), .A3(n2709), .A4(n2710), .ZN(n2693) );
  OR2_X1 U1882 ( .A1(n2711), .A2(n2712), .ZN(n2710) );
  NAND3_X1 U1883 ( .A1(KEYINPUT71), .A2(n2711), .A3(n2712), .ZN(n2709) );
  NOR2_X1 U1884 ( .A1(KEYINPUT74), .A2(n2713), .ZN(n2711) );
  NAND4_X1 U1885 ( .A1(n2552), .A2(n2714), .A3(n2715), .A4(n2716), .ZN(n2692) );
  NOR4_X1 U1886 ( .A1(n2717), .A2(n2718), .A3(n2719), .A4(n2465), .ZN(n2716) );
  NOR2_X1 U1887 ( .A1(n2477), .A2(n2466), .ZN(n2719) );
  NOR2_X1 U1888 ( .A1(n2512), .A2(n2532), .ZN(n2718) );
  INV_X1 U1889 ( .A(G311), .ZN(n2532) );
  NOR2_X1 U1890 ( .A1(n2473), .A2(n2468), .ZN(n2717) );
  NOR3_X1 U1891 ( .A1(n2720), .A2(n2721), .A3(n2722), .ZN(n2715) );
  NOR2_X1 U1892 ( .A1(n2435), .A2(n2474), .ZN(n2722) );
  NOR2_X1 U1893 ( .A1(n2533), .A2(n2475), .ZN(n2721) );
  NOR2_X1 U1894 ( .A1(n2723), .A2(n2478), .ZN(n2720) );
  NAND2_X1 U1895 ( .A1(n2479), .A2(G116), .ZN(n2714) );
  NAND2_X1 U1896 ( .A1(n2480), .A2(G87), .ZN(n2552) );
  NAND3_X1 U1897 ( .A1(n2724), .A2(n2725), .A3(n2726), .ZN(G381) );
  NAND2_X1 U1898 ( .A1(n2727), .A2(n2728), .ZN(n2726) );
  NAND4_X1 U1899 ( .A1(n2729), .A2(n2730), .A3(n2731), .A4(n2732), .ZN(n2725) );
  NOR2_X1 U1900 ( .A1(n2733), .A2(n2409), .ZN(n2732) );
  NOR2_X1 U1901 ( .A1(G68), .A2(n2697), .ZN(n2733) );
  NAND4_X1 U1902 ( .A1(n2734), .A2(n2735), .A3(n2736), .A4(n2737), .ZN(n2731) );
  NOR4_X1 U1903 ( .A1(n2738), .A2(n2739), .A3(n2740), .A4(n2509), .ZN(n2737) );
  NOR2_X1 U1904 ( .A1(n2741), .A2(n2466), .ZN(n2740) );
  NOR2_X1 U1905 ( .A1(n2742), .A2(n2512), .ZN(n2739) );
  NOR2_X1 U1906 ( .A1(n2468), .A2(n2743), .ZN(n2738) );
  NOR3_X1 U1907 ( .A1(n2744), .A2(n2745), .A3(n2746), .ZN(n2736) );
  NOR2_X1 U1908 ( .A1(n2513), .A2(n2474), .ZN(n2746) );
  NOR2_X1 U1909 ( .A1(n2475), .A2(n2559), .ZN(n2745) );
  NOR2_X1 U1910 ( .A1(n2510), .A2(n2478), .ZN(n2744) );
  NAND2_X1 U1911 ( .A1(n2479), .A2(G150), .ZN(n2735) );
  NAND2_X1 U1912 ( .A1(n2480), .A2(G58), .ZN(n2734) );
  NAND4_X1 U1913 ( .A1(KEYINPUT35), .A2(n2708), .A3(n2747), .A4(n2748), .ZN(n2730) );
  OR2_X1 U1914 ( .A1(n2749), .A2(n2750), .ZN(n2748) );
  NAND3_X1 U1915 ( .A1(KEYINPUT76), .A2(n2749), .A3(n2750), .ZN(n2747) );
  NOR2_X1 U1916 ( .A1(KEYINPUT79), .A2(n2751), .ZN(n2749) );
  NAND4_X1 U1917 ( .A1(n2668), .A2(n2752), .A3(n2753), .A4(n2754), .ZN(n2729) );
  NOR4_X1 U1918 ( .A1(n2755), .A2(n2756), .A3(n2757), .A4(n2465), .ZN(n2754) );
  NOR2_X1 U1919 ( .A1(n2533), .A2(n2466), .ZN(n2757) );
  NOR2_X1 U1920 ( .A1(n2473), .A2(n2512), .ZN(n2756) );
  INV_X1 U1921 ( .A(G303), .ZN(n2473) );
  NOR2_X1 U1922 ( .A1(n2477), .A2(n2468), .ZN(n2755) );
  NOR3_X1 U1923 ( .A1(n2514), .A2(n2758), .A3(n2759), .ZN(n2753) );
  NOR2_X1 U1924 ( .A1(n2723), .A2(n2474), .ZN(n2759) );
  NOR2_X1 U1925 ( .A1(n2580), .A2(n2475), .ZN(n2758) );
  NOR2_X1 U1926 ( .A1(n2760), .A2(n2478), .ZN(n2514) );
  NAND2_X1 U1927 ( .A1(n2479), .A2(G107), .ZN(n2752) );
  NAND2_X1 U1928 ( .A1(n2480), .A2(G77), .ZN(n2668) );
  NAND2_X1 U1929 ( .A1(n2761), .A2(n2537), .ZN(n2724) );
  XNOR2_X1 U1930 ( .A(n2762), .B(n2763), .ZN(n2761) );
  NAND3_X1 U1931 ( .A1(n2764), .A2(n2765), .A3(KEYINPUT38), .ZN(n2762) );
  OR2_X1 U1932 ( .A1(n2766), .A2(n2767), .ZN(n2765) );
  NAND3_X1 U1933 ( .A1(KEYINPUT69), .A2(n2766), .A3(n2767), .ZN(n2764) );
  NOR2_X1 U1934 ( .A1(KEYINPUT67), .A2(n2768), .ZN(n2767) );
  NAND3_X1 U1935 ( .A1(n2769), .A2(n2770), .A3(n2771), .ZN(G378) );
  NAND4_X1 U1936 ( .A1(n2772), .A2(n2773), .A3(n2774), .A4(n2775), .ZN(n2771) );
  NOR2_X1 U1937 ( .A1(n2776), .A2(n2409), .ZN(n2775) );
  NOR2_X1 U1938 ( .A1(G58), .A2(n2697), .ZN(n2776) );
  NAND2_X1 U1939 ( .A1(n2777), .A2(n2680), .ZN(n2697) );
  NAND3_X1 U1940 ( .A1(n2778), .A2(n2708), .A3(KEYINPUT82), .ZN(n2774) );
  NAND4_X1 U1941 ( .A1(n2779), .A2(n2780), .A3(n2781), .A4(n2782), .ZN(n2773) );
  NOR4_X1 U1942 ( .A1(n2783), .A2(n2784), .A3(n2785), .A4(n2509), .ZN(n2782) );
  NOR2_X1 U1943 ( .A1(n2466), .A2(n2743), .ZN(n2785) );
  AND2_X1 U1944 ( .A1(n2450), .A2(G125), .ZN(n2784) );
  NOR2_X1 U1945 ( .A1(n2468), .A2(n2742), .ZN(n2783) );
  NOR3_X1 U1946 ( .A1(n2786), .A2(n2787), .A3(n2788), .ZN(n2781) );
  NOR2_X1 U1947 ( .A1(n2511), .A2(n2474), .ZN(n2788) );
  INV_X1 U1948 ( .A(G150), .ZN(n2511) );
  NOR2_X1 U1949 ( .A1(n2475), .A2(n2741), .ZN(n2787) );
  INV_X1 U1950 ( .A(G137), .ZN(n2741) );
  NOR2_X1 U1951 ( .A1(n2513), .A2(n2478), .ZN(n2786) );
  NAND2_X1 U1952 ( .A1(G143), .A2(n2479), .ZN(n2780) );
  NAND2_X1 U1953 ( .A1(n2480), .A2(G50), .ZN(n2779) );
  NAND4_X1 U1954 ( .A1(n2789), .A2(n2790), .A3(n2791), .A4(n2792), .ZN(n2772) );
  NOR4_X1 U1955 ( .A1(n2793), .A2(n2794), .A3(n2795), .A4(n2465), .ZN(n2792) );
  INV_X1 U1956 ( .A(n2654), .ZN(n2465) );
  NOR2_X1 U1957 ( .A1(n2580), .A2(n2466), .ZN(n2795) );
  NOR2_X1 U1958 ( .A1(n2477), .A2(n2512), .ZN(n2794) );
  INV_X1 U1959 ( .A(G294), .ZN(n2477) );
  NOR2_X1 U1960 ( .A1(n2533), .A2(n2468), .ZN(n2793) );
  NOR3_X1 U1961 ( .A1(n2560), .A2(n2796), .A3(n2797), .ZN(n2791) );
  NOR2_X1 U1962 ( .A1(n2760), .A2(n2474), .ZN(n2797) );
  NOR2_X1 U1963 ( .A1(n2435), .A2(n2475), .ZN(n2796) );
  NOR2_X1 U1964 ( .A1(n2437), .A2(n2478), .ZN(n2560) );
  NAND2_X1 U1965 ( .A1(n2479), .A2(G97), .ZN(n2790) );
  NAND2_X1 U1966 ( .A1(n2480), .A2(G68), .ZN(n2789) );
  NAND3_X1 U1967 ( .A1(n2798), .A2(n2409), .A3(n2799), .ZN(n2770) );
  NAND3_X1 U1968 ( .A1(n2800), .A2(n2727), .A3(n2605), .ZN(n2798) );
  NAND4_X1 U1969 ( .A1(n2800), .A2(n2727), .A3(n2537), .A4(n2801), .ZN(n2769) );
  INV_X1 U1970 ( .A(n2799), .ZN(n2801) );
  NAND4_X1 U1971 ( .A1(n2802), .A2(n2803), .A3(n2804), .A4(n2805), .ZN(G375) );
  NAND3_X1 U1972 ( .A1(n2806), .A2(n2807), .A3(n2409), .ZN(n2805) );
  INV_X1 U1973 ( .A(n2415), .ZN(n2409) );
  NAND3_X1 U1974 ( .A1(n2808), .A2(n2809), .A3(KEYINPUT1), .ZN(n2807) );
  NAND2_X1 U1975 ( .A1(n2810), .A2(n2811), .ZN(n2809) );
  NAND2_X1 U1976 ( .A1(n2812), .A2(n2813), .ZN(n2811) );
  INV_X1 U1977 ( .A(n2814), .ZN(n2810) );
  NAND4_X1 U1978 ( .A1(n2812), .A2(n2813), .A3(KEYINPUT5), .A4(n2814), .ZN(n2808) );
  INV_X1 U1979 ( .A(KEYINPUT8), .ZN(n2813) );
  NAND2_X1 U1980 ( .A1(n2605), .A2(n2815), .ZN(n2806) );
  NAND3_X1 U1981 ( .A1(n2727), .A2(n2799), .A3(n2800), .ZN(n2815) );
  NAND3_X1 U1982 ( .A1(n2816), .A2(n2817), .A3(KEYINPUT15), .ZN(n2799) );
  NAND2_X1 U1983 ( .A1(n2818), .A2(n2819), .ZN(n2817) );
  NAND3_X1 U1984 ( .A1(n2820), .A2(n2821), .A3(n2822), .ZN(n2819) );
  XNOR2_X1 U1985 ( .A(n2823), .B(n2824), .ZN(n2818) );
  NAND3_X1 U1986 ( .A1(KEYINPUT23), .A2(n2825), .A3(n2826), .ZN(n2816) );
  AND3_X1 U1987 ( .A1(n2822), .A2(n2821), .A3(n2820), .ZN(n2826) );
  NAND2_X1 U1988 ( .A1(KEYINPUT59), .A2(G330), .ZN(n2820) );
  INV_X1 U1989 ( .A(KEYINPUT22), .ZN(n2821) );
  NAND3_X1 U1990 ( .A1(n2827), .A2(n2688), .A3(n2687), .ZN(n2822) );
  XNOR2_X1 U1991 ( .A(n2823), .B(n2828), .ZN(n2825) );
  NAND3_X1 U1992 ( .A1(n2829), .A2(n2830), .A3(KEYINPUT37), .ZN(n2727) );
  OR2_X1 U1993 ( .A1(n2766), .A2(n2831), .ZN(n2830) );
  NAND3_X1 U1994 ( .A1(KEYINPUT68), .A2(n2766), .A3(n2831), .ZN(n2829) );
  NOR2_X1 U1995 ( .A1(KEYINPUT66), .A2(n2768), .ZN(n2831) );
  OR2_X1 U1996 ( .A1(n2832), .A2(KEYINPUT65), .ZN(n2768) );
  AND2_X1 U1997 ( .A1(n2688), .A2(n2687), .ZN(n2832) );
  XOR2_X1 U1998 ( .A(n2833), .B(n2827), .Z(n2766) );
  INV_X1 U1999 ( .A(n2728), .ZN(n2605) );
  NAND4_X1 U2000 ( .A1(n2834), .A2(n2835), .A3(n2836), .A4(n2415), .ZN(n2804) );
  NOR2_X1 U2001 ( .A1(n2728), .A2(n2537), .ZN(n2415) );
  NAND2_X1 U2002 ( .A1(G1), .A2(n2837), .ZN(n2728) );
  NAND3_X1 U2003 ( .A1(G13), .A2(n2838), .A3(G45), .ZN(n2837) );
  NOR2_X1 U2004 ( .A1(n2839), .A2(n2840), .ZN(n2836) );
  NOR4_X1 U2005 ( .A1(n2841), .A2(n2842), .A3(n2843), .A4(n2509), .ZN(n2840) );
  INV_X1 U2006 ( .A(n2445), .ZN(n2509) );
  NOR2_X1 U2007 ( .A1(n2777), .A2(G33), .ZN(n2445) );
  NOR2_X1 U2008 ( .A1(n2742), .A2(n2466), .ZN(n2843) );
  INV_X1 U2009 ( .A(n2451), .ZN(n2466) );
  INV_X1 U2010 ( .A(G128), .ZN(n2742) );
  NAND3_X1 U2011 ( .A1(n2844), .A2(n2845), .A3(n2846), .ZN(n2842) );
  NAND2_X1 U2012 ( .A1(G124), .A2(n2450), .ZN(n2846) );
  NAND2_X1 U2013 ( .A1(n2480), .A2(G159), .ZN(n2845) );
  NAND2_X1 U2014 ( .A1(G125), .A2(n2449), .ZN(n2844) );
  NAND3_X1 U2015 ( .A1(n2847), .A2(n2848), .A3(n2849), .ZN(n2841) );
  NOR3_X1 U2016 ( .A1(n2850), .A2(G41), .A3(n2851), .ZN(n2849) );
  NOR2_X1 U2017 ( .A1(n2475), .A2(n2743), .ZN(n2851) );
  INV_X1 U2018 ( .A(G132), .ZN(n2743) );
  INV_X1 U2019 ( .A(n2443), .ZN(n2475) );
  NOR2_X1 U2020 ( .A1(n2474), .A2(n2559), .ZN(n2850) );
  INV_X1 U2021 ( .A(G143), .ZN(n2559) );
  NAND2_X1 U2022 ( .A1(n2442), .A2(G150), .ZN(n2848) );
  NAND2_X1 U2023 ( .A1(n2479), .A2(G137), .ZN(n2847) );
  NOR4_X1 U2024 ( .A1(n2852), .A2(n2853), .A3(n2516), .A4(n2854), .ZN(n2839) );
  NOR2_X1 U2025 ( .A1(n2760), .A2(n2438), .ZN(n2854) );
  INV_X1 U2026 ( .A(n2479), .ZN(n2438) );
  NOR2_X1 U2027 ( .A1(n2437), .A2(n2474), .ZN(n2516) );
  NAND4_X1 U2028 ( .A1(G200), .A2(G190), .A3(G20), .A4(n2855), .ZN(n2474) );
  NAND3_X1 U2029 ( .A1(n2669), .A2(n2857), .A3(n2858), .ZN(n2853) );
  NAND2_X1 U2030 ( .A1(n2443), .A2(G97), .ZN(n2858) );
  NOR3_X1 U2031 ( .A1(n2855), .A2(n2859), .A3(n2856), .ZN(n2443) );
  NAND2_X1 U2032 ( .A1(n2442), .A2(G68), .ZN(n2669) );
  INV_X1 U2033 ( .A(n2478), .ZN(n2442) );
  NAND3_X1 U2034 ( .A1(n2855), .A2(n2856), .A3(n2860), .ZN(n2478) );
  NAND2_X1 U2035 ( .A1(G200), .A2(G20), .ZN(n2860) );
  NAND3_X1 U2036 ( .A1(n2654), .A2(n2861), .A3(n2862), .ZN(n2852) );
  NOR3_X1 U2037 ( .A1(n2863), .A2(n2864), .A3(n2865), .ZN(n2862) );
  NOR2_X1 U2038 ( .A1(n2580), .A2(n2468), .ZN(n2865) );
  INV_X1 U2039 ( .A(n2449), .ZN(n2468) );
  NOR3_X1 U2040 ( .A1(n2859), .A2(n2866), .A3(n2855), .ZN(n2449) );
  NOR2_X1 U2041 ( .A1(n2500), .A2(n2436), .ZN(n2864) );
  INV_X1 U2042 ( .A(n2480), .ZN(n2436) );
  INV_X1 U2043 ( .A(G200), .ZN(n2859) );
  NOR2_X1 U2044 ( .A1(n2533), .A2(n2512), .ZN(n2863) );
  INV_X1 U2045 ( .A(n2450), .ZN(n2512) );
  NOR3_X1 U2046 ( .A1(n2867), .A2(G200), .A3(n2856), .ZN(n2450) );
  INV_X1 U2047 ( .A(n2866), .ZN(n2856) );
  INV_X1 U2048 ( .A(G283), .ZN(n2533) );
  NAND2_X1 U2049 ( .A1(n2451), .A2(G107), .ZN(n2861) );
  NOR3_X1 U2050 ( .A1(n2866), .A2(G200), .A3(n2855), .ZN(n2451) );
  INV_X1 U2051 ( .A(n2867), .ZN(n2855) );
  NOR2_X1 U2052 ( .A1(n2868), .A2(n2838), .ZN(n2867) );
  NOR2_X1 U2053 ( .A1(n2838), .A2(G190), .ZN(n2866) );
  NOR2_X1 U2054 ( .A1(n2777), .A2(n2662), .ZN(n2654) );
  NAND3_X1 U2055 ( .A1(n2869), .A2(n2510), .A3(n2680), .ZN(n2835) );
  INV_X1 U2056 ( .A(n2708), .ZN(n2680) );
  NAND2_X1 U2057 ( .A1(n2658), .A2(n2857), .ZN(n2869) );
  INV_X1 U2058 ( .A(n2777), .ZN(n2658) );
  NAND2_X1 U2059 ( .A1(n2870), .A2(n2871), .ZN(n2777) );
  NAND2_X1 U2060 ( .A1(G20), .A2(n2872), .ZN(n2871) );
  NAND3_X1 U2061 ( .A1(KEYINPUT84), .A2(n2873), .A3(n2708), .ZN(n2834) );
  NOR2_X1 U2062 ( .A1(G13), .A2(G33), .ZN(n2708) );
  INV_X1 U2063 ( .A(KEYINPUT39), .ZN(n2803) );
  NAND3_X1 U2064 ( .A1(n2874), .A2(n2763), .A3(n2537), .ZN(n2802) );
  INV_X1 U2065 ( .A(n2800), .ZN(n2763) );
  NOR3_X1 U2066 ( .A1(KEYINPUT0), .A2(n2875), .A3(n2876), .ZN(n2800) );
  NOR2_X1 U2067 ( .A1(n2877), .A2(n2411), .ZN(n2875) );
  NOR2_X1 U2068 ( .A1(KEYINPUT12), .A2(n2878), .ZN(n2877) );
  NAND3_X1 U2069 ( .A1(n2879), .A2(n2880), .A3(KEYINPUT2), .ZN(n2874) );
  OR2_X1 U2070 ( .A1(n2814), .A2(n2881), .ZN(n2880) );
  NAND3_X1 U2071 ( .A1(KEYINPUT6), .A2(n2814), .A3(n2881), .ZN(n2879) );
  NOR2_X1 U2072 ( .A1(KEYINPUT9), .A2(n2882), .ZN(n2881) );
  INV_X1 U2073 ( .A(n2812), .ZN(n2882) );
  NOR2_X1 U2074 ( .A1(KEYINPUT7), .A2(n2883), .ZN(n2812) );
  NOR2_X1 U2075 ( .A1(n2884), .A2(n2411), .ZN(n2883) );
  NOR2_X1 U2076 ( .A1(KEYINPUT20), .A2(n2885), .ZN(n2884) );
  XOR2_X1 U2077 ( .A(n2886), .B(n2887), .Z(n2814) );
  NAND2_X1 U2078 ( .A1(KEYINPUT85), .A2(n2873), .ZN(n2886) );
  XNOR2_X1 U2079 ( .A(n2888), .B(n2889), .ZN(n2873) );
  NOR2_X1 U2080 ( .A1(n2890), .A2(n2891), .ZN(n2889) );
  OR2_X1 U2081 ( .A1(n2892), .A2(KEYINPUT14), .ZN(G372_enc) );
  NOR2_X1 U2082 ( .A1(n2893), .A2(n2894), .ZN(n2892) );
  NAND2_X1 U2083 ( .A1(n2895), .A2(n2896), .ZN(G369) );
  NAND2_X1 U2084 ( .A1(n2897), .A2(n2898), .ZN(n2896) );
  NAND3_X1 U2085 ( .A1(n2899), .A2(n2900), .A3(n2901), .ZN(G367) );
  NAND2_X1 U2086 ( .A1(n2902), .A2(n2903), .ZN(n2901) );
  NAND3_X1 U2087 ( .A1(n2904), .A2(n2905), .A3(n2906), .ZN(n2903) );
  NAND2_X1 U2088 ( .A1(G68), .A2(n2510), .ZN(n2906) );
  NAND4_X1 U2089 ( .A1(G50), .A2(n2563), .A3(G77), .A4(G58), .ZN(n2905) );
  NAND2_X1 U2090 ( .A1(n2499), .A2(n2500), .ZN(n2904) );
  NOR2_X1 U2091 ( .A1(n2563), .A2(n2437), .ZN(n2499) );
  NAND3_X1 U2092 ( .A1(n2907), .A2(n2908), .A3(n2909), .ZN(n2900) );
  NAND2_X1 U2093 ( .A1(KEYINPUT4), .A2(n2910), .ZN(n2907) );
  NAND2_X1 U2094 ( .A1(n2911), .A2(n2912), .ZN(n2910) );
  NAND2_X1 U2095 ( .A1(n2913), .A2(n2914), .ZN(n2912) );
  NAND3_X1 U2096 ( .A1(n2915), .A2(n2916), .A3(KEYINPUT16), .ZN(n2914) );
  XOR2_X1 U2097 ( .A(n2876), .B(n2887), .Z(n2913) );
  NAND3_X1 U2098 ( .A1(n2915), .A2(n2916), .A3(n2917), .ZN(n2911) );
  XNOR2_X1 U2099 ( .A(n2887), .B(n2876), .ZN(n2917) );
  NAND2_X1 U2100 ( .A1(n2895), .A2(n2918), .ZN(n2876) );
  NAND2_X1 U2101 ( .A1(n2691), .A2(n2897), .ZN(n2918) );
  INV_X1 U2102 ( .A(n2893), .ZN(n2897) );
  AND3_X1 U2103 ( .A1(n2919), .A2(n2920), .A3(n2921), .ZN(n2895) );
  NAND2_X1 U2104 ( .A1(n2888), .A2(n2922), .ZN(n2921) );
  NAND2_X1 U2105 ( .A1(n2923), .A2(n2924), .ZN(n2922) );
  NAND2_X1 U2106 ( .A1(n2925), .A2(n2926), .ZN(n2924) );
  NAND2_X1 U2107 ( .A1(n2927), .A2(n2928), .ZN(n2926) );
  NAND2_X1 U2108 ( .A1(n2750), .A2(n2929), .ZN(n2928) );
  NAND2_X1 U2109 ( .A1(n2930), .A2(n2931), .ZN(n2887) );
  NAND2_X1 U2110 ( .A1(n2824), .A2(n2823), .ZN(n2931) );
  NAND2_X1 U2111 ( .A1(n2932), .A2(n2933), .ZN(n2823) );
  NAND2_X1 U2112 ( .A1(n2827), .A2(n2833), .ZN(n2933) );
  NAND2_X1 U2113 ( .A1(n2934), .A2(n2935), .ZN(n2833) );
  NAND2_X1 U2114 ( .A1(n2691), .A2(n2688), .ZN(n2935) );
  NAND2_X1 U2115 ( .A1(n2929), .A2(n2624), .ZN(n2934) );
  INV_X1 U2116 ( .A(n2936), .ZN(n2929) );
  OR2_X1 U2117 ( .A1(n2927), .A2(n2597), .ZN(n2932) );
  OR2_X1 U2118 ( .A1(n2923), .A2(n2937), .ZN(n2930) );
  INV_X1 U2119 ( .A(KEYINPUT17), .ZN(n2916) );
  NAND2_X1 U2120 ( .A1(G330), .A2(n2938), .ZN(n2915) );
  NAND4_X1 U2121 ( .A1(n2939), .A2(n2940), .A3(KEYINPUT18), .A4(n2941), .ZN(n2938) );
  NOR2_X1 U2122 ( .A1(KEYINPUT40), .A2(n2942), .ZN(n2941) );
  INV_X1 U2123 ( .A(KEYINPUT10), .ZN(n2942) );
  NAND3_X1 U2124 ( .A1(KEYINPUT19), .A2(n2943), .A3(n2944), .ZN(n2940) );
  INV_X1 U2125 ( .A(n2945), .ZN(n2944) );
  NAND3_X1 U2126 ( .A1(KEYINPUT11), .A2(n2946), .A3(n2945), .ZN(n2939) );
  NOR3_X1 U2127 ( .A1(KEYINPUT13), .A2(KEYINPUT12), .A3(n2878), .ZN(n2945) );
  NOR2_X1 U2128 ( .A1(n2947), .A2(n2893), .ZN(n2878) );
  NAND4_X1 U2129 ( .A1(n2712), .A2(n2888), .A3(n2925), .A4(n2750), .ZN(n2893) );
  AND3_X1 U2130 ( .A1(n2919), .A2(n2920), .A3(n2948), .ZN(n2888) );
  NAND3_X1 U2131 ( .A1(n2949), .A2(n2950), .A3(n2890), .ZN(n2948) );
  INV_X1 U2132 ( .A(n2951), .ZN(n2890) );
  NAND2_X1 U2133 ( .A1(G200), .A2(n2952), .ZN(n2950) );
  NAND2_X1 U2134 ( .A1(G190), .A2(n2953), .ZN(n2949) );
  NAND3_X1 U2135 ( .A1(n2953), .A2(n2951), .A3(G179), .ZN(n2920) );
  INV_X1 U2136 ( .A(n2952), .ZN(n2953) );
  NAND3_X1 U2137 ( .A1(n2952), .A2(n2951), .A3(G169), .ZN(n2919) );
  NAND4_X1 U2138 ( .A1(n2954), .A2(n2955), .A3(n2956), .A4(n2957), .ZN(n2951) );
  NOR2_X1 U2139 ( .A1(n2958), .A2(n2959), .ZN(n2957) );
  NOR2_X1 U2140 ( .A1(n2960), .A2(n2500), .ZN(n2959) );
  NOR2_X1 U2141 ( .A1(n2961), .A2(n2962), .ZN(n2958) );
  NAND2_X1 U2142 ( .A1(G150), .A2(n2963), .ZN(n2956) );
  NAND2_X1 U2143 ( .A1(n2964), .A2(n2510), .ZN(n2955) );
  INV_X1 U2144 ( .A(G50), .ZN(n2510) );
  NAND2_X1 U2145 ( .A1(n2965), .A2(G50), .ZN(n2954) );
  NAND3_X1 U2146 ( .A1(n2966), .A2(n2967), .A3(n2968), .ZN(n2952) );
  NOR3_X1 U2147 ( .A1(n2969), .A2(n2970), .A3(n2971), .ZN(n2968) );
  NOR2_X1 U2148 ( .A1(n2972), .A2(n2973), .ZN(n2971) );
  NOR2_X1 U2149 ( .A1(n2974), .A2(n2975), .ZN(n2969) );
  INV_X1 U2150 ( .A(G223), .ZN(n2975) );
  NAND2_X1 U2151 ( .A1(G77), .A2(n2976), .ZN(n2967) );
  NAND2_X1 U2152 ( .A1(G222), .A2(n2977), .ZN(n2966) );
  INV_X1 U2153 ( .A(n2943), .ZN(n2946) );
  NOR3_X1 U2154 ( .A1(KEYINPUT21), .A2(KEYINPUT20), .A3(n2885), .ZN(n2943) );
  NOR4_X1 U2155 ( .A1(n2828), .A2(n2978), .A3(n2686), .A4(n2947), .ZN(n2885) );
  INV_X1 U2156 ( .A(n2688), .ZN(n2686) );
  NAND3_X1 U2157 ( .A1(n2979), .A2(n2980), .A3(KEYINPUT34), .ZN(n2688) );
  OR2_X1 U2158 ( .A1(n2981), .A2(n2712), .ZN(n2980) );
  NAND3_X1 U2159 ( .A1(KEYINPUT70), .A2(n2981), .A3(n2712), .ZN(n2979) );
  AND2_X1 U2160 ( .A1(n2982), .A2(n2936), .ZN(n2712) );
  NAND3_X1 U2161 ( .A1(n2983), .A2(n2984), .A3(n2985), .ZN(n2936) );
  NAND2_X1 U2162 ( .A1(n2986), .A2(n2868), .ZN(n2984) );
  NAND2_X1 U2163 ( .A1(n2987), .A2(n2872), .ZN(n2983) );
  NAND3_X1 U2164 ( .A1(n2988), .A2(n2989), .A3(n2990), .ZN(n2982) );
  NAND2_X1 U2165 ( .A1(G200), .A2(n2987), .ZN(n2989) );
  NAND2_X1 U2166 ( .A1(n2986), .A2(G190), .ZN(n2988) );
  INV_X1 U2167 ( .A(n2987), .ZN(n2986) );
  NAND3_X1 U2168 ( .A1(n2991), .A2(n2992), .A3(n2993), .ZN(n2987) );
  NOR3_X1 U2169 ( .A1(n2994), .A2(n2970), .A3(n2995), .ZN(n2993) );
  NOR2_X1 U2170 ( .A1(n2972), .A2(n2996), .ZN(n2995) );
  NOR2_X1 U2171 ( .A1(n2974), .A2(n2997), .ZN(n2994) );
  NAND2_X1 U2172 ( .A1(G107), .A2(n2976), .ZN(n2992) );
  NAND2_X1 U2173 ( .A1(G232), .A2(n2977), .ZN(n2991) );
  NOR2_X1 U2174 ( .A1(KEYINPUT73), .A2(n2713), .ZN(n2981) );
  OR2_X1 U2175 ( .A1(n2998), .A2(KEYINPUT72), .ZN(n2713) );
  NOR2_X1 U2176 ( .A1(n2990), .A2(n2624), .ZN(n2998) );
  INV_X1 U2177 ( .A(n2985), .ZN(n2990) );
  NAND4_X1 U2178 ( .A1(n2999), .A2(n3000), .A3(n3001), .A4(n3002), .ZN(n2985) );
  NAND2_X1 U2179 ( .A1(n2964), .A2(n2437), .ZN(n3002) );
  NAND2_X1 U2180 ( .A1(G77), .A2(n3003), .ZN(n3001) );
  NAND2_X1 U2181 ( .A1(n2962), .A2(n3004), .ZN(n3003) );
  INV_X1 U2182 ( .A(n2965), .ZN(n3004) );
  NAND2_X1 U2183 ( .A1(G87), .A2(n3005), .ZN(n3000) );
  NAND2_X1 U2184 ( .A1(n2963), .A2(G58), .ZN(n2999) );
  INV_X1 U2185 ( .A(n2827), .ZN(n2978) );
  NAND3_X1 U2186 ( .A1(n3006), .A2(n3007), .A3(KEYINPUT36), .ZN(n2827) );
  OR2_X1 U2187 ( .A1(n3008), .A2(n2750), .ZN(n3007) );
  NAND3_X1 U2188 ( .A1(KEYINPUT75), .A2(n3008), .A3(n2750), .ZN(n3006) );
  AND2_X1 U2189 ( .A1(n3009), .A2(n2927), .ZN(n2750) );
  NAND3_X1 U2190 ( .A1(n3010), .A2(n3011), .A3(n3012), .ZN(n2927) );
  NAND2_X1 U2191 ( .A1(n3013), .A2(n2868), .ZN(n3011) );
  NAND2_X1 U2192 ( .A1(n3014), .A2(n2872), .ZN(n3010) );
  NAND3_X1 U2193 ( .A1(n3015), .A2(n3016), .A3(n3017), .ZN(n3009) );
  NAND2_X1 U2194 ( .A1(G200), .A2(n3014), .ZN(n3016) );
  NAND2_X1 U2195 ( .A1(n3013), .A2(G190), .ZN(n3015) );
  INV_X1 U2196 ( .A(n3014), .ZN(n3013) );
  NAND3_X1 U2197 ( .A1(n3018), .A2(n3019), .A3(n3020), .ZN(n3014) );
  NOR3_X1 U2198 ( .A1(n3021), .A2(n2970), .A3(n3022), .ZN(n3020) );
  NOR2_X1 U2199 ( .A1(n2972), .A2(n2997), .ZN(n3022) );
  INV_X1 U2200 ( .A(G238), .ZN(n2997) );
  NOR2_X1 U2201 ( .A1(n2974), .A2(n3023), .ZN(n3021) );
  NAND2_X1 U2202 ( .A1(G97), .A2(n2976), .ZN(n3019) );
  NAND2_X1 U2203 ( .A1(n2977), .A2(G226), .ZN(n3018) );
  NOR2_X1 U2204 ( .A1(KEYINPUT78), .A2(n2751), .ZN(n3008) );
  OR2_X1 U2205 ( .A1(n3024), .A2(KEYINPUT77), .ZN(n2751) );
  NOR2_X1 U2206 ( .A1(n3017), .A2(n2624), .ZN(n3024) );
  INV_X1 U2207 ( .A(n3012), .ZN(n3017) );
  NAND4_X1 U2208 ( .A1(n3025), .A2(n3026), .A3(n3027), .A4(n3028), .ZN(n3012) );
  NAND2_X1 U2209 ( .A1(n2965), .A2(G68), .ZN(n3028) );
  NAND2_X1 U2210 ( .A1(n3029), .A2(n2563), .ZN(n3027) );
  NAND2_X1 U2211 ( .A1(G77), .A2(n3005), .ZN(n3026) );
  NAND2_X1 U2212 ( .A1(G50), .A2(n2963), .ZN(n3025) );
  INV_X1 U2213 ( .A(n2824), .ZN(n2828) );
  NAND2_X1 U2214 ( .A1(KEYINPUT83), .A2(n2778), .ZN(n2824) );
  XNOR2_X1 U2215 ( .A(n2925), .B(n3030), .ZN(n2778) );
  NOR2_X1 U2216 ( .A1(n3031), .A2(n2891), .ZN(n3030) );
  AND2_X1 U2217 ( .A1(n3032), .A2(n2923), .ZN(n2925) );
  NAND3_X1 U2218 ( .A1(n3033), .A2(n3034), .A3(n3035), .ZN(n2923) );
  NAND2_X1 U2219 ( .A1(n3036), .A2(n2868), .ZN(n3034) );
  NAND2_X1 U2220 ( .A1(n3037), .A2(n2872), .ZN(n3033) );
  NAND3_X1 U2221 ( .A1(n3038), .A2(n3039), .A3(n3031), .ZN(n3032) );
  INV_X1 U2222 ( .A(n3035), .ZN(n3031) );
  NAND4_X1 U2223 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n3035) );
  NOR2_X1 U2224 ( .A1(n3044), .A2(n3045), .ZN(n3043) );
  NOR2_X1 U2225 ( .A1(n3046), .A2(n2513), .ZN(n3045) );
  INV_X1 U2226 ( .A(G159), .ZN(n2513) );
  NOR2_X1 U2227 ( .A1(n2960), .A2(n2563), .ZN(n3044) );
  OR2_X1 U2228 ( .A1(n3047), .A2(n2962), .ZN(n3042) );
  NAND2_X1 U2229 ( .A1(n2964), .A2(n2500), .ZN(n3041) );
  NAND2_X1 U2230 ( .A1(n2965), .A2(G58), .ZN(n3040) );
  NOR2_X1 U2231 ( .A1(n3048), .A2(n3049), .ZN(n2965) );
  NAND2_X1 U2232 ( .A1(G200), .A2(n3037), .ZN(n3039) );
  NAND2_X1 U2233 ( .A1(n3036), .A2(G190), .ZN(n3038) );
  INV_X1 U2234 ( .A(n3037), .ZN(n3036) );
  NAND3_X1 U2235 ( .A1(n3050), .A2(n3051), .A3(n3052), .ZN(n3037) );
  NOR3_X1 U2236 ( .A1(n3053), .A2(n2970), .A3(n3054), .ZN(n3052) );
  NOR2_X1 U2237 ( .A1(n2972), .A2(n3023), .ZN(n3054) );
  INV_X1 U2238 ( .A(G232), .ZN(n3023) );
  OR2_X1 U2239 ( .A1(n3055), .A2(n3056), .ZN(n2972) );
  AND2_X1 U2240 ( .A1(G274), .A2(n3055), .ZN(n2970) );
  NAND2_X1 U2241 ( .A1(n3057), .A2(n3058), .ZN(n3055) );
  NAND2_X1 U2242 ( .A1(G41), .A2(n3059), .ZN(n3058) );
  NOR2_X1 U2243 ( .A1(n2973), .A2(n2974), .ZN(n3053) );
  INV_X1 U2244 ( .A(G226), .ZN(n2973) );
  NAND2_X1 U2245 ( .A1(G87), .A2(n2976), .ZN(n3051) );
  NAND2_X1 U2246 ( .A1(n2977), .A2(G223), .ZN(n3050) );
  NAND3_X1 U2247 ( .A1(G116), .A2(n3060), .A3(n3061), .ZN(n2899) );
  NAND3_X1 U2248 ( .A1(n3062), .A2(n3063), .A3(n3064), .ZN(G364) );
  NAND2_X1 U2249 ( .A1(n2428), .A2(n2537), .ZN(n3064) );
  INV_X1 U2250 ( .A(n3065), .ZN(n2428) );
  OR3_X1 U2251 ( .A1(n2501), .A2(n2537), .A3(n3059), .ZN(n3063) );
  NOR2_X1 U2252 ( .A1(n2663), .A2(G41), .ZN(n2537) );
  NAND2_X1 U2253 ( .A1(n3066), .A2(n2580), .ZN(n2501) );
  NAND2_X1 U2254 ( .A1(n2607), .A2(n3059), .ZN(n3062) );
  INV_X1 U2255 ( .A(n2536), .ZN(n2607) );
  NOR2_X1 U2256 ( .A1(n2691), .A2(n2687), .ZN(n2536) );
  NOR2_X1 U2257 ( .A1(n2411), .A2(n2947), .ZN(n2687) );
  NOR3_X1 U2258 ( .A1(n3067), .A2(n3068), .A3(KEYINPUT3), .ZN(n2947) );
  NOR2_X1 U2259 ( .A1(n2624), .A2(n3069), .ZN(n3068) );
  NOR2_X1 U2260 ( .A1(n3070), .A2(n3071), .ZN(n3069) );
  NOR2_X1 U2261 ( .A1(n2868), .A2(n3072), .ZN(n3071) );
  NAND4_X1 U2262 ( .A1(n3073), .A2(n3074), .A3(n3075), .A4(n3076), .ZN(n3072) );
  NOR2_X1 U2263 ( .A1(G179), .A2(n3077), .ZN(n3070) );
  NAND4_X1 U2264 ( .A1(n3078), .A2(n3079), .A3(n3080), .A4(n3081), .ZN(n3077) );
  NOR2_X1 U2265 ( .A1(n2597), .A2(n2894), .ZN(n3067) );
  NAND4_X1 U2266 ( .A1(n2456), .A2(n2602), .A3(n2567), .A4(n2520), .ZN(n2894) );
  AND2_X1 U2267 ( .A1(n3082), .A2(n3083), .ZN(n2456) );
  NAND3_X1 U2268 ( .A1(n3084), .A2(n3085), .A3(n2642), .ZN(n3082) );
  INV_X1 U2269 ( .A(n3086), .ZN(n2642) );
  NAND2_X1 U2270 ( .A1(G200), .A2(n3081), .ZN(n3085) );
  NAND2_X1 U2271 ( .A1(n3073), .A2(G190), .ZN(n3084) );
  INV_X1 U2272 ( .A(n2624), .ZN(n2597) );
  INV_X1 U2273 ( .A(G330), .ZN(n2411) );
  INV_X1 U2274 ( .A(n2689), .ZN(n2691) );
  NAND2_X1 U2275 ( .A1(n2624), .A2(n2898), .ZN(n2689) );
  NAND3_X1 U2276 ( .A1(n3087), .A2(n3088), .A3(n3089), .ZN(n2898) );
  NAND2_X1 U2277 ( .A1(n2602), .A2(n3090), .ZN(n3089) );
  NAND2_X1 U2278 ( .A1(n2598), .A2(n3091), .ZN(n3090) );
  NAND2_X1 U2279 ( .A1(n2567), .A2(n3092), .ZN(n3091) );
  NAND2_X1 U2280 ( .A1(n2627), .A2(n3093), .ZN(n3092) );
  NAND2_X1 U2281 ( .A1(n2520), .A2(n2628), .ZN(n3093) );
  INV_X1 U2282 ( .A(n3083), .ZN(n2628) );
  NAND3_X1 U2283 ( .A1(n3094), .A2(n3095), .A3(n3086), .ZN(n3083) );
  NAND4_X1 U2284 ( .A1(n3096), .A2(n3097), .A3(n3098), .A4(n3099), .ZN(n3086) );
  NAND2_X1 U2285 ( .A1(n2964), .A2(n2580), .ZN(n3099) );
  INV_X1 U2286 ( .A(G116), .ZN(n2580) );
  NAND2_X1 U2287 ( .A1(G116), .A2(n3100), .ZN(n3098) );
  NAND2_X1 U2288 ( .A1(n3101), .A2(n2962), .ZN(n3100) );
  NAND2_X1 U2289 ( .A1(G283), .A2(n3005), .ZN(n3097) );
  NAND2_X1 U2290 ( .A1(G97), .A2(n2963), .ZN(n3096) );
  NAND2_X1 U2291 ( .A1(n3073), .A2(n2868), .ZN(n3095) );
  INV_X1 U2292 ( .A(n3081), .ZN(n3073) );
  NAND2_X1 U2293 ( .A1(n3081), .A2(n2872), .ZN(n3094) );
  NAND3_X1 U2294 ( .A1(n3102), .A2(n3103), .A3(n3104), .ZN(n3081) );
  NOR3_X1 U2295 ( .A1(n3105), .A2(n3106), .A3(n3107), .ZN(n3104) );
  NOR2_X1 U2296 ( .A1(n3108), .A2(n3109), .ZN(n3107) );
  INV_X1 U2297 ( .A(G270), .ZN(n3109) );
  NOR2_X1 U2298 ( .A1(n2974), .A2(n3110), .ZN(n3105) );
  NAND2_X1 U2299 ( .A1(G303), .A2(n2976), .ZN(n3103) );
  NAND2_X1 U2300 ( .A1(G257), .A2(n2977), .ZN(n3102) );
  AND2_X1 U2301 ( .A1(n3111), .A2(n2627), .ZN(n2520) );
  NAND3_X1 U2302 ( .A1(n3112), .A2(n3113), .A3(n2637), .ZN(n3111) );
  INV_X1 U2303 ( .A(n3114), .ZN(n2637) );
  NAND2_X1 U2304 ( .A1(G200), .A2(n3078), .ZN(n3113) );
  NAND2_X1 U2305 ( .A1(n3074), .A2(G190), .ZN(n3112) );
  NAND3_X1 U2306 ( .A1(n3115), .A2(n3116), .A3(n3114), .ZN(n2627) );
  NAND4_X1 U2307 ( .A1(n3117), .A2(n3118), .A3(n3119), .A4(n3120), .ZN(n3114) );
  NAND2_X1 U2308 ( .A1(n3121), .A2(G107), .ZN(n3120) );
  NAND2_X1 U2309 ( .A1(n3029), .A2(n2435), .ZN(n3119) );
  NAND2_X1 U2310 ( .A1(n3122), .A2(n2962), .ZN(n3029) );
  NAND2_X1 U2311 ( .A1(G116), .A2(n3005), .ZN(n3118) );
  NAND2_X1 U2312 ( .A1(G87), .A2(n2963), .ZN(n3117) );
  NAND2_X1 U2313 ( .A1(n3074), .A2(n2868), .ZN(n3116) );
  INV_X1 U2314 ( .A(n3078), .ZN(n3074) );
  NAND2_X1 U2315 ( .A1(n3078), .A2(n2872), .ZN(n3115) );
  NAND3_X1 U2316 ( .A1(n3123), .A2(n3124), .A3(n3125), .ZN(n3078) );
  NOR3_X1 U2317 ( .A1(n3126), .A2(n3106), .A3(n3127), .ZN(n3125) );
  NOR2_X1 U2318 ( .A1(n3108), .A2(n3110), .ZN(n3127) );
  INV_X1 U2319 ( .A(G264), .ZN(n3110) );
  NOR2_X1 U2320 ( .A1(n2974), .A2(n3128), .ZN(n3126) );
  NAND2_X1 U2321 ( .A1(G294), .A2(n2976), .ZN(n3124) );
  NAND2_X1 U2322 ( .A1(G250), .A2(n2977), .ZN(n3123) );
  INV_X1 U2323 ( .A(n2620), .ZN(n2567) );
  NAND2_X1 U2324 ( .A1(n3129), .A2(n2598), .ZN(n2620) );
  NAND3_X1 U2325 ( .A1(n3130), .A2(n3131), .A3(n2623), .ZN(n3129) );
  INV_X1 U2326 ( .A(n3132), .ZN(n2623) );
  NAND2_X1 U2327 ( .A1(G200), .A2(n3079), .ZN(n3131) );
  NAND2_X1 U2328 ( .A1(n3075), .A2(G190), .ZN(n3130) );
  NAND3_X1 U2329 ( .A1(n3133), .A2(n3134), .A3(n3132), .ZN(n2598) );
  NAND4_X1 U2330 ( .A1(n3135), .A2(n3136), .A3(n3137), .A4(n3138), .ZN(n3132) );
  NOR2_X1 U2331 ( .A1(n3139), .A2(n3140), .ZN(n3138) );
  NOR2_X1 U2332 ( .A1(n3046), .A2(n2437), .ZN(n3140) );
  INV_X1 U2333 ( .A(n2963), .ZN(n3046) );
  NOR2_X1 U2334 ( .A1(n2960), .A2(n2435), .ZN(n3139) );
  OR2_X1 U2335 ( .A1(n3060), .A2(n2962), .ZN(n3137) );
  NAND2_X1 U2336 ( .A1(n2964), .A2(n2723), .ZN(n3136) );
  NAND2_X1 U2337 ( .A1(n3121), .A2(G97), .ZN(n3135) );
  NAND2_X1 U2338 ( .A1(n3075), .A2(n2868), .ZN(n3134) );
  INV_X1 U2339 ( .A(G179), .ZN(n2868) );
  INV_X1 U2340 ( .A(n3079), .ZN(n3075) );
  NAND2_X1 U2341 ( .A1(n3079), .A2(n2872), .ZN(n3133) );
  INV_X1 U2342 ( .A(G169), .ZN(n2872) );
  NAND3_X1 U2343 ( .A1(n3141), .A2(n3142), .A3(n3143), .ZN(n3079) );
  NOR3_X1 U2344 ( .A1(n3144), .A2(n3106), .A3(n3145), .ZN(n3143) );
  NOR2_X1 U2345 ( .A1(n3108), .A2(n3128), .ZN(n3145) );
  NAND2_X1 U2346 ( .A1(n3146), .A2(n3147), .ZN(n3108) );
  NAND2_X1 U2347 ( .A1(n3148), .A2(n2857), .ZN(n3147) );
  AND3_X1 U2348 ( .A1(G274), .A2(n2857), .A3(n3148), .ZN(n3106) );
  INV_X1 U2349 ( .A(G41), .ZN(n2857) );
  NOR2_X1 U2350 ( .A1(n2974), .A2(n3149), .ZN(n3144) );
  NAND2_X1 U2351 ( .A1(G283), .A2(n2976), .ZN(n3142) );
  NAND2_X1 U2352 ( .A1(G244), .A2(n2977), .ZN(n3141) );
  AND3_X1 U2353 ( .A1(n3150), .A2(n3088), .A3(n3087), .ZN(n2602) );
  NAND3_X1 U2354 ( .A1(n3151), .A2(n3152), .A3(n2679), .ZN(n3150) );
  INV_X1 U2355 ( .A(n3153), .ZN(n2679) );
  NAND2_X1 U2356 ( .A1(G200), .A2(n3080), .ZN(n3152) );
  NAND2_X1 U2357 ( .A1(n3076), .A2(G190), .ZN(n3151) );
  NAND3_X1 U2358 ( .A1(G179), .A2(n3153), .A3(n3076), .ZN(n3088) );
  INV_X1 U2359 ( .A(n3080), .ZN(n3076) );
  NAND3_X1 U2360 ( .A1(n3153), .A2(n3080), .A3(G169), .ZN(n3087) );
  NAND4_X1 U2361 ( .A1(n3154), .A2(n3155), .A3(n3156), .A4(n3157), .ZN(n3080) );
  NOR2_X1 U2362 ( .A1(n3158), .A2(n3159), .ZN(n3157) );
  AND2_X1 U2363 ( .A1(n2976), .A2(G116), .ZN(n3159) );
  NOR2_X1 U2364 ( .A1(n3146), .A2(n2662), .ZN(n2976) );
  NOR2_X1 U2365 ( .A1(n2974), .A2(n2996), .ZN(n3158) );
  NAND3_X1 U2366 ( .A1(n3056), .A2(n2662), .A3(G1698), .ZN(n2974) );
  INV_X1 U2367 ( .A(n3146), .ZN(n3056) );
  NAND2_X1 U2368 ( .A1(G238), .A2(n2977), .ZN(n3156) );
  NAND3_X1 U2369 ( .A1(G250), .A2(n3146), .A3(n3057), .ZN(n3155) );
  INV_X1 U2370 ( .A(n3148), .ZN(n3057) );
  NAND2_X1 U2371 ( .A1(n2870), .A2(n3160), .ZN(n3146) );
  NAND2_X1 U2372 ( .A1(G41), .A2(G33), .ZN(n3160) );
  NAND2_X1 U2373 ( .A1(n3148), .A2(G274), .ZN(n3154) );
  NOR2_X1 U2374 ( .A1(n2495), .A2(G1), .ZN(n3148) );
  INV_X1 U2375 ( .A(G45), .ZN(n2495) );
  NAND4_X1 U2376 ( .A1(n3161), .A2(n3162), .A3(n3163), .A4(n3164), .ZN(n3153) );
  NOR2_X1 U2377 ( .A1(n3165), .A2(n3166), .ZN(n3164) );
  NOR2_X1 U2378 ( .A1(n2960), .A2(n2723), .ZN(n3166) );
  INV_X1 U2379 ( .A(n3005), .ZN(n2960) );
  NOR3_X1 U2380 ( .A1(n3167), .A2(G20), .A3(n2662), .ZN(n3005) );
  NOR2_X1 U2381 ( .A1(n3066), .A2(n2962), .ZN(n3165) );
  NAND2_X1 U2382 ( .A1(G20), .A2(n3048), .ZN(n2962) );
  INV_X1 U2383 ( .A(n3167), .ZN(n3048) );
  NOR3_X1 U2384 ( .A1(G87), .A2(G97), .A3(G107), .ZN(n3066) );
  NAND2_X1 U2385 ( .A1(G68), .A2(n2963), .ZN(n3163) );
  NOR3_X1 U2386 ( .A1(G20), .A2(G33), .A3(n3167), .ZN(n2963) );
  NAND2_X1 U2387 ( .A1(n2964), .A2(n2760), .ZN(n3162) );
  INV_X1 U2388 ( .A(G87), .ZN(n2760) );
  INV_X1 U2389 ( .A(n3122), .ZN(n2964) );
  NAND2_X1 U2390 ( .A1(n3121), .A2(G87), .ZN(n3161) );
  INV_X1 U2391 ( .A(n3101), .ZN(n3121) );
  NAND3_X1 U2392 ( .A1(n3168), .A2(n3122), .A3(n3167), .ZN(n3101) );
  NOR2_X1 U2393 ( .A1(n3169), .A2(n2870), .ZN(n3167) );
  NOR3_X1 U2394 ( .A1(n2838), .A2(n3059), .A3(n2662), .ZN(n3169) );
  INV_X1 U2395 ( .A(G33), .ZN(n2662) );
  NAND2_X1 U2396 ( .A1(n3049), .A2(G13), .ZN(n3122) );
  NOR2_X1 U2397 ( .A1(n2838), .A2(G1), .ZN(n3049) );
  NAND2_X1 U2398 ( .A1(G33), .A2(n3059), .ZN(n3168) );
  NAND2_X1 U2399 ( .A1(G343), .A2(n2937), .ZN(n2624) );
  INV_X1 U2400 ( .A(n2891), .ZN(n2937) );
  NAND4_X1 U2401 ( .A1(G213), .A2(G13), .A3(n3059), .A4(n2838), .ZN(n2891) );
  NOR3_X1 U2402 ( .A1(n3170), .A2(n3171), .A3(n3172), .ZN(G361) );
  NOR3_X1 U2403 ( .A1(n2663), .A2(n3173), .A3(n3149), .ZN(n3172) );
  INV_X1 U2404 ( .A(G250), .ZN(n3149) );
  NOR2_X1 U2405 ( .A1(G257), .A2(G264), .ZN(n3173) );
  INV_X1 U2406 ( .A(n3174), .ZN(n2663) );
  NOR3_X1 U2407 ( .A1(n3174), .A2(n3061), .A3(n3175), .ZN(n3171) );
  NOR2_X1 U2408 ( .A1(n3176), .A2(n3177), .ZN(n3175) );
  NAND4_X1 U2409 ( .A1(n3178), .A2(n3179), .A3(n3180), .A4(n3181), .ZN(n3177) );
  NAND2_X1 U2410 ( .A1(G238), .A2(G68), .ZN(n3181) );
  NAND2_X1 U2411 ( .A1(G244), .A2(G77), .ZN(n3180) );
  NAND2_X1 U2412 ( .A1(G250), .A2(G87), .ZN(n3179) );
  NAND2_X1 U2413 ( .A1(G257), .A2(G97), .ZN(n3178) );
  NAND4_X1 U2414 ( .A1(n3182), .A2(n3183), .A3(n3184), .A4(n3185), .ZN(n3176) );
  NAND2_X1 U2415 ( .A1(G264), .A2(G107), .ZN(n3185) );
  NAND2_X1 U2416 ( .A1(G270), .A2(G116), .ZN(n3184) );
  NAND2_X1 U2417 ( .A1(G226), .A2(G50), .ZN(n3183) );
  NAND2_X1 U2418 ( .A1(G232), .A2(G58), .ZN(n3182) );
  INV_X1 U2419 ( .A(n2909), .ZN(n3061) );
  NOR2_X1 U2420 ( .A1(n2838), .A2(n2908), .ZN(n3174) );
  INV_X1 U2421 ( .A(n2902), .ZN(n2908) );
  NOR2_X1 U2422 ( .A1(n3059), .A2(G13), .ZN(n2902) );
  INV_X1 U2423 ( .A(G1), .ZN(n3059) );
  INV_X1 U2424 ( .A(G20), .ZN(n2838) );
  NOR2_X1 U2425 ( .A1(n3065), .A2(n2909), .ZN(n3170) );
  NAND2_X1 U2426 ( .A1(n2870), .A2(G20), .ZN(n2909) );
  AND2_X1 U2427 ( .A1(G13), .A2(G1), .ZN(n2870) );
  NAND2_X1 U2428 ( .A1(G50), .A2(n3186), .ZN(n3065) );
  NAND2_X1 U2429 ( .A1(n2500), .A2(n2563), .ZN(n3186) );
  INV_X1 U2430 ( .A(G58), .ZN(n2500) );
  XOR2_X1 U2431 ( .A(n2661), .B(n2496), .Z(G358) );
  XNOR2_X1 U2432 ( .A(n3187), .B(n3188), .ZN(n2496) );
  XNOR2_X1 U2433 ( .A(n2996), .B(G238), .ZN(n3188) );
  INV_X1 U2434 ( .A(G244), .ZN(n2996) );
  XNOR2_X1 U2435 ( .A(G226), .B(G232), .ZN(n3187) );
  XOR2_X1 U2436 ( .A(n3189), .B(n3190), .Z(n2661) );
  XNOR2_X1 U2437 ( .A(n3128), .B(G250), .ZN(n3190) );
  INV_X1 U2438 ( .A(G257), .ZN(n3128) );
  XNOR2_X1 U2439 ( .A(G270), .B(G264), .ZN(n3189) );
  NAND2_X1 U2440 ( .A1(G87), .A2(n3191), .ZN(G355) );
  NAND2_X1 U2441 ( .A1(n2435), .A2(n2723), .ZN(n3191) );
  INV_X1 U2442 ( .A(G107), .ZN(n2435) );
  AND2_X1 U2443 ( .A1(n2437), .A2(n2961), .ZN(G353) );
  NOR3_X1 U2444 ( .A1(G58), .A2(G68), .A3(G50), .ZN(n2961) );
  INV_X1 U2445 ( .A(G77), .ZN(n2437) );
  XOR2_X1 U2446 ( .A(n2551), .B(n2427), .Z(G351) );
  XNOR2_X1 U2447 ( .A(n3192), .B(n3047), .ZN(n2427) );
  XNOR2_X1 U2448 ( .A(G58), .B(n2563), .ZN(n3047) );
  INV_X1 U2449 ( .A(G68), .ZN(n2563) );
  XNOR2_X1 U2450 ( .A(G50), .B(G77), .ZN(n3192) );
  XOR2_X1 U2451 ( .A(n3193), .B(n3060), .Z(n2551) );
  XNOR2_X1 U2452 ( .A(G107), .B(n2723), .ZN(n3060) );
  INV_X1 U2453 ( .A(G97), .ZN(n2723) );
  XNOR2_X1 U2454 ( .A(G116), .B(G87), .ZN(n3193) );
endmodule

