//Key = 0110101010110100100001000101111010100001101000101100000011001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378;

XNOR2_X1 U755 ( .A(G107), .B(n1047), .ZN(G9) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U757 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
NAND2_X1 U758 ( .A1(G952), .A2(n1054), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND4_X1 U760 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1050) );
NAND3_X1 U761 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1058) );
XNOR2_X1 U762 ( .A(n1055), .B(KEYINPUT6), .ZN(n1063) );
AND4_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1055) );
NAND3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1064), .ZN(n1057) );
INV_X1 U765 ( .A(n1070), .ZN(n1064) );
NAND2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND3_X1 U767 ( .A1(n1067), .A2(n1073), .A3(n1066), .ZN(n1072) );
OR2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1076), .ZN(n1071) );
NAND3_X1 U770 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1080), .A2(n1066), .ZN(n1079) );
INV_X1 U772 ( .A(n1081), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1067), .A2(n1082), .ZN(n1077) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR3_X1 U776 ( .A1(n1087), .A2(G953), .A3(n1088), .ZN(n1048) );
INV_X1 U777 ( .A(n1059), .ZN(n1088) );
NAND4_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1059) );
NOR4_X1 U779 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
XOR2_X1 U780 ( .A(G472), .B(n1097), .Z(n1096) );
XNOR2_X1 U781 ( .A(KEYINPUT44), .B(n1098), .ZN(n1095) );
XOR2_X1 U782 ( .A(KEYINPUT3), .B(n1099), .Z(n1094) );
NOR3_X1 U783 ( .A1(n1085), .A2(n1100), .A3(n1062), .ZN(n1091) );
NAND2_X1 U784 ( .A1(n1101), .A2(G478), .ZN(n1090) );
XOR2_X1 U785 ( .A(n1102), .B(KEYINPUT26), .Z(n1101) );
XOR2_X1 U786 ( .A(n1103), .B(n1104), .Z(n1089) );
NAND2_X1 U787 ( .A1(KEYINPUT16), .A2(n1105), .ZN(n1104) );
XNOR2_X1 U788 ( .A(G952), .B(KEYINPUT30), .ZN(n1087) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(G72) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U793 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U794 ( .A(n1116), .B(n1117), .Z(n1112) );
XNOR2_X1 U795 ( .A(G140), .B(n1118), .ZN(n1117) );
NOR2_X1 U796 ( .A1(KEYINPUT50), .A2(n1119), .ZN(n1118) );
NAND2_X1 U797 ( .A1(KEYINPUT28), .A2(G131), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1060), .ZN(n1108) );
XOR2_X1 U799 ( .A(n1121), .B(KEYINPUT59), .Z(n1120) );
NAND2_X1 U800 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U801 ( .A1(G953), .A2(n1124), .ZN(n1106) );
NAND2_X1 U802 ( .A1(G900), .A2(G227), .ZN(n1124) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U804 ( .A1(n1127), .A2(G953), .ZN(n1126) );
XNOR2_X1 U805 ( .A(n1128), .B(n1129), .ZN(n1127) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U807 ( .A1(n1132), .A2(n1060), .ZN(n1125) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1053), .ZN(n1134) );
NAND2_X1 U810 ( .A1(n1128), .A2(n1136), .ZN(n1133) );
XNOR2_X1 U811 ( .A(n1135), .B(KEYINPUT31), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NAND2_X1 U813 ( .A1(G953), .A2(n1131), .ZN(n1138) );
XOR2_X1 U814 ( .A(n1139), .B(n1140), .Z(n1137) );
NAND2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
XOR2_X1 U816 ( .A(n1143), .B(KEYINPUT22), .Z(n1141) );
NOR2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U818 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1150), .ZN(G63) );
XOR2_X1 U821 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U822 ( .A1(n1148), .A2(G478), .ZN(n1151) );
NOR2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(G60) );
XOR2_X1 U824 ( .A(KEYINPUT36), .B(n1144), .Z(n1154) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1153) );
NAND3_X1 U826 ( .A1(n1148), .A2(G475), .A3(KEYINPUT27), .ZN(n1155) );
XNOR2_X1 U827 ( .A(G104), .B(n1157), .ZN(G6) );
NAND3_X1 U828 ( .A1(n1074), .A2(n1158), .A3(n1159), .ZN(n1157) );
XNOR2_X1 U829 ( .A(n1067), .B(KEYINPUT46), .ZN(n1159) );
NOR2_X1 U830 ( .A1(n1144), .A2(n1160), .ZN(G57) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1161) );
XNOR2_X1 U834 ( .A(KEYINPUT32), .B(n1167), .ZN(n1166) );
NAND3_X1 U835 ( .A1(n1148), .A2(G472), .A3(KEYINPUT4), .ZN(n1165) );
NOR2_X1 U836 ( .A1(n1144), .A2(n1168), .ZN(G54) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U838 ( .A(n1164), .B(n1171), .Z(n1170) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(n1169) );
NOR2_X1 U840 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U841 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XNOR2_X1 U842 ( .A(n1178), .B(KEYINPUT33), .ZN(n1177) );
NAND2_X1 U843 ( .A1(n1148), .A2(G469), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1144), .A2(n1179), .ZN(G51) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1180) );
XOR2_X1 U848 ( .A(KEYINPUT43), .B(n1186), .Z(n1185) );
NAND2_X1 U849 ( .A1(n1148), .A2(n1187), .ZN(n1184) );
AND2_X1 U850 ( .A1(G902), .A2(n1188), .ZN(n1148) );
NAND2_X1 U851 ( .A1(n1136), .A2(n1189), .ZN(n1188) );
XNOR2_X1 U852 ( .A(KEYINPUT38), .B(n1052), .ZN(n1189) );
NAND2_X1 U853 ( .A1(n1122), .A2(n1190), .ZN(n1052) );
XNOR2_X1 U854 ( .A(KEYINPUT21), .B(n1123), .ZN(n1190) );
AND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1122) );
AND4_X1 U856 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
NOR4_X1 U857 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1191) );
INV_X1 U858 ( .A(n1201), .ZN(n1200) );
AND4_X1 U859 ( .A1(KEYINPUT9), .A2(n1202), .A3(n1203), .A4(n1056), .ZN(n1198) );
NOR2_X1 U860 ( .A1(KEYINPUT9), .A2(n1204), .ZN(n1197) );
INV_X1 U861 ( .A(n1053), .ZN(n1136) );
NAND4_X1 U862 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1053) );
AND3_X1 U863 ( .A1(n1209), .A2(n1047), .A3(n1210), .ZN(n1208) );
NAND3_X1 U864 ( .A1(n1075), .A2(n1067), .A3(n1158), .ZN(n1047) );
NAND2_X1 U865 ( .A1(n1065), .A2(n1211), .ZN(n1207) );
NAND2_X1 U866 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND3_X1 U867 ( .A1(n1066), .A2(n1214), .A3(n1215), .ZN(n1213) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1158), .ZN(n1212) );
XNOR2_X1 U869 ( .A(n1080), .B(KEYINPUT2), .ZN(n1216) );
NAND3_X1 U870 ( .A1(n1158), .A2(n1067), .A3(n1074), .ZN(n1206) );
NAND2_X1 U871 ( .A1(n1056), .A2(n1217), .ZN(n1205) );
NAND2_X1 U872 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR2_X1 U873 ( .A1(n1060), .A2(G952), .ZN(n1144) );
XNOR2_X1 U874 ( .A(G146), .B(n1196), .ZN(G48) );
NAND3_X1 U875 ( .A1(n1215), .A2(n1074), .A3(n1220), .ZN(n1196) );
XNOR2_X1 U876 ( .A(G143), .B(n1204), .ZN(G45) );
NAND3_X1 U877 ( .A1(n1221), .A2(n1056), .A3(n1202), .ZN(n1204) );
XOR2_X1 U878 ( .A(n1222), .B(n1223), .Z(G42) );
NOR2_X1 U879 ( .A1(KEYINPUT7), .A2(n1224), .ZN(n1223) );
NAND2_X1 U880 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
OR2_X1 U881 ( .A1(n1195), .A2(KEYINPUT15), .ZN(n1226) );
NAND2_X1 U882 ( .A1(n1227), .A2(n1068), .ZN(n1195) );
NAND3_X1 U883 ( .A1(n1227), .A2(n1228), .A3(KEYINPUT15), .ZN(n1225) );
AND3_X1 U884 ( .A1(n1080), .A2(n1074), .A3(n1220), .ZN(n1227) );
NAND3_X1 U885 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(G39) );
OR2_X1 U886 ( .A1(n1201), .A2(G137), .ZN(n1231) );
NAND2_X1 U887 ( .A1(KEYINPUT0), .A2(n1232), .ZN(n1230) );
NAND2_X1 U888 ( .A1(G137), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U889 ( .A(KEYINPUT8), .B(n1201), .ZN(n1233) );
NAND2_X1 U890 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
INV_X1 U891 ( .A(KEYINPUT0), .ZN(n1235) );
NAND2_X1 U892 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
NAND3_X1 U893 ( .A1(KEYINPUT8), .A2(G137), .A3(n1201), .ZN(n1237) );
OR2_X1 U894 ( .A1(n1201), .A2(KEYINPUT8), .ZN(n1236) );
NAND3_X1 U895 ( .A1(n1068), .A2(n1220), .A3(n1238), .ZN(n1201) );
XNOR2_X1 U896 ( .A(G134), .B(n1194), .ZN(G36) );
NAND3_X1 U897 ( .A1(n1202), .A2(n1075), .A3(n1068), .ZN(n1194) );
NAND3_X1 U898 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(G33) );
NAND2_X1 U899 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U900 ( .A1(n1244), .A2(n1245), .ZN(n1240) );
INV_X1 U901 ( .A(KEYINPUT13), .ZN(n1245) );
NAND2_X1 U902 ( .A1(n1246), .A2(G131), .ZN(n1244) );
XNOR2_X1 U903 ( .A(n1242), .B(KEYINPUT5), .ZN(n1246) );
NAND2_X1 U904 ( .A1(KEYINPUT13), .A2(n1247), .ZN(n1239) );
NAND2_X1 U905 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR3_X1 U906 ( .A1(n1243), .A2(n1242), .A3(KEYINPUT5), .ZN(n1249) );
INV_X1 U907 ( .A(G131), .ZN(n1243) );
NAND2_X1 U908 ( .A1(KEYINPUT5), .A2(n1242), .ZN(n1248) );
INV_X1 U909 ( .A(n1193), .ZN(n1242) );
NAND3_X1 U910 ( .A1(n1202), .A2(n1074), .A3(n1068), .ZN(n1193) );
INV_X1 U911 ( .A(n1228), .ZN(n1068) );
NAND2_X1 U912 ( .A1(n1061), .A2(n1250), .ZN(n1228) );
AND3_X1 U913 ( .A1(n1251), .A2(n1252), .A3(n1220), .ZN(n1202) );
XNOR2_X1 U914 ( .A(G128), .B(n1123), .ZN(G30) );
NAND3_X1 U915 ( .A1(n1215), .A2(n1075), .A3(n1220), .ZN(n1123) );
NOR2_X1 U916 ( .A1(n1083), .A2(n1253), .ZN(n1220) );
INV_X1 U917 ( .A(n1254), .ZN(n1083) );
NOR3_X1 U918 ( .A1(n1255), .A2(n1256), .A3(n1251), .ZN(n1215) );
XNOR2_X1 U919 ( .A(G101), .B(n1209), .ZN(G3) );
NAND3_X1 U920 ( .A1(n1251), .A2(n1252), .A3(n1257), .ZN(n1209) );
XNOR2_X1 U921 ( .A(G125), .B(n1258), .ZN(G27) );
NAND2_X1 U922 ( .A1(KEYINPUT1), .A2(n1199), .ZN(n1258) );
AND4_X1 U923 ( .A1(n1080), .A2(n1074), .A3(n1259), .A4(n1066), .ZN(n1199) );
NOR2_X1 U924 ( .A1(n1253), .A2(n1255), .ZN(n1259) );
AND2_X1 U925 ( .A1(n1260), .A2(n1070), .ZN(n1253) );
XOR2_X1 U926 ( .A(n1261), .B(KEYINPUT58), .Z(n1260) );
NAND3_X1 U927 ( .A1(G902), .A2(n1262), .A3(n1110), .ZN(n1261) );
NOR2_X1 U928 ( .A1(n1060), .A2(G900), .ZN(n1110) );
XNOR2_X1 U929 ( .A(G122), .B(n1210), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1056), .A2(n1214), .A3(n1067), .A4(n1263), .ZN(n1210) );
NOR2_X1 U931 ( .A1(n1203), .A2(n1264), .ZN(n1263) );
INV_X1 U932 ( .A(n1221), .ZN(n1203) );
NOR2_X1 U933 ( .A1(n1098), .A2(n1265), .ZN(n1221) );
NOR2_X1 U934 ( .A1(n1252), .A2(n1266), .ZN(n1067) );
XNOR2_X1 U935 ( .A(G119), .B(n1267), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1238), .A2(n1066), .A3(n1268), .A4(n1214), .ZN(n1267) );
XNOR2_X1 U937 ( .A(KEYINPUT51), .B(n1255), .ZN(n1268) );
INV_X1 U938 ( .A(n1264), .ZN(n1066) );
AND3_X1 U939 ( .A1(n1065), .A2(n1252), .A3(n1266), .ZN(n1238) );
XNOR2_X1 U940 ( .A(n1269), .B(n1270), .ZN(G18) );
NOR2_X1 U941 ( .A1(n1271), .A2(n1255), .ZN(n1270) );
INV_X1 U942 ( .A(n1056), .ZN(n1255) );
XOR2_X1 U943 ( .A(n1219), .B(KEYINPUT18), .Z(n1271) );
NAND3_X1 U944 ( .A1(n1075), .A2(n1214), .A3(n1081), .ZN(n1219) );
NOR2_X1 U945 ( .A1(n1272), .A2(n1265), .ZN(n1075) );
XOR2_X1 U946 ( .A(n1273), .B(n1274), .Z(G15) );
NAND2_X1 U947 ( .A1(KEYINPUT57), .A2(G113), .ZN(n1274) );
NAND2_X1 U948 ( .A1(n1056), .A2(n1275), .ZN(n1273) );
XNOR2_X1 U949 ( .A(KEYINPUT55), .B(n1218), .ZN(n1275) );
NAND3_X1 U950 ( .A1(n1074), .A2(n1214), .A3(n1081), .ZN(n1218) );
NOR3_X1 U951 ( .A1(n1266), .A2(n1256), .A3(n1264), .ZN(n1081) );
NAND2_X1 U952 ( .A1(n1086), .A2(n1276), .ZN(n1264) );
INV_X1 U953 ( .A(n1252), .ZN(n1256) );
INV_X1 U954 ( .A(n1251), .ZN(n1266) );
NOR2_X1 U955 ( .A1(n1277), .A2(n1098), .ZN(n1074) );
INV_X1 U956 ( .A(n1272), .ZN(n1098) );
XNOR2_X1 U957 ( .A(G110), .B(n1278), .ZN(G12) );
NAND2_X1 U958 ( .A1(n1080), .A2(n1257), .ZN(n1278) );
AND2_X1 U959 ( .A1(n1065), .A2(n1158), .ZN(n1257) );
AND3_X1 U960 ( .A1(n1254), .A2(n1214), .A3(n1056), .ZN(n1158) );
NOR2_X1 U961 ( .A1(n1061), .A2(n1062), .ZN(n1056) );
INV_X1 U962 ( .A(n1250), .ZN(n1062) );
NAND2_X1 U963 ( .A1(G214), .A2(n1279), .ZN(n1250) );
XNOR2_X1 U964 ( .A(n1099), .B(KEYINPUT20), .ZN(n1061) );
XNOR2_X1 U965 ( .A(n1280), .B(n1187), .ZN(n1099) );
AND2_X1 U966 ( .A1(G210), .A2(n1279), .ZN(n1187) );
NAND2_X1 U967 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
INV_X1 U968 ( .A(G237), .ZN(n1281) );
NAND2_X1 U969 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
XOR2_X1 U970 ( .A(n1285), .B(n1182), .Z(n1284) );
XOR2_X1 U971 ( .A(n1286), .B(n1140), .Z(n1182) );
XNOR2_X1 U972 ( .A(n1287), .B(G122), .ZN(n1140) );
INV_X1 U973 ( .A(G110), .ZN(n1287) );
XOR2_X1 U974 ( .A(n1288), .B(KEYINPUT52), .Z(n1286) );
NAND2_X1 U975 ( .A1(n1142), .A2(n1143), .ZN(n1288) );
NAND2_X1 U976 ( .A1(n1289), .A2(n1290), .ZN(n1143) );
XNOR2_X1 U977 ( .A(n1291), .B(n1292), .ZN(n1290) );
XOR2_X1 U978 ( .A(n1293), .B(n1294), .Z(n1289) );
NAND2_X1 U979 ( .A1(n1295), .A2(n1296), .ZN(n1142) );
XNOR2_X1 U980 ( .A(n1292), .B(n1297), .ZN(n1296) );
XNOR2_X1 U981 ( .A(n1298), .B(n1299), .ZN(n1292) );
NAND2_X1 U982 ( .A1(KEYINPUT29), .A2(n1269), .ZN(n1298) );
INV_X1 U983 ( .A(G116), .ZN(n1269) );
XNOR2_X1 U984 ( .A(n1293), .B(n1294), .ZN(n1295) );
NOR2_X1 U985 ( .A1(KEYINPUT63), .A2(G101), .ZN(n1293) );
NAND2_X1 U986 ( .A1(n1300), .A2(n1301), .ZN(n1285) );
NAND2_X1 U987 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U988 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
OR2_X1 U989 ( .A1(n1183), .A2(KEYINPUT37), .ZN(n1305) );
INV_X1 U990 ( .A(KEYINPUT41), .ZN(n1304) );
NAND2_X1 U991 ( .A1(n1183), .A2(n1306), .ZN(n1300) );
NAND2_X1 U992 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
OR2_X1 U993 ( .A1(n1302), .A2(KEYINPUT41), .ZN(n1308) );
XNOR2_X1 U994 ( .A(n1186), .B(KEYINPUT11), .ZN(n1302) );
NOR2_X1 U995 ( .A1(n1130), .A2(G953), .ZN(n1186) );
INV_X1 U996 ( .A(G224), .ZN(n1130) );
INV_X1 U997 ( .A(KEYINPUT37), .ZN(n1307) );
XOR2_X1 U998 ( .A(n1309), .B(n1119), .Z(n1183) );
NAND2_X1 U999 ( .A1(n1070), .A2(n1310), .ZN(n1214) );
NAND4_X1 U1000 ( .A1(G953), .A2(G902), .A3(n1262), .A4(n1131), .ZN(n1310) );
INV_X1 U1001 ( .A(G898), .ZN(n1131) );
NAND3_X1 U1002 ( .A1(n1262), .A2(n1060), .A3(G952), .ZN(n1070) );
NAND2_X1 U1003 ( .A1(G237), .A2(G234), .ZN(n1262) );
NOR2_X1 U1004 ( .A1(n1086), .A2(n1085), .ZN(n1254) );
INV_X1 U1005 ( .A(n1276), .ZN(n1085) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1311), .ZN(n1276) );
XNOR2_X1 U1007 ( .A(n1103), .B(n1105), .ZN(n1086) );
INV_X1 U1008 ( .A(G469), .ZN(n1105) );
NAND2_X1 U1009 ( .A1(n1312), .A2(n1283), .ZN(n1103) );
XOR2_X1 U1010 ( .A(n1313), .B(n1314), .Z(n1312) );
XOR2_X1 U1011 ( .A(KEYINPUT34), .B(n1315), .Z(n1314) );
NOR2_X1 U1012 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1013 ( .A(KEYINPUT12), .B(n1174), .Z(n1317) );
AND2_X1 U1014 ( .A1(n1176), .A2(n1318), .ZN(n1174) );
NOR2_X1 U1015 ( .A1(n1176), .A2(n1319), .ZN(n1316) );
XNOR2_X1 U1016 ( .A(KEYINPUT56), .B(n1318), .ZN(n1319) );
INV_X1 U1017 ( .A(n1178), .ZN(n1318) );
AND2_X1 U1018 ( .A1(G227), .A2(n1060), .ZN(n1176) );
XOR2_X1 U1019 ( .A(n1320), .B(n1321), .Z(n1313) );
NAND2_X1 U1020 ( .A1(KEYINPUT42), .A2(n1322), .ZN(n1320) );
XNOR2_X1 U1021 ( .A(n1119), .B(n1171), .ZN(n1322) );
XOR2_X1 U1022 ( .A(n1294), .B(n1323), .Z(n1171) );
NOR2_X1 U1023 ( .A1(G101), .A2(KEYINPUT61), .ZN(n1323) );
XOR2_X1 U1024 ( .A(G104), .B(G107), .Z(n1294) );
NOR2_X1 U1025 ( .A1(n1277), .A2(n1272), .ZN(n1065) );
XNOR2_X1 U1026 ( .A(n1324), .B(G475), .ZN(n1272) );
NAND2_X1 U1027 ( .A1(n1156), .A2(n1283), .ZN(n1324) );
XOR2_X1 U1028 ( .A(n1325), .B(n1326), .Z(n1156) );
XOR2_X1 U1029 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1030 ( .A(G146), .B(n1224), .ZN(n1328) );
XOR2_X1 U1031 ( .A(KEYINPUT60), .B(KEYINPUT23), .Z(n1327) );
XOR2_X1 U1032 ( .A(n1329), .B(n1330), .Z(n1325) );
XNOR2_X1 U1033 ( .A(n1331), .B(n1332), .ZN(n1330) );
NOR2_X1 U1034 ( .A1(n1333), .A2(KEYINPUT17), .ZN(n1332) );
NOR2_X1 U1035 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1036 ( .A(KEYINPUT24), .B(n1336), .Z(n1335) );
AND2_X1 U1037 ( .A1(n1299), .A2(n1337), .ZN(n1336) );
NOR2_X1 U1038 ( .A1(n1299), .A2(n1337), .ZN(n1334) );
XOR2_X1 U1039 ( .A(G122), .B(KEYINPUT47), .Z(n1337) );
NAND2_X1 U1040 ( .A1(KEYINPUT49), .A2(n1114), .ZN(n1331) );
XNOR2_X1 U1041 ( .A(G104), .B(n1338), .ZN(n1329) );
NOR2_X1 U1042 ( .A1(KEYINPUT19), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1043 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1044 ( .A(G143), .B(G131), .ZN(n1341) );
NAND2_X1 U1045 ( .A1(n1342), .A2(G214), .ZN(n1340) );
INV_X1 U1046 ( .A(n1265), .ZN(n1277) );
NOR2_X1 U1047 ( .A1(n1343), .A2(n1100), .ZN(n1265) );
NOR2_X1 U1048 ( .A1(n1102), .A2(G478), .ZN(n1100) );
AND2_X1 U1049 ( .A1(n1344), .A2(n1102), .ZN(n1343) );
NAND2_X1 U1050 ( .A1(n1152), .A2(n1283), .ZN(n1102) );
XOR2_X1 U1051 ( .A(n1345), .B(n1346), .Z(n1152) );
XOR2_X1 U1052 ( .A(G107), .B(n1347), .Z(n1346) );
XNOR2_X1 U1053 ( .A(n1348), .B(G116), .ZN(n1347) );
INV_X1 U1054 ( .A(G122), .ZN(n1348) );
XOR2_X1 U1055 ( .A(n1349), .B(n1350), .Z(n1345) );
NOR2_X1 U1056 ( .A1(KEYINPUT35), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1057 ( .A(G128), .B(n1352), .Z(n1351) );
XNOR2_X1 U1058 ( .A(n1353), .B(G134), .ZN(n1352) );
INV_X1 U1059 ( .A(G143), .ZN(n1353) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1354), .ZN(n1349) );
XOR2_X1 U1061 ( .A(KEYINPUT62), .B(G478), .Z(n1344) );
NOR2_X1 U1062 ( .A1(n1251), .A2(n1252), .ZN(n1080) );
XOR2_X1 U1063 ( .A(G472), .B(n1355), .Z(n1252) );
NOR2_X1 U1064 ( .A1(KEYINPUT45), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1065 ( .A(KEYINPUT25), .B(n1097), .Z(n1356) );
AND2_X1 U1066 ( .A1(n1283), .A2(n1357), .ZN(n1097) );
XOR2_X1 U1067 ( .A(n1358), .B(n1163), .Z(n1357) );
XNOR2_X1 U1068 ( .A(n1359), .B(G101), .ZN(n1163) );
NAND2_X1 U1069 ( .A1(n1342), .A2(G210), .ZN(n1359) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1342) );
NOR2_X1 U1071 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
XOR2_X1 U1072 ( .A(n1362), .B(KEYINPUT48), .Z(n1361) );
NAND2_X1 U1073 ( .A1(n1164), .A2(n1167), .ZN(n1362) );
NOR2_X1 U1074 ( .A1(n1164), .A2(n1167), .ZN(n1360) );
NAND2_X1 U1075 ( .A1(n1363), .A2(n1364), .ZN(n1167) );
NAND2_X1 U1076 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1077 ( .A1(KEYINPUT39), .A2(n1367), .ZN(n1366) );
NAND2_X1 U1078 ( .A1(KEYINPUT10), .A2(n1299), .ZN(n1367) );
INV_X1 U1079 ( .A(G113), .ZN(n1299) );
NAND2_X1 U1080 ( .A1(G113), .A2(n1368), .ZN(n1363) );
NAND2_X1 U1081 ( .A1(KEYINPUT10), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1082 ( .A1(n1370), .A2(KEYINPUT39), .ZN(n1369) );
INV_X1 U1083 ( .A(n1365), .ZN(n1370) );
XNOR2_X1 U1084 ( .A(G116), .B(n1297), .ZN(n1365) );
INV_X1 U1085 ( .A(n1291), .ZN(n1297) );
XNOR2_X1 U1086 ( .A(n1321), .B(n1119), .ZN(n1164) );
XNOR2_X1 U1087 ( .A(G143), .B(n1371), .ZN(n1119) );
XOR2_X1 U1088 ( .A(G131), .B(n1115), .Z(n1321) );
XOR2_X1 U1089 ( .A(G134), .B(G137), .Z(n1115) );
XOR2_X1 U1090 ( .A(n1093), .B(KEYINPUT40), .Z(n1251) );
XNOR2_X1 U1091 ( .A(n1372), .B(n1149), .ZN(n1093) );
AND2_X1 U1092 ( .A1(G217), .A2(n1311), .ZN(n1149) );
NAND2_X1 U1093 ( .A1(G234), .A2(n1282), .ZN(n1311) );
INV_X1 U1094 ( .A(G902), .ZN(n1282) );
NAND2_X1 U1095 ( .A1(n1283), .A2(n1147), .ZN(n1372) );
XNOR2_X1 U1096 ( .A(n1373), .B(n1374), .ZN(n1147) );
XOR2_X1 U1097 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1098 ( .A(n1377), .B(n1371), .Z(n1376) );
XOR2_X1 U1099 ( .A(G128), .B(G146), .Z(n1371) );
NAND2_X1 U1100 ( .A1(n1354), .A2(G221), .ZN(n1377) );
AND2_X1 U1101 ( .A1(G234), .A2(n1060), .ZN(n1354) );
INV_X1 U1102 ( .A(G953), .ZN(n1060) );
XNOR2_X1 U1103 ( .A(KEYINPUT23), .B(G137), .ZN(n1375) );
XNOR2_X1 U1104 ( .A(n1178), .B(n1378), .ZN(n1373) );
XNOR2_X1 U1105 ( .A(n1114), .B(n1291), .ZN(n1378) );
XOR2_X1 U1106 ( .A(G119), .B(KEYINPUT53), .Z(n1291) );
INV_X1 U1107 ( .A(n1309), .ZN(n1114) );
XOR2_X1 U1108 ( .A(G125), .B(KEYINPUT54), .Z(n1309) );
XNOR2_X1 U1109 ( .A(G110), .B(n1224), .ZN(n1178) );
INV_X1 U1110 ( .A(G140), .ZN(n1224) );
XNOR2_X1 U1111 ( .A(G902), .B(KEYINPUT14), .ZN(n1283) );
endmodule


