//Key = 1011110010001100111101001100110111001111011010000100010011111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336;

XOR2_X1 U746 ( .A(n1024), .B(G107), .Z(G9) );
NAND2_X1 U747 ( .A1(KEYINPUT28), .A2(n1025), .ZN(n1024) );
NAND2_X1 U748 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U749 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NOR2_X1 U751 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U752 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U753 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR4_X1 U754 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1046), .A2(n1027), .ZN(n1044) );
NOR2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1042) );
XOR2_X1 U759 ( .A(n1051), .B(KEYINPUT40), .Z(n1049) );
AND2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1041) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1038) );
NOR3_X1 U762 ( .A1(n1051), .A2(n1056), .A3(n1045), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR4_X1 U764 ( .A1(n1059), .A2(n1045), .A3(n1051), .A4(n1040), .ZN(n1035) );
INV_X1 U765 ( .A(n1060), .ZN(n1045) );
NOR2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U767 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U768 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1030) );
NOR4_X1 U769 ( .A1(n1067), .A2(n1068), .A3(n1051), .A4(n1069), .ZN(n1066) );
XNOR2_X1 U770 ( .A(G472), .B(n1070), .ZN(n1068) );
NOR2_X1 U771 ( .A1(n1071), .A2(KEYINPUT30), .ZN(n1070) );
XOR2_X1 U772 ( .A(n1072), .B(KEYINPUT13), .Z(n1067) );
NOR3_X1 U773 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1063) );
XOR2_X1 U775 ( .A(KEYINPUT2), .B(G469), .Z(n1077) );
XOR2_X1 U776 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U777 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U779 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U780 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND2_X1 U781 ( .A1(KEYINPUT18), .A2(n1088), .ZN(n1086) );
XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U783 ( .A(G125), .B(n1091), .Z(n1090) );
XOR2_X1 U784 ( .A(KEYINPUT49), .B(KEYINPUT41), .Z(n1089) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1080) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NAND2_X1 U787 ( .A1(G953), .A2(n1096), .ZN(n1078) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1097), .B(n1098), .Z(G69) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR3_X1 U791 ( .A1(n1101), .A2(KEYINPUT34), .A3(n1102), .ZN(n1100) );
NOR2_X1 U792 ( .A1(G898), .A2(n1103), .ZN(n1102) );
XOR2_X1 U793 ( .A(KEYINPUT26), .B(n1104), .Z(n1103) );
XOR2_X1 U794 ( .A(n1105), .B(n1106), .Z(n1101) );
XNOR2_X1 U795 ( .A(KEYINPUT4), .B(KEYINPUT24), .ZN(n1105) );
NAND2_X1 U796 ( .A1(n1093), .A2(n1107), .ZN(n1099) );
NAND2_X1 U797 ( .A1(G953), .A2(n1108), .ZN(n1097) );
NAND2_X1 U798 ( .A1(G898), .A2(G224), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(G66) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
AND2_X1 U804 ( .A1(n1116), .A2(n1115), .ZN(n1111) );
INV_X1 U805 ( .A(KEYINPUT0), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1109), .A2(n1119), .ZN(G63) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U808 ( .A1(n1117), .A2(G478), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1109), .A2(n1122), .ZN(G60) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U811 ( .A1(n1117), .A2(G475), .ZN(n1123) );
XNOR2_X1 U812 ( .A(G104), .B(n1125), .ZN(G6) );
NOR2_X1 U813 ( .A1(n1109), .A2(n1126), .ZN(G57) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U816 ( .A1(KEYINPUT62), .A2(n1131), .ZN(n1130) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U818 ( .A1(KEYINPUT39), .A2(n1134), .ZN(n1132) );
NAND2_X1 U819 ( .A1(n1117), .A2(G472), .ZN(n1129) );
NOR2_X1 U820 ( .A1(n1109), .A2(n1135), .ZN(G54) );
XOR2_X1 U821 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U822 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U823 ( .A(n1140), .B(n1141), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1117), .A2(G469), .ZN(n1140) );
INV_X1 U825 ( .A(n1142), .ZN(n1117) );
XOR2_X1 U826 ( .A(n1143), .B(n1144), .Z(n1136) );
XOR2_X1 U827 ( .A(n1145), .B(KEYINPUT22), .Z(n1144) );
NAND2_X1 U828 ( .A1(KEYINPUT17), .A2(n1146), .ZN(n1145) );
NAND2_X1 U829 ( .A1(KEYINPUT56), .A2(n1134), .ZN(n1143) );
NOR2_X1 U830 ( .A1(n1109), .A2(n1147), .ZN(G51) );
XOR2_X1 U831 ( .A(n1106), .B(n1148), .Z(n1147) );
XOR2_X1 U832 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U833 ( .A1(n1151), .A2(KEYINPUT45), .ZN(n1150) );
NOR2_X1 U834 ( .A1(n1152), .A2(n1142), .ZN(n1151) );
NAND2_X1 U835 ( .A1(G902), .A2(n1032), .ZN(n1142) );
NAND3_X1 U836 ( .A1(n1153), .A2(n1154), .A3(n1094), .ZN(n1032) );
AND4_X1 U837 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1094) );
AND4_X1 U838 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
NOR2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1157) );
NOR4_X1 U840 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1062), .ZN(n1164) );
INV_X1 U841 ( .A(KEYINPUT20), .ZN(n1165) );
NOR2_X1 U842 ( .A1(KEYINPUT20), .A2(n1168), .ZN(n1163) );
NAND2_X1 U843 ( .A1(n1053), .A2(n1169), .ZN(n1155) );
XNOR2_X1 U844 ( .A(KEYINPUT43), .B(n1170), .ZN(n1169) );
XNOR2_X1 U845 ( .A(KEYINPUT33), .B(n1095), .ZN(n1154) );
INV_X1 U846 ( .A(n1107), .ZN(n1153) );
NAND4_X1 U847 ( .A1(n1171), .A2(n1125), .A3(n1172), .A4(n1173), .ZN(n1107) );
AND3_X1 U848 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1027), .A2(n1177), .ZN(n1172) );
NAND3_X1 U850 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
XOR2_X1 U851 ( .A(KEYINPUT53), .B(n1026), .Z(n1180) );
AND3_X1 U852 ( .A1(n1060), .A2(n1061), .A3(n1181), .ZN(n1026) );
OR4_X1 U853 ( .A1(n1182), .A2(n1054), .A3(n1183), .A4(KEYINPUT37), .ZN(n1179) );
XNOR2_X1 U854 ( .A(KEYINPUT19), .B(n1184), .ZN(n1178) );
NAND4_X1 U855 ( .A1(n1062), .A2(n1027), .A3(n1181), .A4(n1060), .ZN(n1125) );
NAND2_X1 U856 ( .A1(n1185), .A2(n1186), .ZN(n1171) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U858 ( .A1(KEYINPUT37), .A2(n1189), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1062), .A2(n1190), .ZN(n1187) );
NOR3_X1 U860 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1149) );
AND3_X1 U861 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1191) );
AND2_X1 U862 ( .A1(n1197), .A2(G953), .ZN(n1109) );
XNOR2_X1 U863 ( .A(G952), .B(KEYINPUT35), .ZN(n1197) );
XOR2_X1 U864 ( .A(n1198), .B(n1156), .Z(G48) );
NAND3_X1 U865 ( .A1(n1199), .A2(n1062), .A3(n1200), .ZN(n1156) );
NAND2_X1 U866 ( .A1(n1201), .A2(n1202), .ZN(G45) );
NAND2_X1 U867 ( .A1(G143), .A2(n1162), .ZN(n1202) );
XOR2_X1 U868 ( .A(KEYINPUT31), .B(n1203), .Z(n1201) );
NOR2_X1 U869 ( .A1(G143), .A2(n1162), .ZN(n1203) );
NAND4_X1 U870 ( .A1(n1200), .A2(n1190), .A3(n1204), .A4(n1069), .ZN(n1162) );
XOR2_X1 U871 ( .A(G140), .B(n1205), .Z(G42) );
NOR2_X1 U872 ( .A1(n1051), .A2(n1170), .ZN(n1205) );
NAND3_X1 U873 ( .A1(n1206), .A2(n1052), .A3(n1062), .ZN(n1170) );
XNOR2_X1 U874 ( .A(G137), .B(n1161), .ZN(G39) );
NAND3_X1 U875 ( .A1(n1206), .A2(n1053), .A3(n1189), .ZN(n1161) );
INV_X1 U876 ( .A(n1182), .ZN(n1189) );
XOR2_X1 U877 ( .A(n1160), .B(n1207), .Z(G36) );
NOR2_X1 U878 ( .A1(G134), .A2(KEYINPUT23), .ZN(n1207) );
NAND2_X1 U879 ( .A1(n1208), .A2(n1061), .ZN(n1160) );
XNOR2_X1 U880 ( .A(G131), .B(n1159), .ZN(G33) );
NAND2_X1 U881 ( .A1(n1062), .A2(n1208), .ZN(n1159) );
AND3_X1 U882 ( .A1(n1206), .A2(n1053), .A3(n1190), .ZN(n1208) );
INV_X1 U883 ( .A(n1051), .ZN(n1053) );
NAND2_X1 U884 ( .A1(n1209), .A2(n1048), .ZN(n1051) );
INV_X1 U885 ( .A(n1210), .ZN(n1062) );
XOR2_X1 U886 ( .A(n1211), .B(n1095), .Z(G30) );
NAND3_X1 U887 ( .A1(n1199), .A2(n1061), .A3(n1200), .ZN(n1095) );
AND2_X1 U888 ( .A1(n1206), .A2(n1027), .ZN(n1200) );
NOR3_X1 U889 ( .A1(n1057), .A2(n1074), .A3(n1167), .ZN(n1206) );
XOR2_X1 U890 ( .A(n1212), .B(n1174), .Z(G3) );
NAND4_X1 U891 ( .A1(n1213), .A2(n1190), .A3(n1027), .A4(n1181), .ZN(n1174) );
XOR2_X1 U892 ( .A(n1214), .B(n1168), .Z(G27) );
OR3_X1 U893 ( .A1(n1210), .A2(n1167), .A3(n1166), .ZN(n1168) );
NAND3_X1 U894 ( .A1(n1027), .A2(n1052), .A3(n1054), .ZN(n1166) );
INV_X1 U895 ( .A(n1040), .ZN(n1054) );
INV_X1 U896 ( .A(n1215), .ZN(n1027) );
AND2_X1 U897 ( .A1(n1034), .A2(n1216), .ZN(n1167) );
NAND3_X1 U898 ( .A1(G902), .A2(n1217), .A3(n1082), .ZN(n1216) );
NOR2_X1 U899 ( .A1(n1104), .A2(G900), .ZN(n1082) );
XNOR2_X1 U900 ( .A(G122), .B(n1176), .ZN(G24) );
NAND4_X1 U901 ( .A1(n1185), .A2(n1060), .A3(n1204), .A4(n1069), .ZN(n1176) );
XOR2_X1 U902 ( .A(G119), .B(n1218), .Z(G21) );
NOR2_X1 U903 ( .A1(n1182), .A2(n1219), .ZN(n1218) );
NAND2_X1 U904 ( .A1(n1199), .A2(n1213), .ZN(n1182) );
AND2_X1 U905 ( .A1(n1220), .A2(n1221), .ZN(n1199) );
XOR2_X1 U906 ( .A(n1222), .B(n1175), .Z(G18) );
NAND3_X1 U907 ( .A1(n1190), .A2(n1061), .A3(n1185), .ZN(n1175) );
AND2_X1 U908 ( .A1(n1223), .A2(n1204), .ZN(n1061) );
XNOR2_X1 U909 ( .A(n1224), .B(KEYINPUT38), .ZN(n1204) );
INV_X1 U910 ( .A(n1050), .ZN(n1190) );
XOR2_X1 U911 ( .A(G113), .B(n1225), .Z(G15) );
NOR4_X1 U912 ( .A1(KEYINPUT9), .A2(n1050), .A3(n1210), .A4(n1219), .ZN(n1225) );
INV_X1 U913 ( .A(n1185), .ZN(n1219) );
NOR3_X1 U914 ( .A1(n1215), .A2(n1183), .A3(n1040), .ZN(n1185) );
NAND2_X1 U915 ( .A1(n1057), .A2(n1058), .ZN(n1040) );
NAND2_X1 U916 ( .A1(n1226), .A2(n1069), .ZN(n1210) );
INV_X1 U917 ( .A(n1223), .ZN(n1069) );
NAND2_X1 U918 ( .A1(n1072), .A2(n1220), .ZN(n1050) );
XOR2_X1 U919 ( .A(n1227), .B(n1228), .Z(G12) );
NOR2_X1 U920 ( .A1(KEYINPUT51), .A2(n1229), .ZN(n1228) );
NOR2_X1 U921 ( .A1(n1215), .A2(n1184), .ZN(n1227) );
NAND3_X1 U922 ( .A1(n1181), .A2(n1052), .A3(n1213), .ZN(n1184) );
INV_X1 U923 ( .A(n1037), .ZN(n1213) );
NAND2_X1 U924 ( .A1(n1223), .A2(n1226), .ZN(n1037) );
XNOR2_X1 U925 ( .A(n1224), .B(KEYINPUT50), .ZN(n1226) );
NAND2_X1 U926 ( .A1(n1230), .A2(n1064), .ZN(n1224) );
NAND3_X1 U927 ( .A1(n1231), .A2(n1232), .A3(n1121), .ZN(n1064) );
XOR2_X1 U928 ( .A(KEYINPUT5), .B(G478), .Z(n1232) );
XNOR2_X1 U929 ( .A(n1073), .B(KEYINPUT14), .ZN(n1230) );
AND2_X1 U930 ( .A1(n1233), .A2(n1234), .ZN(n1073) );
NAND2_X1 U931 ( .A1(n1121), .A2(n1231), .ZN(n1234) );
XOR2_X1 U932 ( .A(n1235), .B(n1236), .Z(n1121) );
XOR2_X1 U933 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U934 ( .A(n1239), .B(G107), .Z(n1238) );
NAND3_X1 U935 ( .A1(G234), .A2(n1093), .A3(G217), .ZN(n1239) );
NAND2_X1 U936 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
NAND2_X1 U937 ( .A1(G143), .A2(n1211), .ZN(n1241) );
XOR2_X1 U938 ( .A(KEYINPUT63), .B(n1242), .Z(n1240) );
NOR2_X1 U939 ( .A1(G143), .A2(n1211), .ZN(n1242) );
XOR2_X1 U940 ( .A(n1222), .B(n1243), .Z(n1235) );
XOR2_X1 U941 ( .A(G134), .B(G122), .Z(n1243) );
XNOR2_X1 U942 ( .A(G478), .B(KEYINPUT5), .ZN(n1233) );
XOR2_X1 U943 ( .A(n1244), .B(G475), .Z(n1223) );
NAND2_X1 U944 ( .A1(n1124), .A2(n1231), .ZN(n1244) );
XOR2_X1 U945 ( .A(n1245), .B(n1246), .Z(n1124) );
XOR2_X1 U946 ( .A(n1247), .B(n1248), .Z(n1246) );
NAND2_X1 U947 ( .A1(G214), .A2(n1249), .ZN(n1248) );
NAND3_X1 U948 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1247) );
NAND2_X1 U949 ( .A1(KEYINPUT55), .A2(n1253), .ZN(n1252) );
OR3_X1 U950 ( .A1(n1253), .A2(KEYINPUT55), .A3(n1254), .ZN(n1251) );
NAND2_X1 U951 ( .A1(n1254), .A2(n1255), .ZN(n1250) );
NAND2_X1 U952 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U953 ( .A(KEYINPUT55), .ZN(n1257) );
XNOR2_X1 U954 ( .A(KEYINPUT52), .B(n1253), .ZN(n1256) );
XNOR2_X1 U955 ( .A(n1258), .B(KEYINPUT7), .ZN(n1253) );
XOR2_X1 U956 ( .A(G113), .B(G122), .Z(n1254) );
XOR2_X1 U957 ( .A(n1259), .B(n1260), .Z(n1245) );
NOR2_X1 U958 ( .A1(KEYINPUT54), .A2(n1261), .ZN(n1260) );
XOR2_X1 U959 ( .A(n1262), .B(n1263), .Z(n1261) );
NAND2_X1 U960 ( .A1(n1264), .A2(KEYINPUT59), .ZN(n1262) );
XOR2_X1 U961 ( .A(n1265), .B(n1091), .Z(n1264) );
XNOR2_X1 U962 ( .A(KEYINPUT6), .B(n1266), .ZN(n1265) );
NOR2_X1 U963 ( .A1(KEYINPUT47), .A2(n1214), .ZN(n1266) );
XNOR2_X1 U964 ( .A(G131), .B(G143), .ZN(n1259) );
NAND2_X1 U965 ( .A1(n1267), .A2(n1268), .ZN(n1052) );
NAND2_X1 U966 ( .A1(n1060), .A2(n1269), .ZN(n1268) );
NOR2_X1 U967 ( .A1(n1221), .A2(n1220), .ZN(n1060) );
INV_X1 U968 ( .A(n1072), .ZN(n1221) );
OR3_X1 U969 ( .A1(n1072), .A2(n1220), .A3(n1269), .ZN(n1267) );
INV_X1 U970 ( .A(KEYINPUT25), .ZN(n1269) );
XOR2_X1 U971 ( .A(n1071), .B(G472), .Z(n1220) );
AND3_X1 U972 ( .A1(n1270), .A2(n1271), .A3(n1231), .ZN(n1071) );
NAND2_X1 U973 ( .A1(n1272), .A2(n1133), .ZN(n1271) );
NAND2_X1 U974 ( .A1(n1273), .A2(n1196), .ZN(n1270) );
INV_X1 U975 ( .A(n1133), .ZN(n1196) );
XNOR2_X1 U976 ( .A(n1272), .B(KEYINPUT48), .ZN(n1273) );
XNOR2_X1 U977 ( .A(n1127), .B(n1274), .ZN(n1272) );
INV_X1 U978 ( .A(n1134), .ZN(n1274) );
XOR2_X1 U979 ( .A(n1275), .B(n1276), .Z(n1127) );
XOR2_X1 U980 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U981 ( .A(KEYINPUT16), .B(KEYINPUT12), .ZN(n1278) );
XOR2_X1 U982 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U983 ( .A(n1281), .B(G116), .Z(n1279) );
NAND2_X1 U984 ( .A1(G210), .A2(n1249), .ZN(n1281) );
NOR2_X1 U985 ( .A1(G953), .A2(G237), .ZN(n1249) );
XOR2_X1 U986 ( .A(n1282), .B(n1118), .Z(n1072) );
AND2_X1 U987 ( .A1(G217), .A2(n1283), .ZN(n1118) );
NAND2_X1 U988 ( .A1(n1231), .A2(n1115), .ZN(n1282) );
NAND2_X1 U989 ( .A1(n1284), .A2(n1285), .ZN(n1115) );
NAND2_X1 U990 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U991 ( .A(n1288), .B(KEYINPUT15), .Z(n1284) );
OR2_X1 U992 ( .A1(n1287), .A2(n1286), .ZN(n1288) );
XNOR2_X1 U993 ( .A(n1289), .B(G137), .ZN(n1286) );
NAND3_X1 U994 ( .A1(G234), .A2(n1093), .A3(G221), .ZN(n1289) );
XNOR2_X1 U995 ( .A(n1290), .B(n1291), .ZN(n1287) );
XOR2_X1 U996 ( .A(n1292), .B(n1293), .Z(n1291) );
INV_X1 U997 ( .A(n1263), .ZN(n1293) );
XOR2_X1 U998 ( .A(n1198), .B(KEYINPUT44), .Z(n1263) );
INV_X1 U999 ( .A(G146), .ZN(n1198) );
NOR2_X1 U1000 ( .A1(KEYINPUT27), .A2(n1091), .ZN(n1292) );
XOR2_X1 U1001 ( .A(n1294), .B(n1295), .Z(n1290) );
XOR2_X1 U1002 ( .A(G125), .B(G110), .Z(n1295) );
NAND2_X1 U1003 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
NAND2_X1 U1004 ( .A1(G119), .A2(n1211), .ZN(n1297) );
XOR2_X1 U1005 ( .A(KEYINPUT58), .B(n1298), .Z(n1296) );
NOR2_X1 U1006 ( .A1(G119), .A2(n1211), .ZN(n1298) );
NOR3_X1 U1007 ( .A1(n1057), .A2(n1074), .A3(n1183), .ZN(n1181) );
AND2_X1 U1008 ( .A1(n1034), .A2(n1299), .ZN(n1183) );
OR4_X1 U1009 ( .A1(n1104), .A2(n1300), .A3(n1301), .A4(G898), .ZN(n1299) );
INV_X1 U1010 ( .A(n1217), .ZN(n1301) );
XNOR2_X1 U1011 ( .A(n1093), .B(KEYINPUT57), .ZN(n1104) );
NAND3_X1 U1012 ( .A1(n1217), .A2(n1093), .A3(G952), .ZN(n1034) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1217) );
INV_X1 U1014 ( .A(n1058), .ZN(n1074) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1283), .ZN(n1058) );
NAND2_X1 U1016 ( .A1(G234), .A2(n1300), .ZN(n1283) );
NOR2_X1 U1017 ( .A1(n1075), .A2(n1302), .ZN(n1057) );
AND2_X1 U1018 ( .A1(n1076), .A2(n1303), .ZN(n1302) );
NOR2_X1 U1019 ( .A1(n1303), .A2(n1076), .ZN(n1075) );
AND2_X1 U1020 ( .A1(n1231), .A2(n1304), .ZN(n1076) );
XOR2_X1 U1021 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1022 ( .A(n1138), .B(n1141), .ZN(n1306) );
XNOR2_X1 U1023 ( .A(n1229), .B(n1307), .ZN(n1141) );
AND2_X1 U1024 ( .A1(n1093), .A2(G227), .ZN(n1307) );
XNOR2_X1 U1025 ( .A(n1308), .B(n1309), .ZN(n1138) );
XOR2_X1 U1026 ( .A(KEYINPUT36), .B(G101), .Z(n1309) );
XNOR2_X1 U1027 ( .A(n1310), .B(n1087), .ZN(n1308) );
XOR2_X1 U1028 ( .A(n1134), .B(n1311), .Z(n1305) );
NOR2_X1 U1029 ( .A1(KEYINPUT11), .A2(n1091), .ZN(n1311) );
INV_X1 U1030 ( .A(n1146), .ZN(n1091) );
XNOR2_X1 U1031 ( .A(G140), .B(KEYINPUT61), .ZN(n1146) );
XNOR2_X1 U1032 ( .A(n1084), .B(KEYINPUT21), .ZN(n1134) );
XOR2_X1 U1033 ( .A(G131), .B(n1312), .Z(n1084) );
XOR2_X1 U1034 ( .A(G137), .B(G134), .Z(n1312) );
INV_X1 U1035 ( .A(G469), .ZN(n1303) );
NAND2_X1 U1036 ( .A1(n1047), .A2(n1048), .ZN(n1215) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1313), .ZN(n1048) );
INV_X1 U1038 ( .A(n1209), .ZN(n1047) );
XNOR2_X1 U1039 ( .A(n1314), .B(n1152), .ZN(n1209) );
NAND2_X1 U1040 ( .A1(G210), .A2(n1313), .ZN(n1152) );
NAND2_X1 U1041 ( .A1(n1315), .A2(n1300), .ZN(n1313) );
INV_X1 U1042 ( .A(G237), .ZN(n1315) );
NAND2_X1 U1043 ( .A1(n1316), .A2(n1231), .ZN(n1314) );
XOR2_X1 U1044 ( .A(n1300), .B(KEYINPUT10), .Z(n1231) );
INV_X1 U1045 ( .A(G902), .ZN(n1300) );
XOR2_X1 U1046 ( .A(n1317), .B(n1106), .Z(n1316) );
XNOR2_X1 U1047 ( .A(n1318), .B(n1319), .ZN(n1106) );
XNOR2_X1 U1048 ( .A(n1320), .B(n1280), .ZN(n1319) );
XNOR2_X1 U1049 ( .A(n1212), .B(G113), .ZN(n1280) );
INV_X1 U1050 ( .A(G101), .ZN(n1212) );
NAND3_X1 U1051 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(n1320) );
OR2_X1 U1052 ( .A1(n1222), .A2(KEYINPUT32), .ZN(n1323) );
NAND3_X1 U1053 ( .A1(KEYINPUT32), .A2(n1222), .A3(G119), .ZN(n1322) );
INV_X1 U1054 ( .A(G116), .ZN(n1222) );
NAND2_X1 U1055 ( .A1(n1324), .A2(n1277), .ZN(n1321) );
INV_X1 U1056 ( .A(G119), .ZN(n1277) );
NAND2_X1 U1057 ( .A1(KEYINPUT32), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1058 ( .A(KEYINPUT8), .B(G116), .Z(n1325) );
XOR2_X1 U1059 ( .A(n1326), .B(n1327), .Z(n1318) );
NOR2_X1 U1060 ( .A1(KEYINPUT46), .A2(n1310), .ZN(n1327) );
XNOR2_X1 U1061 ( .A(n1328), .B(n1258), .ZN(n1310) );
XOR2_X1 U1062 ( .A(G104), .B(KEYINPUT3), .Z(n1258) );
INV_X1 U1063 ( .A(G107), .ZN(n1328) );
XOR2_X1 U1064 ( .A(n1229), .B(G122), .Z(n1326) );
INV_X1 U1065 ( .A(G110), .ZN(n1229) );
XOR2_X1 U1066 ( .A(n1329), .B(KEYINPUT42), .Z(n1317) );
NAND4_X1 U1067 ( .A1(n1330), .A2(n1331), .A3(n1332), .A4(n1333), .ZN(n1329) );
OR3_X1 U1068 ( .A1(n1195), .A2(KEYINPUT29), .A3(n1194), .ZN(n1333) );
NAND3_X1 U1069 ( .A1(n1334), .A2(n1195), .A3(n1194), .ZN(n1332) );
NAND2_X1 U1070 ( .A1(KEYINPUT29), .A2(n1133), .ZN(n1334) );
INV_X1 U1071 ( .A(n1193), .ZN(n1331) );
NOR3_X1 U1072 ( .A1(n1194), .A2(n1133), .A3(n1195), .ZN(n1193) );
NAND2_X1 U1073 ( .A1(n1192), .A2(KEYINPUT29), .ZN(n1330) );
AND2_X1 U1074 ( .A1(n1335), .A2(n1133), .ZN(n1192) );
XNOR2_X1 U1075 ( .A(n1087), .B(KEYINPUT1), .ZN(n1133) );
XNOR2_X1 U1076 ( .A(n1211), .B(n1336), .ZN(n1087) );
XOR2_X1 U1077 ( .A(G146), .B(G143), .Z(n1336) );
INV_X1 U1078 ( .A(G128), .ZN(n1211) );
XOR2_X1 U1079 ( .A(n1195), .B(n1194), .Z(n1335) );
XNOR2_X1 U1080 ( .A(n1214), .B(KEYINPUT60), .ZN(n1194) );
INV_X1 U1081 ( .A(G125), .ZN(n1214) );
NAND2_X1 U1082 ( .A1(G224), .A2(n1093), .ZN(n1195) );
INV_X1 U1083 ( .A(G953), .ZN(n1093) );
endmodule


