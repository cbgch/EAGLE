//Key = 0011000100110001010101110011110001101101100100001000001010101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395;

XOR2_X1 U756 ( .A(n1050), .B(n1051), .Z(G9) );
NAND4_X1 U757 ( .A1(KEYINPUT26), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1051) );
NOR2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U759 ( .A1(G953), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1056) );
NOR2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U763 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1064) );
AND3_X1 U764 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT63), .ZN(n1068) );
NOR2_X1 U765 ( .A1(n1071), .A2(n1069), .ZN(n1067) );
NOR3_X1 U766 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1052), .A2(n1077), .ZN(n1075) );
AND3_X1 U769 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1073) );
NOR2_X1 U770 ( .A1(KEYINPUT63), .A2(n1081), .ZN(n1072) );
NOR3_X1 U771 ( .A1(n1082), .A2(n1083), .A3(n1076), .ZN(n1066) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR4_X1 U774 ( .A1(n1088), .A2(n1076), .A3(n1082), .A4(n1069), .ZN(n1062) );
NOR2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U776 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1055) );
AND4_X1 U777 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1057) );
NOR4_X1 U778 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
INV_X1 U779 ( .A(n1087), .ZN(n1097) );
NOR3_X1 U780 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1093) );
NOR2_X1 U781 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U782 ( .A(KEYINPUT41), .ZN(n1103) );
NOR3_X1 U783 ( .A1(n1104), .A2(n1078), .A3(n1105), .ZN(n1102) );
NOR2_X1 U784 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
INV_X1 U785 ( .A(G469), .ZN(n1104) );
NOR2_X1 U786 ( .A1(KEYINPUT41), .A2(n1108), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1109), .B(n1110), .Z(n1099) );
XOR2_X1 U788 ( .A(n1111), .B(n1112), .Z(n1091) );
XOR2_X1 U789 ( .A(n1113), .B(n1114), .Z(G72) );
NOR2_X1 U790 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1117), .B(KEYINPUT57), .Z(n1116) );
NOR2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U793 ( .A1(n1120), .A2(n1121), .ZN(n1113) );
NAND3_X1 U794 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
INV_X1 U795 ( .A(n1125), .ZN(n1124) );
NAND2_X1 U796 ( .A1(G953), .A2(n1119), .ZN(n1123) );
NAND2_X1 U797 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
XOR2_X1 U798 ( .A(n1128), .B(KEYINPUT5), .Z(n1120) );
NAND3_X1 U799 ( .A1(n1126), .A2(n1127), .A3(n1125), .ZN(n1128) );
XOR2_X1 U800 ( .A(n1129), .B(n1130), .Z(n1125) );
XOR2_X1 U801 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND2_X1 U802 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U803 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U804 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U805 ( .A1(KEYINPUT36), .A2(G134), .ZN(n1138) );
NAND2_X1 U806 ( .A1(n1139), .A2(n1140), .ZN(n1133) );
NAND2_X1 U807 ( .A1(KEYINPUT36), .A2(n1141), .ZN(n1139) );
NAND2_X1 U808 ( .A1(n1142), .A2(n1137), .ZN(n1141) );
INV_X1 U809 ( .A(KEYINPUT1), .ZN(n1137) );
XNOR2_X1 U810 ( .A(n1143), .B(n1144), .ZN(n1129) );
NAND2_X1 U811 ( .A1(n1145), .A2(n1146), .ZN(n1126) );
XOR2_X1 U812 ( .A(n1147), .B(KEYINPUT31), .Z(n1145) );
XOR2_X1 U813 ( .A(n1148), .B(n1149), .Z(G69) );
XOR2_X1 U814 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U815 ( .A1(n1152), .A2(G953), .ZN(n1151) );
NOR3_X1 U816 ( .A1(n1153), .A2(KEYINPUT44), .A3(n1154), .ZN(n1150) );
NOR2_X1 U817 ( .A1(G898), .A2(n1127), .ZN(n1154) );
NAND3_X1 U818 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1153) );
NAND2_X1 U819 ( .A1(KEYINPUT24), .A2(n1158), .ZN(n1157) );
OR3_X1 U820 ( .A1(n1158), .A2(KEYINPUT24), .A3(n1159), .ZN(n1156) );
NAND2_X1 U821 ( .A1(n1159), .A2(n1160), .ZN(n1155) );
NAND2_X1 U822 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
INV_X1 U823 ( .A(KEYINPUT24), .ZN(n1162) );
XNOR2_X1 U824 ( .A(n1158), .B(KEYINPUT6), .ZN(n1161) );
INV_X1 U825 ( .A(n1163), .ZN(n1159) );
NOR2_X1 U826 ( .A1(n1164), .A2(n1117), .ZN(n1148) );
XOR2_X1 U827 ( .A(n1127), .B(KEYINPUT32), .Z(n1117) );
NOR2_X1 U828 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NOR2_X1 U829 ( .A1(n1167), .A2(n1168), .ZN(G66) );
XNOR2_X1 U830 ( .A(n1169), .B(n1170), .ZN(n1168) );
NOR3_X1 U831 ( .A1(n1171), .A2(KEYINPUT59), .A3(n1172), .ZN(n1170) );
NOR2_X1 U832 ( .A1(n1167), .A2(n1173), .ZN(G63) );
XOR2_X1 U833 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U834 ( .A1(n1112), .A2(n1171), .ZN(n1174) );
NOR2_X1 U835 ( .A1(n1167), .A2(n1176), .ZN(G60) );
NOR2_X1 U836 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U837 ( .A(KEYINPUT0), .B(n1179), .Z(n1178) );
AND2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U839 ( .A1(n1181), .A2(n1180), .ZN(n1177) );
NAND3_X1 U840 ( .A1(n1182), .A2(n1059), .A3(G475), .ZN(n1180) );
XOR2_X1 U841 ( .A(KEYINPUT13), .B(G902), .Z(n1182) );
XNOR2_X1 U842 ( .A(n1183), .B(n1184), .ZN(G6) );
NAND2_X1 U843 ( .A1(KEYINPUT2), .A2(G104), .ZN(n1184) );
NOR2_X1 U844 ( .A1(n1167), .A2(n1185), .ZN(G57) );
XOR2_X1 U845 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U846 ( .A(KEYINPUT60), .B(G101), .Z(n1187) );
XNOR2_X1 U847 ( .A(n1188), .B(n1189), .ZN(n1186) );
NAND2_X1 U848 ( .A1(KEYINPUT39), .A2(n1190), .ZN(n1189) );
NAND2_X1 U849 ( .A1(n1191), .A2(KEYINPUT58), .ZN(n1188) );
XOR2_X1 U850 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U851 ( .A(n1194), .B(n1195), .Z(n1192) );
NOR2_X1 U852 ( .A1(n1196), .A2(n1171), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1167), .A2(n1197), .ZN(G54) );
XOR2_X1 U854 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U855 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U856 ( .A1(n1171), .A2(n1202), .ZN(n1201) );
XOR2_X1 U857 ( .A(KEYINPUT21), .B(G469), .Z(n1202) );
NOR2_X1 U858 ( .A1(KEYINPUT45), .A2(n1203), .ZN(n1200) );
XNOR2_X1 U859 ( .A(n1204), .B(n1205), .ZN(n1203) );
XOR2_X1 U860 ( .A(n1206), .B(n1207), .Z(n1198) );
NOR2_X1 U861 ( .A1(G140), .A2(KEYINPUT46), .ZN(n1207) );
NOR2_X1 U862 ( .A1(n1167), .A2(n1208), .ZN(G51) );
XOR2_X1 U863 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U864 ( .A1(n1109), .A2(n1171), .ZN(n1210) );
NAND2_X1 U865 ( .A1(G902), .A2(n1059), .ZN(n1171) );
NAND3_X1 U866 ( .A1(n1146), .A2(n1147), .A3(n1152), .ZN(n1059) );
AND4_X1 U867 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1152) );
NOR4_X1 U868 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR2_X1 U869 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U870 ( .A1(n1221), .A2(n1222), .ZN(n1217) );
XOR2_X1 U871 ( .A(n1223), .B(KEYINPUT50), .Z(n1221) );
NOR2_X1 U872 ( .A1(n1224), .A2(n1065), .ZN(n1216) );
NOR2_X1 U873 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
AND2_X1 U874 ( .A1(n1054), .A2(n1052), .ZN(n1226) );
INV_X1 U875 ( .A(n1227), .ZN(n1054) );
NOR4_X1 U876 ( .A1(n1228), .A2(n1076), .A3(n1229), .A4(n1230), .ZN(n1225) );
NAND3_X1 U877 ( .A1(n1222), .A2(n1220), .A3(n1231), .ZN(n1228) );
INV_X1 U878 ( .A(KEYINPUT54), .ZN(n1220) );
NOR4_X1 U879 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1215) );
NOR2_X1 U880 ( .A1(n1236), .A2(n1237), .ZN(n1233) );
NOR2_X1 U881 ( .A1(n1238), .A2(n1085), .ZN(n1236) );
NOR2_X1 U882 ( .A1(n1239), .A2(n1240), .ZN(n1232) );
NOR2_X1 U883 ( .A1(n1076), .A2(n1237), .ZN(n1240) );
INV_X1 U884 ( .A(KEYINPUT47), .ZN(n1237) );
NOR2_X1 U885 ( .A1(n1183), .A2(n1241), .ZN(n1213) );
NOR3_X1 U886 ( .A1(n1065), .A2(n1227), .A3(n1235), .ZN(n1183) );
INV_X1 U887 ( .A(n1053), .ZN(n1065) );
NAND3_X1 U888 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1147) );
XOR2_X1 U889 ( .A(n1069), .B(KEYINPUT28), .Z(n1244) );
AND4_X1 U890 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1146) );
AND4_X1 U891 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1248) );
NAND2_X1 U892 ( .A1(KEYINPUT22), .A2(n1253), .ZN(n1209) );
XOR2_X1 U893 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND3_X1 U894 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1254) );
OR2_X1 U895 ( .A1(n1259), .A2(G125), .ZN(n1258) );
NAND2_X1 U896 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
INV_X1 U897 ( .A(KEYINPUT62), .ZN(n1261) );
NAND2_X1 U898 ( .A1(n1262), .A2(n1259), .ZN(n1260) );
XOR2_X1 U899 ( .A(KEYINPUT19), .B(n1131), .Z(n1262) );
NAND2_X1 U900 ( .A1(KEYINPUT62), .A2(n1263), .ZN(n1256) );
NAND2_X1 U901 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
OR2_X1 U902 ( .A1(G125), .A2(KEYINPUT19), .ZN(n1265) );
NAND3_X1 U903 ( .A1(G125), .A2(n1259), .A3(KEYINPUT19), .ZN(n1264) );
AND2_X1 U904 ( .A1(n1266), .A2(G953), .ZN(n1167) );
XNOR2_X1 U905 ( .A(G952), .B(KEYINPUT55), .ZN(n1266) );
XOR2_X1 U906 ( .A(n1245), .B(n1267), .Z(G48) );
NAND2_X1 U907 ( .A1(KEYINPUT17), .A2(G146), .ZN(n1267) );
NAND3_X1 U908 ( .A1(n1077), .A2(n1085), .A3(n1268), .ZN(n1245) );
XNOR2_X1 U909 ( .A(G143), .B(n1246), .ZN(G45) );
NAND4_X1 U910 ( .A1(n1269), .A2(n1085), .A3(n1270), .A4(n1098), .ZN(n1246) );
XOR2_X1 U911 ( .A(n1271), .B(n1272), .Z(G42) );
NAND4_X1 U912 ( .A1(KEYINPUT34), .A2(n1242), .A3(n1273), .A4(n1243), .ZN(n1272) );
XNOR2_X1 U913 ( .A(G137), .B(n1252), .ZN(G39) );
NAND3_X1 U914 ( .A1(n1268), .A2(n1079), .A3(n1273), .ZN(n1252) );
XOR2_X1 U915 ( .A(n1140), .B(n1251), .Z(G36) );
NAND3_X1 U916 ( .A1(n1269), .A2(n1052), .A3(n1273), .ZN(n1251) );
XNOR2_X1 U917 ( .A(G131), .B(n1250), .ZN(G33) );
NAND3_X1 U918 ( .A1(n1269), .A2(n1077), .A3(n1273), .ZN(n1250) );
INV_X1 U919 ( .A(n1069), .ZN(n1273) );
NAND2_X1 U920 ( .A1(n1274), .A2(n1087), .ZN(n1069) );
AND3_X1 U921 ( .A1(n1243), .A2(n1275), .A3(n1090), .ZN(n1269) );
XOR2_X1 U922 ( .A(n1276), .B(n1249), .Z(G30) );
NAND3_X1 U923 ( .A1(n1052), .A2(n1085), .A3(n1268), .ZN(n1249) );
AND4_X1 U924 ( .A1(n1243), .A2(n1277), .A3(n1275), .A4(n1278), .ZN(n1268) );
NAND2_X1 U925 ( .A1(n1279), .A2(n1280), .ZN(G3) );
OR2_X1 U926 ( .A1(n1281), .A2(n1241), .ZN(n1280) );
XOR2_X1 U927 ( .A(n1282), .B(KEYINPUT53), .Z(n1279) );
NAND2_X1 U928 ( .A1(n1241), .A2(n1281), .ZN(n1282) );
NOR3_X1 U929 ( .A1(n1234), .A2(n1227), .A3(n1082), .ZN(n1241) );
NAND3_X1 U930 ( .A1(n1085), .A2(n1231), .A3(n1243), .ZN(n1227) );
XOR2_X1 U931 ( .A(n1283), .B(G125), .Z(G27) );
NAND2_X1 U932 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND4_X1 U933 ( .A1(n1286), .A2(n1089), .A3(n1287), .A4(n1288), .ZN(n1285) );
NOR3_X1 U934 ( .A1(n1235), .A2(n1222), .A3(n1076), .ZN(n1287) );
INV_X1 U935 ( .A(n1275), .ZN(n1286) );
OR2_X1 U936 ( .A1(n1247), .A2(n1288), .ZN(n1284) );
INV_X1 U937 ( .A(KEYINPUT29), .ZN(n1288) );
NAND3_X1 U938 ( .A1(n1108), .A2(n1085), .A3(n1242), .ZN(n1247) );
AND3_X1 U939 ( .A1(n1077), .A2(n1275), .A3(n1089), .ZN(n1242) );
NAND2_X1 U940 ( .A1(n1061), .A2(n1289), .ZN(n1275) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1290), .A4(n1119), .ZN(n1289) );
INV_X1 U942 ( .A(G900), .ZN(n1119) );
INV_X1 U943 ( .A(n1222), .ZN(n1085) );
INV_X1 U944 ( .A(n1076), .ZN(n1108) );
XOR2_X1 U945 ( .A(n1291), .B(n1219), .Z(G24) );
NAND4_X1 U946 ( .A1(n1239), .A2(n1053), .A3(n1270), .A4(n1098), .ZN(n1219) );
NOR2_X1 U947 ( .A1(n1278), .A2(n1277), .ZN(n1053) );
XNOR2_X1 U948 ( .A(G119), .B(n1211), .ZN(G21) );
NAND4_X1 U949 ( .A1(n1079), .A2(n1239), .A3(n1277), .A4(n1278), .ZN(n1211) );
INV_X1 U950 ( .A(n1292), .ZN(n1277) );
XNOR2_X1 U951 ( .A(G116), .B(n1212), .ZN(G18) );
NAND3_X1 U952 ( .A1(n1239), .A2(n1052), .A3(n1090), .ZN(n1212) );
NOR2_X1 U953 ( .A1(n1098), .A2(n1230), .ZN(n1052) );
XNOR2_X1 U954 ( .A(G113), .B(n1293), .ZN(G15) );
NAND4_X1 U955 ( .A1(KEYINPUT15), .A2(n1090), .A3(n1239), .A4(n1294), .ZN(n1293) );
XOR2_X1 U956 ( .A(KEYINPUT38), .B(n1077), .Z(n1294) );
INV_X1 U957 ( .A(n1235), .ZN(n1077) );
NAND2_X1 U958 ( .A1(n1230), .A2(n1098), .ZN(n1235) );
INV_X1 U959 ( .A(n1229), .ZN(n1098) );
NOR3_X1 U960 ( .A1(n1222), .A2(n1238), .A3(n1076), .ZN(n1239) );
NAND2_X1 U961 ( .A1(n1080), .A2(n1295), .ZN(n1076) );
INV_X1 U962 ( .A(n1231), .ZN(n1238) );
INV_X1 U963 ( .A(n1234), .ZN(n1090) );
NAND2_X1 U964 ( .A1(n1292), .A2(n1278), .ZN(n1234) );
XOR2_X1 U965 ( .A(G110), .B(n1296), .Z(G12) );
NOR2_X1 U966 ( .A1(n1222), .A2(n1223), .ZN(n1296) );
NAND3_X1 U967 ( .A1(n1089), .A2(n1231), .A3(n1070), .ZN(n1223) );
INV_X1 U968 ( .A(n1081), .ZN(n1070) );
NAND2_X1 U969 ( .A1(n1079), .A2(n1243), .ZN(n1081) );
NOR2_X1 U970 ( .A1(n1080), .A2(n1078), .ZN(n1243) );
INV_X1 U971 ( .A(n1295), .ZN(n1078) );
NAND2_X1 U972 ( .A1(G221), .A2(n1297), .ZN(n1295) );
XOR2_X1 U973 ( .A(n1298), .B(G469), .Z(n1080) );
OR2_X1 U974 ( .A1(n1107), .A2(n1106), .ZN(n1298) );
XNOR2_X1 U975 ( .A(n1299), .B(n1143), .ZN(n1107) );
XNOR2_X1 U976 ( .A(n1205), .B(G140), .ZN(n1143) );
NAND2_X1 U977 ( .A1(KEYINPUT11), .A2(n1300), .ZN(n1205) );
XOR2_X1 U978 ( .A(n1204), .B(n1301), .Z(n1299) );
INV_X1 U979 ( .A(n1206), .ZN(n1301) );
XOR2_X1 U980 ( .A(n1302), .B(n1303), .Z(n1206) );
NOR2_X1 U981 ( .A1(G953), .A2(n1118), .ZN(n1303) );
INV_X1 U982 ( .A(G227), .ZN(n1118) );
XOR2_X1 U983 ( .A(n1304), .B(n1305), .Z(n1204) );
INV_X1 U984 ( .A(n1082), .ZN(n1079) );
NAND2_X1 U985 ( .A1(n1229), .A2(n1230), .ZN(n1082) );
INV_X1 U986 ( .A(n1270), .ZN(n1230) );
XOR2_X1 U987 ( .A(n1306), .B(n1111), .Z(n1270) );
NOR2_X1 U988 ( .A1(n1175), .A2(n1106), .ZN(n1111) );
INV_X1 U989 ( .A(n1307), .ZN(n1106) );
XNOR2_X1 U990 ( .A(n1308), .B(n1309), .ZN(n1175) );
NOR2_X1 U991 ( .A1(n1310), .A2(n1172), .ZN(n1309) );
INV_X1 U992 ( .A(G217), .ZN(n1172) );
NAND2_X1 U993 ( .A1(n1311), .A2(KEYINPUT7), .ZN(n1308) );
XOR2_X1 U994 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U995 ( .A(G107), .B(n1314), .Z(n1313) );
NOR2_X1 U996 ( .A1(KEYINPUT12), .A2(n1315), .ZN(n1314) );
XOR2_X1 U997 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U998 ( .A(n1276), .B(G134), .Z(n1316) );
XOR2_X1 U999 ( .A(G116), .B(n1291), .Z(n1312) );
NAND2_X1 U1000 ( .A1(KEYINPUT48), .A2(n1112), .ZN(n1306) );
INV_X1 U1001 ( .A(G478), .ZN(n1112) );
XOR2_X1 U1002 ( .A(n1318), .B(G475), .Z(n1229) );
NAND2_X1 U1003 ( .A1(n1307), .A2(n1181), .ZN(n1318) );
XOR2_X1 U1004 ( .A(n1319), .B(n1320), .Z(n1181) );
XOR2_X1 U1005 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1006 ( .A(G122), .B(G113), .Z(n1322) );
XOR2_X1 U1007 ( .A(G146), .B(G131), .Z(n1321) );
XOR2_X1 U1008 ( .A(n1323), .B(n1324), .Z(n1319) );
XOR2_X1 U1009 ( .A(n1325), .B(n1317), .Z(n1324) );
AND3_X1 U1010 ( .A1(G214), .A2(n1127), .A3(n1326), .ZN(n1325) );
XOR2_X1 U1011 ( .A(n1327), .B(G104), .Z(n1323) );
NAND3_X1 U1012 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1013 ( .A1(KEYINPUT14), .A2(G140), .ZN(n1330) );
NAND3_X1 U1014 ( .A1(n1271), .A2(n1331), .A3(G125), .ZN(n1329) );
NAND2_X1 U1015 ( .A1(n1332), .A2(n1131), .ZN(n1328) );
NAND2_X1 U1016 ( .A1(n1333), .A2(n1331), .ZN(n1332) );
INV_X1 U1017 ( .A(KEYINPUT14), .ZN(n1331) );
XOR2_X1 U1018 ( .A(n1271), .B(KEYINPUT51), .Z(n1333) );
INV_X1 U1019 ( .A(G140), .ZN(n1271) );
NAND2_X1 U1020 ( .A1(n1334), .A2(n1335), .ZN(n1231) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1290), .A4(n1166), .ZN(n1335) );
INV_X1 U1022 ( .A(G898), .ZN(n1166) );
XOR2_X1 U1023 ( .A(n1061), .B(KEYINPUT16), .Z(n1334) );
NAND3_X1 U1024 ( .A1(n1290), .A2(n1127), .A3(G952), .ZN(n1061) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1290) );
NOR2_X1 U1026 ( .A1(n1278), .A2(n1292), .ZN(n1089) );
XOR2_X1 U1027 ( .A(n1092), .B(KEYINPUT30), .Z(n1292) );
XOR2_X1 U1028 ( .A(n1336), .B(n1337), .Z(n1092) );
AND2_X1 U1029 ( .A1(n1297), .A2(G217), .ZN(n1337) );
NAND2_X1 U1030 ( .A1(G234), .A2(n1338), .ZN(n1297) );
NAND2_X1 U1031 ( .A1(n1307), .A2(n1169), .ZN(n1336) );
XNOR2_X1 U1032 ( .A(n1339), .B(n1340), .ZN(n1169) );
XOR2_X1 U1033 ( .A(n1341), .B(n1135), .Z(n1340) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1342), .ZN(n1341) );
INV_X1 U1035 ( .A(n1310), .ZN(n1342) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1127), .ZN(n1310) );
XOR2_X1 U1037 ( .A(n1343), .B(n1344), .Z(n1339) );
NOR2_X1 U1038 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1039 ( .A(n1347), .B(KEYINPUT3), .Z(n1346) );
NAND2_X1 U1040 ( .A1(G119), .A2(n1276), .ZN(n1347) );
NOR2_X1 U1041 ( .A1(G119), .A2(n1276), .ZN(n1345) );
INV_X1 U1042 ( .A(G128), .ZN(n1276) );
XOR2_X1 U1043 ( .A(n1348), .B(G110), .Z(n1343) );
NAND2_X1 U1044 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1045 ( .A1(G146), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1046 ( .A(KEYINPUT27), .B(n1352), .Z(n1349) );
NOR2_X1 U1047 ( .A1(G146), .A2(n1351), .ZN(n1352) );
XOR2_X1 U1048 ( .A(G140), .B(G125), .Z(n1351) );
NAND3_X1 U1049 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1278) );
INV_X1 U1050 ( .A(n1095), .ZN(n1355) );
NOR2_X1 U1051 ( .A1(n1356), .A2(G472), .ZN(n1095) );
NAND2_X1 U1052 ( .A1(KEYINPUT61), .A2(n1196), .ZN(n1354) );
INV_X1 U1053 ( .A(G472), .ZN(n1196) );
NAND2_X1 U1054 ( .A1(n1096), .A2(n1357), .ZN(n1353) );
INV_X1 U1055 ( .A(KEYINPUT61), .ZN(n1357) );
AND2_X1 U1056 ( .A1(G472), .A2(n1356), .ZN(n1096) );
NAND2_X1 U1057 ( .A1(n1307), .A2(n1358), .ZN(n1356) );
XNOR2_X1 U1058 ( .A(n1193), .B(n1359), .ZN(n1358) );
XNOR2_X1 U1059 ( .A(n1305), .B(n1190), .ZN(n1359) );
AND3_X1 U1060 ( .A1(n1326), .A2(n1127), .A3(G210), .ZN(n1190) );
INV_X1 U1061 ( .A(G953), .ZN(n1127) );
XOR2_X1 U1062 ( .A(n1281), .B(n1194), .Z(n1305) );
XOR2_X1 U1063 ( .A(n1360), .B(n1144), .Z(n1194) );
XOR2_X1 U1064 ( .A(G131), .B(n1361), .Z(n1144) );
NAND2_X1 U1065 ( .A1(n1362), .A2(KEYINPUT56), .ZN(n1360) );
XOR2_X1 U1066 ( .A(n1140), .B(n1142), .Z(n1362) );
INV_X1 U1067 ( .A(n1135), .ZN(n1142) );
XNOR2_X1 U1068 ( .A(G137), .B(KEYINPUT33), .ZN(n1135) );
INV_X1 U1069 ( .A(G134), .ZN(n1140) );
XOR2_X1 U1070 ( .A(n1363), .B(n1364), .Z(n1193) );
NAND2_X1 U1071 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
NAND2_X1 U1072 ( .A1(G113), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1073 ( .A(KEYINPUT40), .B(n1368), .Z(n1365) );
NOR2_X1 U1074 ( .A1(G113), .A2(n1367), .ZN(n1368) );
NAND2_X1 U1075 ( .A1(n1086), .A2(n1087), .ZN(n1222) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1369), .ZN(n1087) );
INV_X1 U1077 ( .A(n1274), .ZN(n1086) );
XOR2_X1 U1078 ( .A(n1109), .B(n1370), .Z(n1274) );
NOR2_X1 U1079 ( .A1(KEYINPUT8), .A2(n1110), .ZN(n1370) );
NAND2_X1 U1080 ( .A1(n1371), .A2(n1307), .ZN(n1110) );
XOR2_X1 U1081 ( .A(n1338), .B(KEYINPUT35), .Z(n1307) );
XOR2_X1 U1082 ( .A(n1255), .B(n1372), .Z(n1371) );
NOR2_X1 U1083 ( .A1(KEYINPUT18), .A2(n1373), .ZN(n1372) );
XOR2_X1 U1084 ( .A(n1131), .B(n1374), .Z(n1373) );
NAND2_X1 U1085 ( .A1(KEYINPUT43), .A2(n1259), .ZN(n1374) );
XOR2_X1 U1086 ( .A(n1364), .B(n1361), .Z(n1259) );
XOR2_X1 U1087 ( .A(G128), .B(G146), .Z(n1361) );
NAND2_X1 U1088 ( .A1(KEYINPUT37), .A2(n1317), .ZN(n1364) );
INV_X1 U1089 ( .A(n1300), .ZN(n1317) );
XNOR2_X1 U1090 ( .A(G143), .B(KEYINPUT25), .ZN(n1300) );
INV_X1 U1091 ( .A(G125), .ZN(n1131) );
XNOR2_X1 U1092 ( .A(n1158), .B(n1375), .ZN(n1255) );
XOR2_X1 U1093 ( .A(n1376), .B(n1377), .Z(n1375) );
NOR2_X1 U1094 ( .A1(KEYINPUT4), .A2(n1163), .ZN(n1377) );
XOR2_X1 U1095 ( .A(n1378), .B(n1379), .Z(n1163) );
NOR3_X1 U1096 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1379) );
NOR2_X1 U1097 ( .A1(n1383), .A2(n1367), .ZN(n1382) );
AND3_X1 U1098 ( .A1(n1367), .A2(n1384), .A3(n1383), .ZN(n1381) );
AND2_X1 U1099 ( .A1(KEYINPUT23), .A2(n1385), .ZN(n1383) );
XOR2_X1 U1100 ( .A(G116), .B(G119), .Z(n1367) );
NOR2_X1 U1101 ( .A1(n1385), .A2(n1384), .ZN(n1380) );
INV_X1 U1102 ( .A(KEYINPUT49), .ZN(n1384) );
XOR2_X1 U1103 ( .A(G113), .B(KEYINPUT10), .Z(n1385) );
NAND2_X1 U1104 ( .A1(n1386), .A2(n1387), .ZN(n1378) );
NAND2_X1 U1105 ( .A1(n1388), .A2(n1281), .ZN(n1387) );
INV_X1 U1106 ( .A(G101), .ZN(n1281) );
XOR2_X1 U1107 ( .A(n1389), .B(KEYINPUT52), .Z(n1386) );
NAND2_X1 U1108 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
XOR2_X1 U1109 ( .A(KEYINPUT20), .B(G101), .Z(n1391) );
INV_X1 U1110 ( .A(n1388), .ZN(n1390) );
NAND2_X1 U1111 ( .A1(n1392), .A2(n1393), .ZN(n1388) );
NAND2_X1 U1112 ( .A1(n1304), .A2(n1394), .ZN(n1393) );
INV_X1 U1113 ( .A(KEYINPUT9), .ZN(n1394) );
XOR2_X1 U1114 ( .A(n1050), .B(n1395), .Z(n1304) );
NAND3_X1 U1115 ( .A1(n1395), .A2(n1050), .A3(KEYINPUT9), .ZN(n1392) );
INV_X1 U1116 ( .A(G107), .ZN(n1050) );
XOR2_X1 U1117 ( .A(G104), .B(KEYINPUT42), .Z(n1395) );
NOR2_X1 U1118 ( .A1(G953), .A2(n1165), .ZN(n1376) );
INV_X1 U1119 ( .A(G224), .ZN(n1165) );
XOR2_X1 U1120 ( .A(n1302), .B(n1291), .Z(n1158) );
INV_X1 U1121 ( .A(G122), .ZN(n1291) );
INV_X1 U1122 ( .A(G110), .ZN(n1302) );
NAND2_X1 U1123 ( .A1(G210), .A2(n1369), .ZN(n1109) );
NAND2_X1 U1124 ( .A1(n1326), .A2(n1338), .ZN(n1369) );
INV_X1 U1125 ( .A(G902), .ZN(n1338) );
INV_X1 U1126 ( .A(G237), .ZN(n1326) );
endmodule


