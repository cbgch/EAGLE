//Key = 11100111111100001110110101100101
module c1355 ( G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, 
        G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, 
        G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, 
        G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, 
        G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, 
        G233gat, G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, 
        G1330gat, G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, 
        G1337gat, G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, 
        G1344gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, 
        G1351gat, G1352gat, G1353gat, G1354gat, G1355gat, KEYINPUT0, KEYINPUT1, 
        KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, 
        KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, 
        KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, 
        KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, 
        KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31
 );
  input G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
         G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
         G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
         G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
         G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat,
         G231gat, G232gat, G233gat, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3,
         KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9,
         KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
         KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
         KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
         KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
         KEYINPUT30, KEYINPUT31;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
         G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
         G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
         G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
         G1352gat, G1353gat, G1354gat, G1355gat;
  wire   n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054;

  XOR2_X1 U640 ( .A(G218gat), .B(n836), .Z(G1355gat) );
  NOR2_X1 U641 ( .A1(n837), .A2(n838), .ZN(n836) );
  XOR2_X1 U642 ( .A(G211gat), .B(n839), .Z(G1354gat) );
  NOR2_X1 U643 ( .A1(n840), .A2(n838), .ZN(n839) );
  XOR2_X1 U644 ( .A(G204gat), .B(n841), .Z(G1353gat) );
  NOR2_X1 U645 ( .A1(n842), .A2(n838), .ZN(n841) );
  XNOR2_X1 U646 ( .A(G197gat), .B(n843), .ZN(G1352gat) );
  NAND3_X1 U647 ( .A1(KEYINPUT6), .A2(n844), .A3(n845), .ZN(n843) );
  XOR2_X1 U648 ( .A(n846), .B(KEYINPUT24), .Z(n845) );
  INV_X1 U649 ( .A(n838), .ZN(n844) );
  NAND4_X1 U650 ( .A1(n847), .A2(n848), .A3(n849), .A4(n850), .ZN(n838) );
  NOR2_X1 U651 ( .A1(n851), .A2(n852), .ZN(n850) );
  XOR2_X1 U652 ( .A(G190gat), .B(n853), .Z(G1351gat) );
  NOR2_X1 U653 ( .A1(n837), .A2(n854), .ZN(n853) );
  XNOR2_X1 U654 ( .A(G183gat), .B(n855), .ZN(G1350gat) );
  NAND2_X1 U655 ( .A1(n856), .A2(n857), .ZN(n855) );
  XOR2_X1 U656 ( .A(n854), .B(KEYINPUT7), .Z(n856) );
  XOR2_X1 U657 ( .A(G176gat), .B(n858), .Z(G1349gat) );
  NOR2_X1 U658 ( .A1(n842), .A2(n854), .ZN(n858) );
  XOR2_X1 U659 ( .A(G169gat), .B(n859), .Z(G1348gat) );
  NOR2_X1 U660 ( .A1(n860), .A2(n854), .ZN(n859) );
  NAND4_X1 U661 ( .A1(n861), .A2(n862), .A3(n863), .A4(n848), .ZN(n854) );
  XOR2_X1 U662 ( .A(G162gat), .B(n864), .Z(G1347gat) );
  NOR2_X1 U663 ( .A1(n837), .A2(n865), .ZN(n864) );
  XOR2_X1 U664 ( .A(G155gat), .B(n866), .Z(G1346gat) );
  NOR2_X1 U665 ( .A1(n840), .A2(n865), .ZN(n866) );
  XOR2_X1 U666 ( .A(G148gat), .B(n867), .Z(G1345gat) );
  NOR2_X1 U667 ( .A1(n842), .A2(n865), .ZN(n867) );
  XOR2_X1 U668 ( .A(G141gat), .B(n868), .Z(G1344gat) );
  NOR2_X1 U669 ( .A1(n860), .A2(n865), .ZN(n868) );
  NAND4_X1 U670 ( .A1(n869), .A2(n870), .A3(n871), .A4(n848), .ZN(n865) );
  XOR2_X1 U671 ( .A(G134gat), .B(n872), .Z(G1343gat) );
  NOR2_X1 U672 ( .A1(n837), .A2(n873), .ZN(n872) );
  XOR2_X1 U673 ( .A(n874), .B(n875), .Z(G1342gat) );
  XOR2_X1 U674 ( .A(KEYINPUT27), .B(G127gat), .Z(n875) );
  NOR2_X1 U675 ( .A1(n840), .A2(n873), .ZN(n874) );
  NAND2_X1 U676 ( .A1(n876), .A2(n877), .ZN(G1341gat) );
  OR3_X1 U677 ( .A1(n842), .A2(n878), .A3(n873), .ZN(n877) );
  XOR2_X1 U678 ( .A(n879), .B(KEYINPUT4), .Z(n876) );
  NAND2_X1 U679 ( .A1(G120gat), .A2(n880), .ZN(n879) );
  XOR2_X1 U680 ( .A(KEYINPUT5), .B(n878), .Z(n880) );
  NOR3_X1 U681 ( .A1(n842), .A2(n881), .A3(n873), .ZN(n878) );
  XOR2_X1 U682 ( .A(G113gat), .B(n882), .Z(G1340gat) );
  NOR2_X1 U683 ( .A1(n860), .A2(n873), .ZN(n882) );
  NAND4_X1 U684 ( .A1(n852), .A2(n848), .A3(n851), .A4(n883), .ZN(n873) );
  NOR2_X1 U685 ( .A1(n847), .A2(n849), .ZN(n883) );
  NAND2_X1 U686 ( .A1(n884), .A2(n885), .ZN(n848) );
  NAND3_X1 U687 ( .A1(n842), .A2(n860), .A3(n886), .ZN(n885) );
  XOR2_X1 U688 ( .A(n840), .B(n837), .Z(n886) );
  NAND3_X1 U689 ( .A1(n840), .A2(n837), .A3(n887), .ZN(n884) );
  XNOR2_X1 U690 ( .A(n842), .B(n888), .ZN(n887) );
  NOR2_X1 U691 ( .A1(KEYINPUT19), .A2(n860), .ZN(n888) );
  NAND2_X1 U692 ( .A1(n889), .A2(n890), .ZN(G1339gat) );
  NAND3_X1 U693 ( .A1(n849), .A2(n891), .A3(n892), .ZN(n890) );
  NAND2_X1 U694 ( .A1(n893), .A2(G106gat), .ZN(n889) );
  XOR2_X1 U695 ( .A(n891), .B(KEYINPUT15), .Z(n893) );
  NAND3_X1 U696 ( .A1(G106gat), .A2(n849), .A3(n892), .ZN(n891) );
  INV_X1 U697 ( .A(n894), .ZN(n892) );
  XOR2_X1 U698 ( .A(G99gat), .B(n895), .Z(G1338gat) );
  NOR2_X1 U699 ( .A1(n871), .A2(n894), .ZN(n895) );
  XOR2_X1 U700 ( .A(G92gat), .B(n896), .Z(G1337gat) );
  NOR2_X1 U701 ( .A1(n869), .A2(n894), .ZN(n896) );
  XOR2_X1 U702 ( .A(G85gat), .B(n897), .Z(G1336gat) );
  NOR2_X1 U703 ( .A1(n863), .A2(n894), .ZN(n897) );
  NAND4_X1 U704 ( .A1(n898), .A2(n860), .A3(n840), .A4(n899), .ZN(n894) );
  NOR2_X1 U705 ( .A1(n837), .A2(n842), .ZN(n899) );
  XNOR2_X1 U706 ( .A(KEYINPUT31), .B(n900), .ZN(n898) );
  NAND2_X1 U707 ( .A1(n901), .A2(n902), .ZN(G1335gat) );
  NAND3_X1 U708 ( .A1(n849), .A2(n903), .A3(n904), .ZN(n902) );
  NAND2_X1 U709 ( .A1(G78gat), .A2(n905), .ZN(n901) );
  XNOR2_X1 U710 ( .A(KEYINPUT29), .B(n903), .ZN(n905) );
  NAND3_X1 U711 ( .A1(G78gat), .A2(n849), .A3(n904), .ZN(n903) );
  XNOR2_X1 U712 ( .A(G71gat), .B(n906), .ZN(G1334gat) );
  NAND2_X1 U713 ( .A1(n904), .A2(n852), .ZN(n906) );
  NAND2_X1 U714 ( .A1(n907), .A2(n908), .ZN(G1333gat) );
  NAND2_X1 U715 ( .A1(G64gat), .A2(n909), .ZN(n908) );
  XOR2_X1 U716 ( .A(KEYINPUT10), .B(n910), .Z(n907) );
  NOR2_X1 U717 ( .A1(G64gat), .A2(n909), .ZN(n910) );
  NAND2_X1 U718 ( .A1(n904), .A2(n847), .ZN(n909) );
  XOR2_X1 U719 ( .A(n911), .B(n912), .Z(G1332gat) );
  NOR2_X1 U720 ( .A1(G57gat), .A2(KEYINPUT13), .ZN(n912) );
  NAND2_X1 U721 ( .A1(n904), .A2(n851), .ZN(n911) );
  NOR3_X1 U722 ( .A1(n842), .A2(n846), .A3(n913), .ZN(n904) );
  XOR2_X1 U723 ( .A(G50gat), .B(n914), .Z(G1331gat) );
  NOR2_X1 U724 ( .A1(n861), .A2(n915), .ZN(n914) );
  XOR2_X1 U725 ( .A(G43gat), .B(n916), .Z(G1330gat) );
  NOR2_X1 U726 ( .A1(n871), .A2(n915), .ZN(n916) );
  XOR2_X1 U727 ( .A(n917), .B(n918), .Z(G1329gat) );
  NOR2_X1 U728 ( .A1(KEYINPUT12), .A2(n919), .ZN(n918) );
  NOR2_X1 U729 ( .A1(n869), .A2(n915), .ZN(n917) );
  XOR2_X1 U730 ( .A(G29gat), .B(n920), .Z(G1328gat) );
  NOR2_X1 U731 ( .A1(n863), .A2(n915), .ZN(n920) );
  NAND4_X1 U732 ( .A1(n842), .A2(n900), .A3(n840), .A4(n921), .ZN(n915) );
  NOR2_X1 U733 ( .A1(n837), .A2(n860), .ZN(n921) );
  XOR2_X1 U734 ( .A(n922), .B(G22gat), .Z(G1327gat) );
  NAND2_X1 U735 ( .A1(KEYINPUT26), .A2(n923), .ZN(n922) );
  NAND2_X1 U736 ( .A1(n924), .A2(n849), .ZN(n923) );
  XOR2_X1 U737 ( .A(n925), .B(n926), .Z(G1326gat) );
  NAND2_X1 U738 ( .A1(n924), .A2(n852), .ZN(n926) );
  XOR2_X1 U739 ( .A(n927), .B(n928), .Z(G1325gat) );
  NAND2_X1 U740 ( .A1(n924), .A2(n847), .ZN(n928) );
  XOR2_X1 U741 ( .A(n929), .B(n930), .Z(G1324gat) );
  NAND2_X1 U742 ( .A1(n924), .A2(n851), .ZN(n930) );
  NOR3_X1 U743 ( .A1(n860), .A2(n931), .A3(n913), .ZN(n924) );
  NAND3_X1 U744 ( .A1(n837), .A2(n900), .A3(n857), .ZN(n913) );
  INV_X1 U745 ( .A(n840), .ZN(n857) );
  XOR2_X1 U746 ( .A(n932), .B(n933), .Z(n840) );
  XOR2_X1 U747 ( .A(n934), .B(n935), .Z(n933) );
  XOR2_X1 U748 ( .A(n936), .B(G127gat), .Z(n935) );
  NAND3_X1 U749 ( .A1(G233gat), .A2(n937), .A3(G231gat), .ZN(n936) );
  INV_X1 U750 ( .A(KEYINPUT30), .ZN(n937) );
  XNOR2_X1 U751 ( .A(G183gat), .B(G211gat), .ZN(n934) );
  XOR2_X1 U752 ( .A(n938), .B(n939), .Z(n932) );
  XNOR2_X1 U753 ( .A(n940), .B(n941), .ZN(n938) );
  NAND2_X1 U754 ( .A1(KEYINPUT9), .A2(n942), .ZN(n940) );
  INV_X1 U755 ( .A(G155gat), .ZN(n942) );
  NAND2_X1 U756 ( .A1(n943), .A2(n944), .ZN(n900) );
  OR3_X1 U757 ( .A1(n852), .A2(n870), .A3(n847), .ZN(n944) );
  INV_X1 U758 ( .A(n869), .ZN(n847) );
  NOR2_X1 U759 ( .A1(n863), .A2(n861), .ZN(n870) );
  INV_X1 U760 ( .A(n871), .ZN(n852) );
  OR3_X1 U761 ( .A1(n851), .A2(n862), .A3(n849), .ZN(n943) );
  INV_X1 U762 ( .A(n861), .ZN(n849) );
  XOR2_X1 U763 ( .A(n945), .B(n946), .Z(n861) );
  XOR2_X1 U764 ( .A(n947), .B(n948), .Z(n946) );
  XOR2_X1 U765 ( .A(G141gat), .B(G106gat), .Z(n948) );
  XOR2_X1 U766 ( .A(G50gat), .B(G22gat), .Z(n947) );
  XOR2_X1 U767 ( .A(n949), .B(n950), .Z(n945) );
  XOR2_X1 U768 ( .A(n951), .B(n952), .Z(n950) );
  NAND2_X1 U769 ( .A1(KEYINPUT20), .A2(G78gat), .ZN(n952) );
  XOR2_X1 U770 ( .A(n953), .B(n954), .Z(n949) );
  NAND2_X1 U771 ( .A1(G228gat), .A2(G233gat), .ZN(n953) );
  NOR2_X1 U772 ( .A1(n871), .A2(n869), .ZN(n862) );
  XOR2_X1 U773 ( .A(n955), .B(n956), .Z(n869) );
  XOR2_X1 U774 ( .A(n957), .B(n958), .Z(n956) );
  XOR2_X1 U775 ( .A(G64gat), .B(n959), .Z(n958) );
  NOR2_X1 U776 ( .A1(KEYINPUT22), .A2(n919), .ZN(n959) );
  INV_X1 U777 ( .A(G36gat), .ZN(n919) );
  XOR2_X1 U778 ( .A(G92gat), .B(G8gat), .Z(n957) );
  XNOR2_X1 U779 ( .A(n960), .B(n961), .ZN(n955) );
  XOR2_X1 U780 ( .A(n962), .B(n951), .Z(n961) );
  NAND2_X1 U781 ( .A1(n963), .A2(n964), .ZN(n951) );
  NAND2_X1 U782 ( .A1(n965), .A2(n966), .ZN(n964) );
  XOR2_X1 U783 ( .A(n967), .B(n968), .Z(n966) );
  INV_X1 U784 ( .A(G204gat), .ZN(n967) );
  XOR2_X1 U785 ( .A(G218gat), .B(G211gat), .Z(n965) );
  NAND2_X1 U786 ( .A1(n969), .A2(n970), .ZN(n963) );
  XOR2_X1 U787 ( .A(n968), .B(G204gat), .Z(n970) );
  NAND2_X1 U788 ( .A1(KEYINPUT21), .A2(G197gat), .ZN(n968) );
  XNOR2_X1 U789 ( .A(G211gat), .B(G218gat), .ZN(n969) );
  NAND2_X1 U790 ( .A1(G226gat), .A2(G233gat), .ZN(n962) );
  XOR2_X1 U791 ( .A(n971), .B(n972), .Z(n871) );
  NOR2_X1 U792 ( .A1(n973), .A2(n974), .ZN(n972) );
  NOR2_X1 U793 ( .A1(n975), .A2(n976), .ZN(n974) );
  XOR2_X1 U794 ( .A(n925), .B(G43gat), .Z(n976) );
  XOR2_X1 U795 ( .A(n977), .B(G99gat), .Z(n975) );
  NOR2_X1 U796 ( .A1(n978), .A2(n979), .ZN(n973) );
  XOR2_X1 U797 ( .A(G43gat), .B(G15gat), .Z(n979) );
  XOR2_X1 U798 ( .A(n980), .B(n977), .Z(n978) );
  NAND2_X1 U799 ( .A1(KEYINPUT11), .A2(G71gat), .ZN(n977) );
  INV_X1 U800 ( .A(G99gat), .ZN(n980) );
  NAND2_X1 U801 ( .A1(n981), .A2(n982), .ZN(n971) );
  NAND2_X1 U802 ( .A1(n983), .A2(n984), .ZN(n982) );
  XOR2_X1 U803 ( .A(n985), .B(n986), .Z(n983) );
  NAND2_X1 U804 ( .A1(n987), .A2(n988), .ZN(n981) );
  XNOR2_X1 U805 ( .A(n986), .B(n985), .ZN(n988) );
  XOR2_X1 U806 ( .A(n989), .B(G113gat), .Z(n985) );
  NAND2_X1 U807 ( .A1(KEYINPUT25), .A2(n960), .ZN(n989) );
  XNOR2_X1 U808 ( .A(n990), .B(n991), .ZN(n960) );
  XOR2_X1 U809 ( .A(G190gat), .B(G183gat), .Z(n991) );
  XOR2_X1 U810 ( .A(n992), .B(G176gat), .Z(n990) );
  NAND2_X1 U811 ( .A1(KEYINPUT1), .A2(G169gat), .ZN(n992) );
  XOR2_X1 U812 ( .A(n984), .B(KEYINPUT17), .Z(n987) );
  NAND2_X1 U813 ( .A1(G233gat), .A2(n993), .ZN(n984) );
  XOR2_X1 U814 ( .A(KEYINPUT14), .B(G227gat), .Z(n993) );
  INV_X1 U815 ( .A(n863), .ZN(n851) );
  XOR2_X1 U816 ( .A(n994), .B(n995), .Z(n863) );
  XOR2_X1 U817 ( .A(n996), .B(n997), .Z(n995) );
  NAND2_X1 U818 ( .A1(n998), .A2(KEYINPUT16), .ZN(n997) );
  XOR2_X1 U819 ( .A(n999), .B(n1000), .Z(n998) );
  XOR2_X1 U820 ( .A(n1001), .B(n1002), .Z(n1000) );
  NAND2_X1 U821 ( .A1(G225gat), .A2(G233gat), .ZN(n1001) );
  XNOR2_X1 U822 ( .A(n986), .B(n954), .ZN(n999) );
  XOR2_X1 U823 ( .A(G148gat), .B(n1003), .Z(n954) );
  XOR2_X1 U824 ( .A(G162gat), .B(G155gat), .Z(n1003) );
  XNOR2_X1 U825 ( .A(n881), .B(n1004), .ZN(n986) );
  XOR2_X1 U826 ( .A(G134gat), .B(G127gat), .Z(n1004) );
  INV_X1 U827 ( .A(G120gat), .ZN(n881) );
  NAND2_X1 U828 ( .A1(n1005), .A2(n1006), .ZN(n996) );
  NAND2_X1 U829 ( .A1(G29gat), .A2(n929), .ZN(n1006) );
  XOR2_X1 U830 ( .A(n1007), .B(KEYINPUT3), .Z(n1005) );
  OR2_X1 U831 ( .A1(n929), .A2(G29gat), .ZN(n1007) );
  XNOR2_X1 U832 ( .A(G57gat), .B(G85gat), .ZN(n994) );
  XNOR2_X1 U833 ( .A(n1008), .B(n1009), .ZN(n837) );
  XOR2_X1 U834 ( .A(G162gat), .B(n1010), .Z(n1009) );
  XOR2_X1 U835 ( .A(G218gat), .B(G190gat), .Z(n1010) );
  XOR2_X1 U836 ( .A(n1011), .B(n1012), .Z(n1008) );
  XNOR2_X1 U837 ( .A(G134gat), .B(n1013), .ZN(n1012) );
  NAND3_X1 U838 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
  NAND2_X1 U839 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
  NAND2_X1 U840 ( .A1(KEYINPUT28), .A2(n1019), .ZN(n1015) );
  NAND2_X1 U841 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
  XOR2_X1 U842 ( .A(KEYINPUT8), .B(n1018), .Z(n1020) );
  INV_X1 U843 ( .A(n1022), .ZN(n1018) );
  NAND2_X1 U844 ( .A1(n1023), .A2(n1024), .ZN(n1014) );
  INV_X1 U845 ( .A(KEYINPUT28), .ZN(n1024) );
  NAND2_X1 U846 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
  NAND3_X1 U847 ( .A1(KEYINPUT8), .A2(n1021), .A3(n1022), .ZN(n1026) );
  INV_X1 U848 ( .A(n1017), .ZN(n1021) );
  OR2_X1 U849 ( .A1(n1022), .A2(KEYINPUT8), .ZN(n1025) );
  NAND2_X1 U850 ( .A1(G233gat), .A2(G232gat), .ZN(n1011) );
  INV_X1 U851 ( .A(n842), .ZN(n931) );
  XNOR2_X1 U852 ( .A(n1027), .B(n1028), .ZN(n842) );
  XOR2_X1 U853 ( .A(G148gat), .B(n1029), .Z(n1028) );
  XOR2_X1 U854 ( .A(G204gat), .B(G176gat), .Z(n1029) );
  XOR2_X1 U855 ( .A(n1030), .B(G120gat), .Z(n1027) );
  NAND2_X1 U856 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
  NAND2_X1 U857 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
  XOR2_X1 U858 ( .A(KEYINPUT2), .B(n1035), .Z(n1031) );
  NOR2_X1 U859 ( .A1(n1033), .A2(n1034), .ZN(n1035) );
  NAND2_X1 U860 ( .A1(G230gat), .A2(G233gat), .ZN(n1034) );
  XOR2_X1 U861 ( .A(n941), .B(n1022), .Z(n1033) );
  XOR2_X1 U862 ( .A(n1036), .B(n1037), .Z(n1022) );
  XOR2_X1 U863 ( .A(G99gat), .B(G92gat), .Z(n1037) );
  XNOR2_X1 U864 ( .A(G85gat), .B(G106gat), .ZN(n1036) );
  XOR2_X1 U865 ( .A(n1038), .B(n1039), .Z(n941) );
  XOR2_X1 U866 ( .A(G78gat), .B(G71gat), .Z(n1039) );
  XNOR2_X1 U867 ( .A(G57gat), .B(G64gat), .ZN(n1038) );
  INV_X1 U868 ( .A(n846), .ZN(n860) );
  XOR2_X1 U869 ( .A(n1040), .B(n1041), .Z(n846) );
  XOR2_X1 U870 ( .A(n1042), .B(n1043), .Z(n1041) );
  XNOR2_X1 U871 ( .A(G169gat), .B(G197gat), .ZN(n1043) );
  NAND2_X1 U872 ( .A1(G229gat), .A2(G233gat), .ZN(n1042) );
  XOR2_X1 U873 ( .A(n1044), .B(n1045), .Z(n1040) );
  INV_X1 U874 ( .A(n1002), .ZN(n1045) );
  XNOR2_X1 U875 ( .A(G113gat), .B(G141gat), .ZN(n1002) );
  XOR2_X1 U876 ( .A(n1017), .B(n939), .Z(n1044) );
  XNOR2_X1 U877 ( .A(n1046), .B(n1047), .ZN(n939) );
  XOR2_X1 U878 ( .A(n925), .B(n1048), .Z(n1047) );
  NAND2_X1 U879 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
  NAND2_X1 U880 ( .A1(G1gat), .A2(n927), .ZN(n1050) );
  XOR2_X1 U881 ( .A(KEYINPUT18), .B(n1051), .Z(n1049) );
  NOR2_X1 U882 ( .A1(G1gat), .A2(n927), .ZN(n1051) );
  INV_X1 U883 ( .A(G8gat), .ZN(n927) );
  INV_X1 U884 ( .A(G15gat), .ZN(n925) );
  NAND2_X1 U885 ( .A1(KEYINPUT23), .A2(G22gat), .ZN(n1046) );
  XOR2_X1 U886 ( .A(n1052), .B(n1053), .Z(n1017) );
  XOR2_X1 U887 ( .A(G36gat), .B(G29gat), .Z(n1053) );
  NAND2_X1 U888 ( .A1(KEYINPUT0), .A2(n1054), .ZN(n1052) );
  XOR2_X1 U889 ( .A(G50gat), .B(G43gat), .Z(n1054) );
  INV_X1 U890 ( .A(G1gat), .ZN(n929) );
endmodule

