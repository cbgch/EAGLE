//Key = 0011011101000101001111001000011111111101100011011001100000111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;

XOR2_X1 U748 ( .A(G107), .B(n1031), .Z(G9) );
NAND3_X1 U749 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(G75) );
NAND2_X1 U750 ( .A1(G952), .A2(n1035), .ZN(n1034) );
NAND4_X1 U751 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND4_X1 U752 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND3_X1 U757 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1050) );
NAND2_X1 U759 ( .A1(n1041), .A2(n1057), .ZN(n1046) );
INV_X1 U760 ( .A(n1058), .ZN(n1041) );
XOR2_X1 U761 ( .A(KEYINPUT23), .B(n1059), .Z(n1037) );
NOR4_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
NOR3_X1 U763 ( .A1(n1058), .A2(n1064), .A3(n1065), .ZN(n1063) );
NOR3_X1 U764 ( .A1(n1058), .A2(n1066), .A3(n1067), .ZN(n1062) );
NAND3_X1 U765 ( .A1(n1054), .A2(n1068), .A3(n1055), .ZN(n1058) );
NOR4_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1061) );
XOR2_X1 U767 ( .A(KEYINPUT15), .B(n1044), .Z(n1072) );
AND4_X1 U768 ( .A1(n1073), .A2(n1044), .A3(n1054), .A4(n1048), .ZN(n1060) );
INV_X1 U769 ( .A(n1071), .ZN(n1048) );
NAND2_X1 U770 ( .A1(n1043), .A2(n1068), .ZN(n1071) );
NAND4_X1 U771 ( .A1(n1074), .A2(n1044), .A3(n1075), .A4(n1076), .ZN(n1032) );
NOR4_X1 U772 ( .A1(n1052), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1076) );
XNOR2_X1 U773 ( .A(G478), .B(n1080), .ZN(n1079) );
NOR2_X1 U774 ( .A1(n1081), .A2(KEYINPUT26), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1078) );
XOR2_X1 U776 ( .A(KEYINPUT19), .B(G475), .Z(n1083) );
INV_X1 U777 ( .A(n1084), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1075) );
XOR2_X1 U779 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U780 ( .A(n1089), .B(n1090), .Z(n1085) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1074) );
NOR2_X1 U782 ( .A1(KEYINPUT8), .A2(n1093), .ZN(n1092) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(G72) );
XOR2_X1 U784 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U787 ( .A(G125), .B(n1102), .Z(n1101) );
NOR2_X1 U788 ( .A1(G140), .A2(KEYINPUT53), .ZN(n1102) );
XNOR2_X1 U789 ( .A(n1103), .B(n1104), .ZN(n1100) );
NOR3_X1 U790 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NOR2_X1 U791 ( .A1(G131), .A2(n1108), .ZN(n1107) );
AND3_X1 U792 ( .A1(n1108), .A2(n1109), .A3(G131), .ZN(n1106) );
INV_X1 U793 ( .A(KEYINPUT25), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1110), .A2(n1109), .ZN(n1105) );
XOR2_X1 U795 ( .A(G134), .B(G137), .Z(n1109) );
NOR2_X1 U796 ( .A1(KEYINPUT25), .A2(n1111), .ZN(n1110) );
XOR2_X1 U797 ( .A(KEYINPUT33), .B(G131), .Z(n1111) );
NAND2_X1 U798 ( .A1(n1112), .A2(n1033), .ZN(n1096) );
NAND3_X1 U799 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND2_X1 U800 ( .A1(G953), .A2(n1116), .ZN(n1094) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1116) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1033), .ZN(n1118) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U805 ( .A1(n1122), .A2(G953), .ZN(n1117) );
NAND2_X1 U806 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U807 ( .A1(n1120), .A2(n1125), .ZN(n1124) );
NAND2_X1 U808 ( .A1(G224), .A2(n1126), .ZN(n1123) );
NAND2_X1 U809 ( .A1(G898), .A2(n1120), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1120) );
NAND2_X1 U811 ( .A1(G953), .A2(n1129), .ZN(n1128) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1127) );
XOR2_X1 U813 ( .A(KEYINPUT27), .B(n1132), .Z(n1131) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U815 ( .A(KEYINPUT0), .B(n1135), .Z(n1134) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U817 ( .A(KEYINPUT10), .B(n1138), .Z(n1137) );
AND2_X1 U818 ( .A1(n1138), .A2(n1136), .ZN(n1133) );
NOR2_X1 U819 ( .A1(KEYINPUT43), .A2(n1139), .ZN(n1130) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U821 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U822 ( .A1(n1093), .A2(n1144), .ZN(n1143) );
NAND2_X1 U823 ( .A1(KEYINPUT18), .A2(n1145), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1140), .A2(n1146), .ZN(G63) );
NOR3_X1 U825 ( .A1(n1081), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR3_X1 U826 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
AND2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
NAND2_X1 U828 ( .A1(n1152), .A2(G478), .ZN(n1149) );
XNOR2_X1 U829 ( .A(n1036), .B(KEYINPUT57), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1153), .ZN(G60) );
XOR2_X1 U831 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U832 ( .A1(n1156), .A2(G475), .A3(KEYINPUT21), .ZN(n1154) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(G6) );
NOR2_X1 U834 ( .A1(KEYINPUT42), .A2(n1159), .ZN(n1158) );
INV_X1 U835 ( .A(G104), .ZN(n1159) );
NOR2_X1 U836 ( .A1(n1140), .A2(n1160), .ZN(G57) );
XOR2_X1 U837 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U838 ( .A(KEYINPUT51), .B(n1163), .Z(n1162) );
NOR2_X1 U839 ( .A1(n1087), .A2(n1144), .ZN(n1163) );
NOR2_X1 U840 ( .A1(n1140), .A2(n1164), .ZN(G54) );
XOR2_X1 U841 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U842 ( .A1(n1089), .A2(n1144), .ZN(n1166) );
INV_X1 U843 ( .A(n1156), .ZN(n1144) );
NAND3_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1165) );
OR2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND3_X1 U846 ( .A1(n1171), .A2(n1170), .A3(KEYINPUT13), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1172), .B(KEYINPUT61), .ZN(n1170) );
NOR2_X1 U848 ( .A1(KEYINPUT41), .A2(n1173), .ZN(n1171) );
NAND2_X1 U849 ( .A1(n1173), .A2(n1174), .ZN(n1167) );
INV_X1 U850 ( .A(KEYINPUT13), .ZN(n1174) );
XNOR2_X1 U851 ( .A(n1175), .B(n1176), .ZN(n1173) );
NOR2_X1 U852 ( .A1(n1140), .A2(n1177), .ZN(G51) );
XOR2_X1 U853 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U854 ( .A1(KEYINPUT14), .A2(n1180), .ZN(n1179) );
NAND2_X1 U855 ( .A1(n1156), .A2(G210), .ZN(n1178) );
NOR2_X1 U856 ( .A1(n1151), .A2(n1036), .ZN(n1156) );
AND4_X1 U857 ( .A1(n1181), .A2(n1115), .A3(n1121), .A4(n1114), .ZN(n1036) );
NAND2_X1 U858 ( .A1(n1182), .A2(n1183), .ZN(n1114) );
XNOR2_X1 U859 ( .A(n1056), .B(KEYINPUT31), .ZN(n1182) );
AND4_X1 U860 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1121) );
NOR4_X1 U861 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1157), .ZN(n1187) );
AND3_X1 U862 ( .A1(n1191), .A2(n1043), .A3(n1192), .ZN(n1157) );
NOR2_X1 U863 ( .A1(n1193), .A2(n1066), .ZN(n1190) );
XOR2_X1 U864 ( .A(n1194), .B(KEYINPUT56), .Z(n1193) );
NOR2_X1 U865 ( .A1(n1031), .A2(n1195), .ZN(n1186) );
AND3_X1 U866 ( .A1(n1056), .A2(n1043), .A3(n1191), .ZN(n1031) );
NAND3_X1 U867 ( .A1(n1196), .A2(n1197), .A3(n1054), .ZN(n1185) );
NAND2_X1 U868 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
NAND4_X1 U869 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
INV_X1 U870 ( .A(KEYINPUT40), .ZN(n1203) );
NAND2_X1 U871 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NAND2_X1 U872 ( .A1(KEYINPUT40), .A2(n1206), .ZN(n1184) );
AND4_X1 U873 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1115) );
AND3_X1 U874 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
XOR2_X1 U875 ( .A(n1113), .B(KEYINPUT17), .Z(n1181) );
NAND3_X1 U876 ( .A1(n1204), .A2(n1214), .A3(n1215), .ZN(n1113) );
XOR2_X1 U877 ( .A(n1216), .B(KEYINPUT22), .Z(n1215) );
NOR2_X1 U878 ( .A1(n1033), .A2(G952), .ZN(n1140) );
XOR2_X1 U879 ( .A(n1211), .B(n1217), .Z(G48) );
NAND2_X1 U880 ( .A1(KEYINPUT30), .A2(G146), .ZN(n1217) );
NAND2_X1 U881 ( .A1(n1183), .A2(n1192), .ZN(n1211) );
NAND2_X1 U882 ( .A1(n1218), .A2(n1219), .ZN(G45) );
NAND2_X1 U883 ( .A1(G143), .A2(n1213), .ZN(n1219) );
XOR2_X1 U884 ( .A(KEYINPUT29), .B(n1220), .Z(n1218) );
NOR2_X1 U885 ( .A1(G143), .A2(n1213), .ZN(n1220) );
NAND4_X1 U886 ( .A1(n1221), .A2(n1073), .A3(n1201), .A4(n1222), .ZN(n1213) );
NOR3_X1 U887 ( .A1(n1066), .A2(n1223), .A3(n1224), .ZN(n1222) );
XNOR2_X1 U888 ( .A(G140), .B(n1212), .ZN(G42) );
NAND2_X1 U889 ( .A1(n1214), .A2(n1225), .ZN(n1212) );
NAND2_X1 U890 ( .A1(n1226), .A2(n1227), .ZN(G39) );
OR2_X1 U891 ( .A1(n1209), .A2(G137), .ZN(n1227) );
XOR2_X1 U892 ( .A(n1228), .B(KEYINPUT49), .Z(n1226) );
NAND2_X1 U893 ( .A1(G137), .A2(n1209), .ZN(n1228) );
NAND3_X1 U894 ( .A1(n1225), .A2(n1205), .A3(n1054), .ZN(n1209) );
XNOR2_X1 U895 ( .A(G134), .B(n1207), .ZN(G36) );
NAND3_X1 U896 ( .A1(n1201), .A2(n1056), .A3(n1225), .ZN(n1207) );
XOR2_X1 U897 ( .A(n1229), .B(n1208), .Z(G33) );
NAND3_X1 U898 ( .A1(n1201), .A2(n1192), .A3(n1225), .ZN(n1208) );
NOR3_X1 U899 ( .A1(n1202), .A2(n1224), .A3(n1064), .ZN(n1225) );
INV_X1 U900 ( .A(n1044), .ZN(n1064) );
NOR2_X1 U901 ( .A1(n1230), .A2(n1040), .ZN(n1044) );
INV_X1 U902 ( .A(n1216), .ZN(n1224) );
INV_X1 U903 ( .A(n1073), .ZN(n1202) );
NAND2_X1 U904 ( .A1(n1231), .A2(n1232), .ZN(G30) );
NAND4_X1 U905 ( .A1(n1183), .A2(n1056), .A3(n1233), .A4(n1234), .ZN(n1232) );
NAND2_X1 U906 ( .A1(KEYINPUT20), .A2(G128), .ZN(n1234) );
OR2_X1 U907 ( .A1(G128), .A2(KEYINPUT62), .ZN(n1233) );
NAND3_X1 U908 ( .A1(G128), .A2(n1235), .A3(KEYINPUT20), .ZN(n1231) );
NAND3_X1 U909 ( .A1(n1183), .A2(n1056), .A3(KEYINPUT62), .ZN(n1235) );
AND4_X1 U910 ( .A1(n1073), .A2(n1236), .A3(n1205), .A4(n1216), .ZN(n1183) );
XOR2_X1 U911 ( .A(G101), .B(n1206), .Z(G3) );
AND3_X1 U912 ( .A1(n1201), .A2(n1191), .A3(n1054), .ZN(n1206) );
XOR2_X1 U913 ( .A(n1237), .B(n1238), .Z(G27) );
NAND3_X1 U914 ( .A1(n1214), .A2(n1216), .A3(n1204), .ZN(n1238) );
NAND2_X1 U915 ( .A1(n1239), .A2(n1240), .ZN(n1216) );
NAND3_X1 U916 ( .A1(G902), .A2(n1068), .A3(n1098), .ZN(n1240) );
NOR2_X1 U917 ( .A1(n1033), .A2(G900), .ZN(n1098) );
AND2_X1 U918 ( .A1(n1057), .A2(n1192), .ZN(n1214) );
XOR2_X1 U919 ( .A(G122), .B(n1241), .Z(G24) );
NOR2_X1 U920 ( .A1(n1066), .A2(n1194), .ZN(n1241) );
NAND3_X1 U921 ( .A1(n1055), .A2(n1043), .A3(n1242), .ZN(n1194) );
NOR3_X1 U922 ( .A1(n1243), .A2(n1223), .A3(n1244), .ZN(n1242) );
INV_X1 U923 ( .A(n1067), .ZN(n1043) );
NAND2_X1 U924 ( .A1(n1245), .A2(n1246), .ZN(n1067) );
INV_X1 U925 ( .A(n1070), .ZN(n1055) );
XOR2_X1 U926 ( .A(n1247), .B(n1248), .Z(G21) );
NAND4_X1 U927 ( .A1(n1204), .A2(n1054), .A3(n1249), .A4(n1205), .ZN(n1248) );
NAND2_X1 U928 ( .A1(n1250), .A2(n1251), .ZN(n1205) );
NAND2_X1 U929 ( .A1(n1057), .A2(n1252), .ZN(n1251) );
INV_X1 U930 ( .A(KEYINPUT5), .ZN(n1252) );
NAND3_X1 U931 ( .A1(n1253), .A2(n1254), .A3(KEYINPUT5), .ZN(n1250) );
NOR2_X1 U932 ( .A1(KEYINPUT38), .A2(n1244), .ZN(n1249) );
INV_X1 U933 ( .A(n1197), .ZN(n1244) );
XOR2_X1 U934 ( .A(G116), .B(n1195), .Z(G18) );
AND4_X1 U935 ( .A1(n1204), .A2(n1201), .A3(n1056), .A4(n1197), .ZN(n1195) );
NOR2_X1 U936 ( .A1(n1255), .A2(n1243), .ZN(n1056) );
INV_X1 U937 ( .A(n1065), .ZN(n1201) );
NOR2_X1 U938 ( .A1(n1070), .A2(n1066), .ZN(n1204) );
XOR2_X1 U939 ( .A(G113), .B(n1189), .Z(G15) );
AND4_X1 U940 ( .A1(n1200), .A2(n1197), .A3(n1192), .A4(n1256), .ZN(n1189) );
NOR2_X1 U941 ( .A1(n1065), .A2(n1070), .ZN(n1256) );
NAND2_X1 U942 ( .A1(n1257), .A2(n1053), .ZN(n1070) );
XNOR2_X1 U943 ( .A(n1052), .B(KEYINPUT28), .ZN(n1257) );
NAND2_X1 U944 ( .A1(n1254), .A2(n1245), .ZN(n1065) );
XNOR2_X1 U945 ( .A(n1253), .B(KEYINPUT50), .ZN(n1245) );
INV_X1 U946 ( .A(n1069), .ZN(n1192) );
NAND2_X1 U947 ( .A1(n1243), .A2(n1255), .ZN(n1069) );
INV_X1 U948 ( .A(n1221), .ZN(n1243) );
XOR2_X1 U949 ( .A(n1258), .B(n1188), .Z(G12) );
AND3_X1 U950 ( .A1(n1057), .A2(n1191), .A3(n1054), .ZN(n1188) );
NOR2_X1 U951 ( .A1(n1255), .A2(n1221), .ZN(n1054) );
XNOR2_X1 U952 ( .A(n1081), .B(n1259), .ZN(n1221) );
XOR2_X1 U953 ( .A(KEYINPUT44), .B(G478), .Z(n1259) );
AND2_X1 U954 ( .A1(n1150), .A2(n1151), .ZN(n1081) );
XNOR2_X1 U955 ( .A(n1260), .B(n1261), .ZN(n1150) );
XOR2_X1 U956 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U957 ( .A(G128), .B(G116), .Z(n1263) );
XOR2_X1 U958 ( .A(G143), .B(G134), .Z(n1262) );
XOR2_X1 U959 ( .A(n1264), .B(n1265), .Z(n1260) );
NOR2_X1 U960 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U961 ( .A(G217), .ZN(n1267) );
XNOR2_X1 U962 ( .A(G107), .B(n1268), .ZN(n1264) );
NOR2_X1 U963 ( .A1(KEYINPUT63), .A2(n1269), .ZN(n1268) );
INV_X1 U964 ( .A(G122), .ZN(n1269) );
INV_X1 U965 ( .A(n1223), .ZN(n1255) );
NOR2_X1 U966 ( .A1(n1270), .A2(n1077), .ZN(n1223) );
NOR2_X1 U967 ( .A1(n1084), .A2(G475), .ZN(n1077) );
AND2_X1 U968 ( .A1(G475), .A2(n1084), .ZN(n1270) );
NAND2_X1 U969 ( .A1(n1155), .A2(n1151), .ZN(n1084) );
XNOR2_X1 U970 ( .A(n1271), .B(n1272), .ZN(n1155) );
XOR2_X1 U971 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U972 ( .A(G122), .B(G113), .Z(n1274) );
XOR2_X1 U973 ( .A(G143), .B(G131), .Z(n1273) );
XOR2_X1 U974 ( .A(n1275), .B(n1276), .Z(n1271) );
NOR2_X1 U975 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
AND2_X1 U976 ( .A1(KEYINPUT32), .A2(n1279), .ZN(n1278) );
NOR2_X1 U977 ( .A1(KEYINPUT45), .A2(n1279), .ZN(n1277) );
XOR2_X1 U978 ( .A(n1237), .B(n1280), .Z(n1279) );
XOR2_X1 U979 ( .A(G146), .B(G140), .Z(n1280) );
INV_X1 U980 ( .A(G125), .ZN(n1237) );
XOR2_X1 U981 ( .A(n1281), .B(G104), .Z(n1275) );
NAND2_X1 U982 ( .A1(n1282), .A2(G214), .ZN(n1281) );
AND3_X1 U983 ( .A1(n1200), .A2(n1197), .A3(n1073), .ZN(n1191) );
NOR2_X1 U984 ( .A1(n1053), .A2(n1283), .ZN(n1073) );
XNOR2_X1 U985 ( .A(KEYINPUT60), .B(n1052), .ZN(n1283) );
AND2_X1 U986 ( .A1(G221), .A2(n1284), .ZN(n1052) );
XOR2_X1 U987 ( .A(n1285), .B(n1090), .Z(n1053) );
NAND2_X1 U988 ( .A1(n1286), .A2(n1151), .ZN(n1090) );
XOR2_X1 U989 ( .A(n1287), .B(n1172), .Z(n1286) );
XOR2_X1 U990 ( .A(n1288), .B(n1289), .Z(n1172) );
XOR2_X1 U991 ( .A(G140), .B(G110), .Z(n1289) );
NAND2_X1 U992 ( .A1(G227), .A2(n1033), .ZN(n1288) );
NAND4_X1 U993 ( .A1(KEYINPUT52), .A2(n1290), .A3(n1291), .A4(n1292), .ZN(n1287) );
NAND3_X1 U994 ( .A1(KEYINPUT58), .A2(n1293), .A3(n1176), .ZN(n1292) );
INV_X1 U995 ( .A(n1294), .ZN(n1293) );
OR2_X1 U996 ( .A1(n1176), .A2(KEYINPUT58), .ZN(n1291) );
NAND2_X1 U997 ( .A1(n1294), .A2(n1295), .ZN(n1290) );
NAND2_X1 U998 ( .A1(n1296), .A2(KEYINPUT58), .ZN(n1295) );
XNOR2_X1 U999 ( .A(n1176), .B(KEYINPUT34), .ZN(n1296) );
XNOR2_X1 U1000 ( .A(n1297), .B(KEYINPUT47), .ZN(n1176) );
XOR2_X1 U1001 ( .A(n1175), .B(KEYINPUT46), .Z(n1294) );
XNOR2_X1 U1002 ( .A(n1138), .B(n1103), .ZN(n1175) );
XNOR2_X1 U1003 ( .A(n1298), .B(n1299), .ZN(n1103) );
XOR2_X1 U1004 ( .A(G128), .B(n1300), .Z(n1299) );
NOR2_X1 U1005 ( .A1(KEYINPUT1), .A2(n1301), .ZN(n1300) );
NAND2_X1 U1006 ( .A1(KEYINPUT2), .A2(n1089), .ZN(n1285) );
INV_X1 U1007 ( .A(G469), .ZN(n1089) );
NAND2_X1 U1008 ( .A1(n1239), .A2(n1302), .ZN(n1197) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1068), .A4(n1129), .ZN(n1302) );
INV_X1 U1010 ( .A(G898), .ZN(n1129) );
NAND3_X1 U1011 ( .A1(n1303), .A2(n1033), .A3(G952), .ZN(n1239) );
XNOR2_X1 U1012 ( .A(KEYINPUT9), .B(n1068), .ZN(n1303) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1068) );
XOR2_X1 U1014 ( .A(n1066), .B(KEYINPUT7), .Z(n1200) );
INV_X1 U1015 ( .A(n1236), .ZN(n1066) );
NOR2_X1 U1016 ( .A1(n1042), .A2(n1040), .ZN(n1236) );
AND2_X1 U1017 ( .A1(G214), .A2(n1304), .ZN(n1040) );
NAND2_X1 U1018 ( .A1(n1151), .A2(n1305), .ZN(n1304) );
INV_X1 U1019 ( .A(n1230), .ZN(n1042) );
NAND2_X1 U1020 ( .A1(n1306), .A2(n1307), .ZN(n1230) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1308), .ZN(n1307) );
NAND2_X1 U1022 ( .A1(n1151), .A2(n1309), .ZN(n1308) );
OR2_X1 U1023 ( .A1(n1310), .A2(n1305), .ZN(n1309) );
INV_X1 U1024 ( .A(G237), .ZN(n1305) );
NAND3_X1 U1025 ( .A1(n1311), .A2(n1151), .A3(n1310), .ZN(n1306) );
XOR2_X1 U1026 ( .A(n1180), .B(KEYINPUT6), .Z(n1310) );
XNOR2_X1 U1027 ( .A(n1312), .B(n1313), .ZN(n1180) );
XNOR2_X1 U1028 ( .A(n1139), .B(n1138), .ZN(n1313) );
XOR2_X1 U1029 ( .A(G101), .B(n1314), .Z(n1138) );
XOR2_X1 U1030 ( .A(G107), .B(G104), .Z(n1314) );
XOR2_X1 U1031 ( .A(n1315), .B(n1316), .Z(n1139) );
XOR2_X1 U1032 ( .A(KEYINPUT37), .B(G110), .Z(n1316) );
NAND2_X1 U1033 ( .A1(KEYINPUT24), .A2(G122), .ZN(n1315) );
XOR2_X1 U1034 ( .A(n1317), .B(n1318), .Z(n1312) );
XOR2_X1 U1035 ( .A(G125), .B(n1319), .Z(n1318) );
NOR2_X1 U1036 ( .A1(G953), .A2(n1125), .ZN(n1319) );
INV_X1 U1037 ( .A(G224), .ZN(n1125) );
NAND2_X1 U1038 ( .A1(G210), .A2(G237), .ZN(n1311) );
AND2_X1 U1039 ( .A1(n1246), .A2(n1253), .ZN(n1057) );
XOR2_X1 U1040 ( .A(n1091), .B(n1093), .Z(n1253) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1284), .ZN(n1093) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1151), .ZN(n1284) );
NAND2_X1 U1043 ( .A1(n1145), .A2(n1151), .ZN(n1091) );
XOR2_X1 U1044 ( .A(n1320), .B(n1321), .Z(n1145) );
XOR2_X1 U1045 ( .A(n1322), .B(n1323), .Z(n1321) );
NOR2_X1 U1046 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1323) );
NOR2_X1 U1047 ( .A1(KEYINPUT4), .A2(n1324), .ZN(n1322) );
NOR2_X1 U1048 ( .A1(n1325), .A2(n1266), .ZN(n1324) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1033), .ZN(n1266) );
INV_X1 U1050 ( .A(G953), .ZN(n1033) );
INV_X1 U1051 ( .A(G221), .ZN(n1325) );
XOR2_X1 U1052 ( .A(n1326), .B(n1327), .Z(n1320) );
XOR2_X1 U1053 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1054 ( .A(G146), .B(G137), .Z(n1329) );
XOR2_X1 U1055 ( .A(KEYINPUT54), .B(KEYINPUT39), .Z(n1328) );
XOR2_X1 U1056 ( .A(n1330), .B(n1331), .Z(n1326) );
XOR2_X1 U1057 ( .A(G128), .B(G125), .Z(n1331) );
XOR2_X1 U1058 ( .A(n1247), .B(G110), .Z(n1330) );
INV_X1 U1059 ( .A(G119), .ZN(n1247) );
INV_X1 U1060 ( .A(n1254), .ZN(n1246) );
XNOR2_X1 U1061 ( .A(n1332), .B(n1088), .ZN(n1254) );
NAND2_X1 U1062 ( .A1(n1161), .A2(n1151), .ZN(n1088) );
INV_X1 U1063 ( .A(G902), .ZN(n1151) );
XOR2_X1 U1064 ( .A(n1333), .B(n1334), .Z(n1161) );
XNOR2_X1 U1065 ( .A(G101), .B(n1335), .ZN(n1334) );
NAND2_X1 U1066 ( .A1(n1282), .A2(G210), .ZN(n1335) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1282) );
XOR2_X1 U1068 ( .A(n1317), .B(n1336), .Z(n1333) );
INV_X1 U1069 ( .A(n1297), .ZN(n1336) );
XOR2_X1 U1070 ( .A(n1229), .B(n1337), .Z(n1297) );
NOR2_X1 U1071 ( .A1(KEYINPUT12), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1072 ( .A(n1339), .B(G134), .Z(n1338) );
NAND2_X1 U1073 ( .A1(KEYINPUT35), .A2(n1340), .ZN(n1339) );
INV_X1 U1074 ( .A(G137), .ZN(n1340) );
INV_X1 U1075 ( .A(G131), .ZN(n1229) );
XOR2_X1 U1076 ( .A(n1341), .B(n1136), .Z(n1317) );
XOR2_X1 U1077 ( .A(G113), .B(n1342), .Z(n1136) );
XOR2_X1 U1078 ( .A(G119), .B(G116), .Z(n1342) );
NAND2_X1 U1079 ( .A1(n1343), .A2(n1344), .ZN(n1341) );
NAND2_X1 U1080 ( .A1(n1345), .A2(G128), .ZN(n1344) );
XOR2_X1 U1081 ( .A(KEYINPUT36), .B(n1346), .Z(n1343) );
NOR2_X1 U1082 ( .A1(G128), .A2(n1345), .ZN(n1346) );
XOR2_X1 U1083 ( .A(n1347), .B(n1348), .Z(n1345) );
INV_X1 U1084 ( .A(n1298), .ZN(n1348) );
XNOR2_X1 U1085 ( .A(G143), .B(KEYINPUT55), .ZN(n1298) );
NAND2_X1 U1086 ( .A1(n1349), .A2(KEYINPUT48), .ZN(n1347) );
XOR2_X1 U1087 ( .A(n1301), .B(KEYINPUT11), .Z(n1349) );
INV_X1 U1088 ( .A(G146), .ZN(n1301) );
NAND2_X1 U1089 ( .A1(KEYINPUT59), .A2(n1087), .ZN(n1332) );
INV_X1 U1090 ( .A(G472), .ZN(n1087) );
XNOR2_X1 U1091 ( .A(G110), .B(KEYINPUT3), .ZN(n1258) );
endmodule


