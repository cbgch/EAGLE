//Key = 0000111010101010111100011010100011110011101010010000001011011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430;

XOR2_X1 U788 ( .A(n1090), .B(n1091), .Z(G9) );
NOR2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND4_X1 U790 ( .A1(KEYINPUT61), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1093) );
NOR2_X1 U791 ( .A1(KEYINPUT61), .A2(n1097), .ZN(n1092) );
NOR2_X1 U792 ( .A1(n1098), .A2(n1099), .ZN(G75) );
NOR2_X1 U793 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U794 ( .A(n1102), .ZN(n1100) );
NOR3_X1 U795 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1098) );
INV_X1 U796 ( .A(n1106), .ZN(n1105) );
NOR3_X1 U797 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR3_X1 U799 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR3_X1 U800 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1110) );
NOR4_X1 U801 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1117) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1114), .ZN(n1121) );
NOR3_X1 U803 ( .A1(n1123), .A2(n1124), .A3(n1112), .ZN(n1120) );
NAND3_X1 U804 ( .A1(n1102), .A2(n1125), .A3(n1126), .ZN(n1103) );
NAND4_X1 U805 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
NOR3_X1 U806 ( .A1(n1107), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR3_X1 U807 ( .A1(n1116), .A2(n1133), .A3(n1134), .ZN(n1132) );
NOR2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
NAND4_X1 U809 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1102) );
NOR4_X1 U810 ( .A1(n1116), .A2(n1141), .A3(n1109), .A4(n1142), .ZN(n1140) );
INV_X1 U811 ( .A(n1123), .ZN(n1141) );
INV_X1 U812 ( .A(n1136), .ZN(n1116) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1139) );
NAND2_X1 U814 ( .A1(n1145), .A2(KEYINPUT34), .ZN(n1143) );
XOR2_X1 U815 ( .A(n1146), .B(KEYINPUT12), .Z(n1145) );
XOR2_X1 U816 ( .A(n1147), .B(G469), .Z(n1138) );
XOR2_X1 U817 ( .A(n1148), .B(n1149), .Z(n1137) );
NOR2_X1 U818 ( .A1(KEYINPUT13), .A2(n1150), .ZN(n1149) );
INV_X1 U819 ( .A(G478), .ZN(n1150) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(G72) );
NOR2_X1 U821 ( .A1(n1153), .A2(n1125), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
NAND2_X1 U824 ( .A1(n1158), .A2(n1125), .ZN(n1157) );
XOR2_X1 U825 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND3_X1 U826 ( .A1(G900), .A2(n1160), .A3(G953), .ZN(n1156) );
XNOR2_X1 U827 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U828 ( .A(G131), .B(n1163), .Z(n1162) );
XOR2_X1 U829 ( .A(KEYINPUT50), .B(G134), .Z(n1163) );
XOR2_X1 U830 ( .A(n1164), .B(n1165), .Z(n1161) );
XOR2_X1 U831 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U832 ( .A(n1168), .B(n1169), .Z(G69) );
XOR2_X1 U833 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U834 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U835 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U836 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U837 ( .A1(KEYINPUT47), .A2(n1178), .ZN(n1176) );
XOR2_X1 U838 ( .A(KEYINPUT32), .B(n1179), .Z(n1174) );
NOR2_X1 U839 ( .A1(G898), .A2(n1125), .ZN(n1172) );
NOR2_X1 U840 ( .A1(G953), .A2(n1180), .ZN(n1170) );
NOR2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U842 ( .A(n1097), .B(KEYINPUT33), .Z(n1181) );
NOR2_X1 U843 ( .A1(n1183), .A2(n1125), .ZN(n1168) );
AND2_X1 U844 ( .A1(G224), .A2(G898), .ZN(n1183) );
NOR2_X1 U845 ( .A1(n1184), .A2(n1185), .ZN(G66) );
XOR2_X1 U846 ( .A(n1186), .B(n1187), .Z(n1185) );
NAND3_X1 U847 ( .A1(n1188), .A2(G217), .A3(KEYINPUT54), .ZN(n1186) );
NOR2_X1 U848 ( .A1(n1184), .A2(n1189), .ZN(G63) );
XOR2_X1 U849 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U850 ( .A1(n1188), .A2(G478), .ZN(n1190) );
NOR2_X1 U851 ( .A1(n1184), .A2(n1192), .ZN(G60) );
NOR3_X1 U852 ( .A1(n1193), .A2(n1144), .A3(n1194), .ZN(n1192) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NOR2_X1 U854 ( .A1(n1106), .A2(n1146), .ZN(n1195) );
INV_X1 U855 ( .A(G475), .ZN(n1146) );
XOR2_X1 U856 ( .A(n1197), .B(KEYINPUT16), .Z(n1193) );
NAND3_X1 U857 ( .A1(n1188), .A2(G475), .A3(n1196), .ZN(n1197) );
XOR2_X1 U858 ( .A(n1198), .B(n1199), .Z(G6) );
XOR2_X1 U859 ( .A(KEYINPUT21), .B(G104), .Z(n1199) );
NOR2_X1 U860 ( .A1(n1113), .A2(n1200), .ZN(n1198) );
NOR3_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(G57) );
NOR2_X1 U862 ( .A1(n1101), .A2(n1204), .ZN(n1203) );
AND2_X1 U863 ( .A1(n1204), .A2(n1184), .ZN(n1202) );
INV_X1 U864 ( .A(KEYINPUT22), .ZN(n1204) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(n1201) );
XOR2_X1 U866 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U867 ( .A(n1209), .B(n1210), .ZN(n1208) );
NAND2_X1 U868 ( .A1(KEYINPUT18), .A2(n1211), .ZN(n1209) );
XOR2_X1 U869 ( .A(n1212), .B(n1213), .Z(n1205) );
XOR2_X1 U870 ( .A(G101), .B(n1214), .Z(n1213) );
NOR2_X1 U871 ( .A1(KEYINPUT46), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U872 ( .A(n1216), .B(KEYINPUT56), .ZN(n1215) );
NAND2_X1 U873 ( .A1(n1188), .A2(G472), .ZN(n1212) );
NOR2_X1 U874 ( .A1(n1184), .A2(n1217), .ZN(G54) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1217) );
XNOR2_X1 U876 ( .A(n1210), .B(n1220), .ZN(n1219) );
XOR2_X1 U877 ( .A(n1221), .B(n1222), .Z(n1220) );
AND2_X1 U878 ( .A1(G469), .A2(n1188), .ZN(n1222) );
NOR3_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1221) );
AND2_X1 U880 ( .A1(n1226), .A2(KEYINPUT30), .ZN(n1225) );
NOR3_X1 U881 ( .A1(KEYINPUT30), .A2(n1226), .A3(n1227), .ZN(n1224) );
XOR2_X1 U882 ( .A(n1164), .B(n1228), .Z(n1218) );
NOR3_X1 U883 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(G51) );
AND2_X1 U884 ( .A1(n1184), .A2(KEYINPUT4), .ZN(n1231) );
NOR2_X1 U885 ( .A1(n1125), .A2(G952), .ZN(n1184) );
NOR2_X1 U886 ( .A1(KEYINPUT4), .A2(n1101), .ZN(n1230) );
OR2_X1 U887 ( .A1(G952), .A2(G953), .ZN(n1101) );
XOR2_X1 U888 ( .A(n1232), .B(n1233), .Z(n1229) );
NOR2_X1 U889 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NOR2_X1 U890 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NOR2_X1 U891 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
AND2_X1 U892 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR3_X1 U893 ( .A1(n1241), .A2(n1242), .A3(n1240), .ZN(n1238) );
NOR2_X1 U894 ( .A1(n1243), .A2(n1244), .ZN(n1234) );
NOR2_X1 U895 ( .A1(n1242), .A2(n1245), .ZN(n1244) );
XOR2_X1 U896 ( .A(n1241), .B(n1240), .Z(n1245) );
INV_X1 U897 ( .A(KEYINPUT59), .ZN(n1240) );
INV_X1 U898 ( .A(n1237), .ZN(n1243) );
XOR2_X1 U899 ( .A(n1246), .B(n1247), .Z(n1232) );
NOR2_X1 U900 ( .A1(KEYINPUT27), .A2(n1248), .ZN(n1247) );
NAND2_X1 U901 ( .A1(n1188), .A2(n1249), .ZN(n1246) );
NOR2_X1 U902 ( .A1(n1250), .A2(n1106), .ZN(n1188) );
NOR3_X1 U903 ( .A1(n1182), .A2(n1251), .A3(n1159), .ZN(n1106) );
NAND4_X1 U904 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1159) );
NOR3_X1 U905 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1255) );
INV_X1 U906 ( .A(n1259), .ZN(n1257) );
NAND2_X1 U907 ( .A1(n1094), .A2(n1260), .ZN(n1254) );
NAND3_X1 U908 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
XOR2_X1 U909 ( .A(n1264), .B(KEYINPUT31), .Z(n1263) );
NAND3_X1 U910 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1262) );
NAND2_X1 U911 ( .A1(n1268), .A2(n1269), .ZN(n1265) );
NAND3_X1 U912 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1269) );
INV_X1 U913 ( .A(KEYINPUT41), .ZN(n1271) );
NAND2_X1 U914 ( .A1(n1273), .A2(n1133), .ZN(n1268) );
NAND2_X1 U915 ( .A1(KEYINPUT41), .A2(n1274), .ZN(n1261) );
NAND2_X1 U916 ( .A1(n1275), .A2(n1272), .ZN(n1274) );
INV_X1 U917 ( .A(n1097), .ZN(n1251) );
NAND2_X1 U918 ( .A1(n1276), .A2(n1095), .ZN(n1097) );
NOR3_X1 U919 ( .A1(n1122), .A2(n1109), .A3(n1277), .ZN(n1095) );
INV_X1 U920 ( .A(n1272), .ZN(n1122) );
NAND4_X1 U921 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1182) );
NOR3_X1 U922 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1281) );
NOR2_X1 U923 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NOR3_X1 U924 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1285) );
NOR4_X1 U925 ( .A1(KEYINPUT44), .A2(n1267), .A3(n1290), .A4(n1112), .ZN(n1289) );
NOR3_X1 U926 ( .A1(n1291), .A2(n1109), .A3(n1114), .ZN(n1288) );
INV_X1 U927 ( .A(n1135), .ZN(n1109) );
AND2_X1 U928 ( .A1(n1119), .A2(n1133), .ZN(n1287) );
NOR2_X1 U929 ( .A1(n1113), .A2(n1292), .ZN(n1283) );
XNOR2_X1 U930 ( .A(KEYINPUT23), .B(n1200), .ZN(n1292) );
NAND4_X1 U931 ( .A1(n1293), .A2(n1267), .A3(n1135), .A4(n1294), .ZN(n1200) );
NOR2_X1 U932 ( .A1(n1295), .A2(n1296), .ZN(n1282) );
INV_X1 U933 ( .A(KEYINPUT44), .ZN(n1296) );
NAND4_X1 U934 ( .A1(n1118), .A2(n1133), .A3(n1297), .A4(n1298), .ZN(n1280) );
OR2_X1 U935 ( .A1(n1276), .A2(KEYINPUT36), .ZN(n1298) );
NAND2_X1 U936 ( .A1(KEYINPUT36), .A2(n1299), .ZN(n1297) );
NAND2_X1 U937 ( .A1(n1094), .A2(n1096), .ZN(n1299) );
INV_X1 U938 ( .A(n1294), .ZN(n1096) );
XOR2_X1 U939 ( .A(n1300), .B(n1301), .Z(G48) );
NOR2_X1 U940 ( .A1(KEYINPUT3), .A2(n1302), .ZN(n1301) );
NOR2_X1 U941 ( .A1(n1113), .A2(n1264), .ZN(n1300) );
NAND2_X1 U942 ( .A1(n1275), .A2(n1293), .ZN(n1264) );
AND3_X1 U943 ( .A1(n1270), .A2(n1266), .A3(n1267), .ZN(n1275) );
NAND2_X1 U944 ( .A1(n1303), .A2(n1304), .ZN(G45) );
NAND2_X1 U945 ( .A1(G143), .A2(n1305), .ZN(n1304) );
XOR2_X1 U946 ( .A(n1306), .B(KEYINPUT43), .Z(n1303) );
OR2_X1 U947 ( .A1(n1305), .A2(G143), .ZN(n1306) );
NAND3_X1 U948 ( .A1(n1273), .A2(n1133), .A3(n1307), .ZN(n1305) );
NOR3_X1 U949 ( .A1(n1113), .A2(n1308), .A3(n1277), .ZN(n1307) );
XOR2_X1 U950 ( .A(n1266), .B(KEYINPUT35), .Z(n1308) );
XNOR2_X1 U951 ( .A(G140), .B(n1252), .ZN(G42) );
NAND3_X1 U952 ( .A1(n1134), .A2(n1293), .A3(n1309), .ZN(n1252) );
XOR2_X1 U953 ( .A(n1253), .B(n1310), .Z(G39) );
NAND2_X1 U954 ( .A1(KEYINPUT17), .A2(G137), .ZN(n1310) );
NAND3_X1 U955 ( .A1(n1309), .A2(n1270), .A3(n1129), .ZN(n1253) );
XOR2_X1 U956 ( .A(G134), .B(n1256), .Z(G36) );
AND3_X1 U957 ( .A1(n1309), .A2(n1272), .A3(n1133), .ZN(n1256) );
XOR2_X1 U958 ( .A(n1258), .B(n1311), .Z(G33) );
NOR2_X1 U959 ( .A1(KEYINPUT0), .A2(n1312), .ZN(n1311) );
INV_X1 U960 ( .A(G131), .ZN(n1312) );
AND3_X1 U961 ( .A1(n1309), .A2(n1293), .A3(n1133), .ZN(n1258) );
AND4_X1 U962 ( .A1(n1267), .A2(n1128), .A3(n1266), .A4(n1136), .ZN(n1309) );
INV_X1 U963 ( .A(n1115), .ZN(n1128) );
XOR2_X1 U964 ( .A(n1313), .B(KEYINPUT57), .Z(n1115) );
XOR2_X1 U965 ( .A(G128), .B(n1314), .Z(G30) );
NOR3_X1 U966 ( .A1(n1315), .A2(n1113), .A3(n1316), .ZN(n1314) );
XOR2_X1 U967 ( .A(KEYINPUT5), .B(n1267), .Z(n1316) );
INV_X1 U968 ( .A(n1277), .ZN(n1267) );
NAND3_X1 U969 ( .A1(n1270), .A2(n1266), .A3(n1272), .ZN(n1315) );
NAND2_X1 U970 ( .A1(n1317), .A2(n1318), .ZN(G3) );
OR2_X1 U971 ( .A1(n1319), .A2(G101), .ZN(n1318) );
XOR2_X1 U972 ( .A(n1320), .B(KEYINPUT53), .Z(n1317) );
NAND2_X1 U973 ( .A1(G101), .A2(n1319), .ZN(n1320) );
NAND3_X1 U974 ( .A1(n1133), .A2(n1276), .A3(n1118), .ZN(n1319) );
XOR2_X1 U975 ( .A(n1321), .B(n1259), .Z(G27) );
NAND4_X1 U976 ( .A1(n1119), .A2(n1134), .A3(n1094), .A4(n1266), .ZN(n1259) );
NAND2_X1 U977 ( .A1(n1107), .A2(n1322), .ZN(n1266) );
NAND4_X1 U978 ( .A1(G953), .A2(G902), .A3(n1323), .A4(n1155), .ZN(n1322) );
INV_X1 U979 ( .A(G900), .ZN(n1155) );
AND2_X1 U980 ( .A1(n1127), .A2(n1293), .ZN(n1119) );
XNOR2_X1 U981 ( .A(G122), .B(n1324), .ZN(G24) );
NAND4_X1 U982 ( .A1(n1273), .A2(n1276), .A3(n1135), .A4(n1325), .ZN(n1324) );
XOR2_X1 U983 ( .A(KEYINPUT2), .B(n1127), .Z(n1325) );
INV_X1 U984 ( .A(n1114), .ZN(n1127) );
NOR2_X1 U985 ( .A1(n1326), .A2(n1327), .ZN(n1135) );
INV_X1 U986 ( .A(n1291), .ZN(n1273) );
NAND2_X1 U987 ( .A1(n1328), .A2(n1329), .ZN(n1291) );
XNOR2_X1 U988 ( .A(G119), .B(n1278), .ZN(G21) );
NAND3_X1 U989 ( .A1(n1129), .A2(n1270), .A3(n1330), .ZN(n1278) );
NAND2_X1 U990 ( .A1(n1331), .A2(n1332), .ZN(n1270) );
NAND3_X1 U991 ( .A1(n1327), .A2(n1326), .A3(n1333), .ZN(n1332) );
INV_X1 U992 ( .A(KEYINPUT11), .ZN(n1333) );
INV_X1 U993 ( .A(n1334), .ZN(n1327) );
NAND2_X1 U994 ( .A1(KEYINPUT11), .A2(n1133), .ZN(n1331) );
XOR2_X1 U995 ( .A(n1335), .B(n1279), .Z(G18) );
NAND3_X1 U996 ( .A1(n1133), .A2(n1272), .A3(n1330), .ZN(n1279) );
NOR2_X1 U997 ( .A1(n1329), .A2(n1336), .ZN(n1272) );
XNOR2_X1 U998 ( .A(G113), .B(n1337), .ZN(G15) );
NAND4_X1 U999 ( .A1(KEYINPUT63), .A2(n1330), .A3(n1133), .A4(n1293), .ZN(n1337) );
AND2_X1 U1000 ( .A1(n1336), .A2(n1329), .ZN(n1293) );
NOR2_X1 U1001 ( .A1(n1326), .A2(n1334), .ZN(n1133) );
NOR2_X1 U1002 ( .A1(n1114), .A2(n1286), .ZN(n1330) );
NAND2_X1 U1003 ( .A1(n1123), .A2(n1338), .ZN(n1114) );
XOR2_X1 U1004 ( .A(n1339), .B(n1295), .Z(G12) );
NAND3_X1 U1005 ( .A1(n1134), .A2(n1276), .A3(n1118), .ZN(n1295) );
NOR2_X1 U1006 ( .A1(n1112), .A2(n1277), .ZN(n1118) );
NAND2_X1 U1007 ( .A1(n1124), .A2(n1123), .ZN(n1277) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1340), .ZN(n1123) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1250), .ZN(n1340) );
INV_X1 U1010 ( .A(n1338), .ZN(n1124) );
NAND3_X1 U1011 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1338) );
NAND2_X1 U1012 ( .A1(G469), .A2(n1344), .ZN(n1343) );
OR3_X1 U1013 ( .A1(n1344), .A2(G469), .A3(KEYINPUT1), .ZN(n1342) );
NAND2_X1 U1014 ( .A1(KEYINPUT39), .A2(n1147), .ZN(n1344) );
NAND2_X1 U1015 ( .A1(n1345), .A2(KEYINPUT1), .ZN(n1341) );
INV_X1 U1016 ( .A(n1147), .ZN(n1345) );
NAND2_X1 U1017 ( .A1(n1346), .A2(n1250), .ZN(n1147) );
XOR2_X1 U1018 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1019 ( .A(n1164), .B(n1210), .ZN(n1348) );
XOR2_X1 U1020 ( .A(n1349), .B(G128), .Z(n1164) );
NAND2_X1 U1021 ( .A1(KEYINPUT60), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1022 ( .A(G143), .B(n1351), .Z(n1350) );
NOR2_X1 U1023 ( .A1(KEYINPUT45), .A2(n1302), .ZN(n1351) );
XOR2_X1 U1024 ( .A(n1352), .B(n1353), .Z(n1347) );
NOR2_X1 U1025 ( .A1(n1354), .A2(n1223), .ZN(n1353) );
AND2_X1 U1026 ( .A1(n1226), .A2(n1227), .ZN(n1223) );
NOR2_X1 U1027 ( .A1(n1226), .A2(n1227), .ZN(n1354) );
XOR2_X1 U1028 ( .A(n1339), .B(G140), .Z(n1227) );
NOR2_X1 U1029 ( .A1(n1154), .A2(G953), .ZN(n1226) );
INV_X1 U1030 ( .A(G227), .ZN(n1154) );
NAND2_X1 U1031 ( .A1(KEYINPUT8), .A2(n1228), .ZN(n1352) );
INV_X1 U1032 ( .A(n1177), .ZN(n1228) );
INV_X1 U1033 ( .A(n1129), .ZN(n1112) );
NOR2_X1 U1034 ( .A1(n1328), .A2(n1329), .ZN(n1129) );
XOR2_X1 U1035 ( .A(n1144), .B(G475), .Z(n1329) );
NOR2_X1 U1036 ( .A1(n1196), .A2(G902), .ZN(n1144) );
XOR2_X1 U1037 ( .A(n1355), .B(n1356), .Z(n1196) );
XOR2_X1 U1038 ( .A(n1357), .B(n1358), .Z(n1356) );
XNOR2_X1 U1039 ( .A(n1359), .B(n1360), .ZN(n1358) );
NOR2_X1 U1040 ( .A1(G131), .A2(KEYINPUT15), .ZN(n1360) );
NOR2_X1 U1041 ( .A1(KEYINPUT25), .A2(n1361), .ZN(n1359) );
XNOR2_X1 U1042 ( .A(n1167), .B(n1362), .ZN(n1361) );
NOR2_X1 U1043 ( .A1(KEYINPUT37), .A2(n1302), .ZN(n1362) );
INV_X1 U1044 ( .A(G146), .ZN(n1302) );
XOR2_X1 U1045 ( .A(G140), .B(G125), .Z(n1167) );
NAND3_X1 U1046 ( .A1(n1363), .A2(n1125), .A3(G214), .ZN(n1357) );
XOR2_X1 U1047 ( .A(n1364), .B(n1365), .Z(n1355) );
XNOR2_X1 U1048 ( .A(n1366), .B(n1367), .ZN(n1364) );
INV_X1 U1049 ( .A(n1336), .ZN(n1328) );
XOR2_X1 U1050 ( .A(n1148), .B(G478), .Z(n1336) );
NAND2_X1 U1051 ( .A1(n1191), .A2(n1250), .ZN(n1148) );
XOR2_X1 U1052 ( .A(n1368), .B(n1369), .Z(n1191) );
XOR2_X1 U1053 ( .A(G116), .B(n1370), .Z(n1369) );
XOR2_X1 U1054 ( .A(G134), .B(G128), .Z(n1370) );
XOR2_X1 U1055 ( .A(n1371), .B(n1366), .Z(n1368) );
XOR2_X1 U1056 ( .A(G143), .B(n1372), .Z(n1366) );
XOR2_X1 U1057 ( .A(n1373), .B(G107), .Z(n1371) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1374), .ZN(n1373) );
INV_X1 U1059 ( .A(n1286), .ZN(n1276) );
NAND2_X1 U1060 ( .A1(n1094), .A2(n1294), .ZN(n1286) );
NAND2_X1 U1061 ( .A1(n1107), .A2(n1375), .ZN(n1294) );
NAND4_X1 U1062 ( .A1(G953), .A2(G902), .A3(n1323), .A4(n1376), .ZN(n1375) );
INV_X1 U1063 ( .A(G898), .ZN(n1376) );
NAND3_X1 U1064 ( .A1(n1323), .A2(n1125), .A3(G952), .ZN(n1107) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1323) );
INV_X1 U1066 ( .A(n1113), .ZN(n1094) );
NAND2_X1 U1067 ( .A1(n1142), .A2(n1136), .ZN(n1113) );
NAND2_X1 U1068 ( .A1(G214), .A2(n1377), .ZN(n1136) );
INV_X1 U1069 ( .A(n1313), .ZN(n1142) );
XOR2_X1 U1070 ( .A(n1378), .B(n1249), .Z(n1313) );
AND2_X1 U1071 ( .A1(G210), .A2(n1377), .ZN(n1249) );
NAND2_X1 U1072 ( .A1(n1363), .A2(n1250), .ZN(n1377) );
NAND2_X1 U1073 ( .A1(n1379), .A2(n1250), .ZN(n1378) );
XOR2_X1 U1074 ( .A(n1380), .B(n1381), .Z(n1379) );
XOR2_X1 U1075 ( .A(n1237), .B(n1248), .Z(n1381) );
XNOR2_X1 U1076 ( .A(n1382), .B(n1178), .ZN(n1248) );
XOR2_X1 U1077 ( .A(n1383), .B(n1372), .Z(n1178) );
XOR2_X1 U1078 ( .A(G122), .B(KEYINPUT14), .Z(n1372) );
NAND2_X1 U1079 ( .A1(KEYINPUT26), .A2(n1339), .ZN(n1383) );
XOR2_X1 U1080 ( .A(n1384), .B(n1179), .Z(n1382) );
AND2_X1 U1081 ( .A1(n1385), .A2(n1386), .ZN(n1179) );
NAND2_X1 U1082 ( .A1(n1367), .A2(n1387), .ZN(n1386) );
OR2_X1 U1083 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
XOR2_X1 U1084 ( .A(KEYINPUT40), .B(n1390), .Z(n1385) );
NOR3_X1 U1085 ( .A1(n1391), .A2(n1389), .A3(n1388), .ZN(n1390) );
NOR2_X1 U1086 ( .A1(n1392), .A2(G119), .ZN(n1389) );
XOR2_X1 U1087 ( .A(G116), .B(n1393), .Z(n1392) );
XNOR2_X1 U1088 ( .A(KEYINPUT58), .B(KEYINPUT49), .ZN(n1393) );
XNOR2_X1 U1089 ( .A(n1367), .B(KEYINPUT6), .ZN(n1391) );
NAND2_X1 U1090 ( .A1(KEYINPUT28), .A2(n1177), .ZN(n1384) );
XOR2_X1 U1091 ( .A(n1394), .B(n1365), .Z(n1177) );
XOR2_X1 U1092 ( .A(G104), .B(KEYINPUT55), .Z(n1365) );
XOR2_X1 U1093 ( .A(n1090), .B(G101), .Z(n1394) );
INV_X1 U1094 ( .A(G107), .ZN(n1090) );
NAND2_X1 U1095 ( .A1(G224), .A2(n1125), .ZN(n1237) );
XOR2_X1 U1096 ( .A(n1395), .B(n1396), .Z(n1380) );
XOR2_X1 U1097 ( .A(KEYINPUT42), .B(KEYINPUT29), .Z(n1396) );
NOR2_X1 U1098 ( .A1(KEYINPUT9), .A2(n1397), .ZN(n1395) );
NOR2_X1 U1099 ( .A1(n1242), .A2(n1241), .ZN(n1397) );
AND2_X1 U1100 ( .A1(n1216), .A2(n1321), .ZN(n1241) );
NOR2_X1 U1101 ( .A1(n1321), .A2(n1216), .ZN(n1242) );
INV_X1 U1102 ( .A(n1290), .ZN(n1134) );
NAND2_X1 U1103 ( .A1(n1334), .A2(n1326), .ZN(n1290) );
NAND3_X1 U1104 ( .A1(n1398), .A2(n1399), .A3(n1400), .ZN(n1326) );
OR2_X1 U1105 ( .A1(n1401), .A2(n1187), .ZN(n1400) );
NAND3_X1 U1106 ( .A1(n1187), .A2(n1401), .A3(n1250), .ZN(n1399) );
NAND2_X1 U1107 ( .A1(G217), .A2(n1402), .ZN(n1401) );
XOR2_X1 U1108 ( .A(n1403), .B(n1404), .Z(n1187) );
XNOR2_X1 U1109 ( .A(n1405), .B(n1406), .ZN(n1404) );
XOR2_X1 U1110 ( .A(n1407), .B(n1408), .Z(n1406) );
NOR2_X1 U1111 ( .A1(n1409), .A2(n1410), .ZN(n1408) );
XOR2_X1 U1112 ( .A(n1411), .B(KEYINPUT38), .Z(n1410) );
NAND2_X1 U1113 ( .A1(n1166), .A2(n1412), .ZN(n1411) );
NAND2_X1 U1114 ( .A1(n1374), .A2(G221), .ZN(n1412) );
INV_X1 U1115 ( .A(n1413), .ZN(n1166) );
AND3_X1 U1116 ( .A1(n1413), .A2(G221), .A3(n1374), .ZN(n1409) );
NOR2_X1 U1117 ( .A1(n1402), .A2(G953), .ZN(n1374) );
INV_X1 U1118 ( .A(G234), .ZN(n1402) );
NAND2_X1 U1119 ( .A1(n1414), .A2(n1415), .ZN(n1407) );
NAND2_X1 U1120 ( .A1(G140), .A2(n1321), .ZN(n1415) );
XOR2_X1 U1121 ( .A(n1416), .B(KEYINPUT48), .Z(n1414) );
OR2_X1 U1122 ( .A1(n1321), .A2(G140), .ZN(n1416) );
INV_X1 U1123 ( .A(G125), .ZN(n1321) );
XOR2_X1 U1124 ( .A(n1339), .B(n1417), .Z(n1403) );
XOR2_X1 U1125 ( .A(KEYINPUT7), .B(G119), .Z(n1417) );
NAND2_X1 U1126 ( .A1(G217), .A2(G902), .ZN(n1398) );
XOR2_X1 U1127 ( .A(n1418), .B(G472), .Z(n1334) );
NAND2_X1 U1128 ( .A1(n1419), .A2(n1250), .ZN(n1418) );
INV_X1 U1129 ( .A(G902), .ZN(n1250) );
XOR2_X1 U1130 ( .A(n1420), .B(n1421), .Z(n1419) );
XNOR2_X1 U1131 ( .A(n1422), .B(n1216), .ZN(n1421) );
XOR2_X1 U1132 ( .A(G143), .B(n1405), .Z(n1216) );
XOR2_X1 U1133 ( .A(G128), .B(G146), .Z(n1405) );
NAND2_X1 U1134 ( .A1(KEYINPUT24), .A2(n1207), .ZN(n1422) );
XNOR2_X1 U1135 ( .A(n1367), .B(n1423), .ZN(n1207) );
NOR2_X1 U1136 ( .A1(KEYINPUT20), .A2(n1424), .ZN(n1423) );
NOR2_X1 U1137 ( .A1(n1425), .A2(n1388), .ZN(n1424) );
AND2_X1 U1138 ( .A1(G119), .A2(n1335), .ZN(n1388) );
NOR2_X1 U1139 ( .A1(G119), .A2(n1335), .ZN(n1425) );
INV_X1 U1140 ( .A(G116), .ZN(n1335) );
XOR2_X1 U1141 ( .A(G113), .B(KEYINPUT51), .Z(n1367) );
XOR2_X1 U1142 ( .A(n1426), .B(n1427), .Z(n1420) );
XOR2_X1 U1143 ( .A(G101), .B(n1211), .Z(n1427) );
AND3_X1 U1144 ( .A1(n1363), .A2(n1125), .A3(G210), .ZN(n1211) );
INV_X1 U1145 ( .A(G953), .ZN(n1125) );
INV_X1 U1146 ( .A(G237), .ZN(n1363) );
NAND2_X1 U1147 ( .A1(KEYINPUT19), .A2(n1210), .ZN(n1426) );
XOR2_X1 U1148 ( .A(n1428), .B(n1429), .Z(n1210) );
NOR2_X1 U1149 ( .A1(KEYINPUT52), .A2(n1413), .ZN(n1429) );
XNOR2_X1 U1150 ( .A(G137), .B(KEYINPUT10), .ZN(n1413) );
XOR2_X1 U1151 ( .A(n1430), .B(G134), .Z(n1428) );
NAND2_X1 U1152 ( .A1(KEYINPUT62), .A2(G131), .ZN(n1430) );
INV_X1 U1153 ( .A(G110), .ZN(n1339) );
endmodule


