//Key = 1111010010111001100011101110010100100001111101011000110000110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389;

XOR2_X1 U762 ( .A(G107), .B(n1059), .Z(G9) );
NOR3_X1 U763 ( .A1(n1060), .A2(KEYINPUT54), .A3(n1061), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(G75) );
XOR2_X1 U765 ( .A(KEYINPUT13), .B(n1064), .Z(n1063) );
NOR3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1065) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1073) );
NAND3_X1 U772 ( .A1(n1078), .A2(n1080), .A3(n1071), .ZN(n1069) );
AND3_X1 U773 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1071) );
NAND3_X1 U774 ( .A1(n1083), .A2(n1084), .A3(n1076), .ZN(n1068) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1087), .A2(n1082), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1078), .A2(n1088), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1091), .ZN(n1090) );
NAND2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1082), .A2(n1094), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
INV_X1 U784 ( .A(n1099), .ZN(n1083) );
NOR2_X1 U785 ( .A1(G952), .A2(n1066), .ZN(n1062) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1066) );
NAND4_X1 U787 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
NOR4_X1 U788 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
XOR2_X1 U789 ( .A(KEYINPUT60), .B(n1110), .Z(n1109) );
XOR2_X1 U790 ( .A(n1111), .B(n1112), .Z(n1106) );
NOR3_X1 U791 ( .A1(n1113), .A2(n1097), .A3(n1077), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1114), .A2(n1115), .ZN(n1103) );
XOR2_X1 U793 ( .A(n1116), .B(n1117), .Z(n1102) );
NOR2_X1 U794 ( .A1(G475), .A2(KEYINPUT7), .ZN(n1117) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(G72) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1100), .ZN(n1119) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND3_X1 U798 ( .A1(KEYINPUT47), .A2(n1123), .A3(n1124), .ZN(n1118) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U800 ( .A1(n1127), .A2(G953), .ZN(n1126) );
OR2_X1 U801 ( .A1(n1128), .A2(KEYINPUT17), .ZN(n1125) );
NAND2_X1 U802 ( .A1(KEYINPUT17), .A2(n1128), .ZN(n1123) );
NAND2_X1 U803 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U804 ( .A1(G953), .A2(n1122), .ZN(n1130) );
XOR2_X1 U805 ( .A(n1131), .B(n1132), .Z(n1129) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U807 ( .A(n1135), .B(KEYINPUT61), .Z(n1134) );
NAND3_X1 U808 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1133) );
NAND2_X1 U809 ( .A1(KEYINPUT30), .A2(G125), .ZN(n1138) );
OR3_X1 U810 ( .A1(G125), .A2(KEYINPUT30), .A3(n1139), .ZN(n1137) );
NAND2_X1 U811 ( .A1(n1140), .A2(n1139), .ZN(n1136) );
NAND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U813 ( .A(KEYINPUT30), .ZN(n1142) );
XOR2_X1 U814 ( .A(KEYINPUT16), .B(G125), .Z(n1141) );
XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(n1131) );
XOR2_X1 U816 ( .A(n1145), .B(n1146), .Z(n1143) );
NAND2_X1 U817 ( .A1(KEYINPUT39), .A2(n1147), .ZN(n1145) );
NAND2_X1 U818 ( .A1(n1148), .A2(n1149), .ZN(G69) );
NAND2_X1 U819 ( .A1(G953), .A2(n1150), .ZN(n1149) );
NAND2_X1 U820 ( .A1(n1151), .A2(G898), .ZN(n1150) );
XOR2_X1 U821 ( .A(n1152), .B(G224), .Z(n1151) );
NAND2_X1 U822 ( .A1(n1153), .A2(n1100), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1154), .B(n1155), .Z(n1153) );
INV_X1 U824 ( .A(n1152), .ZN(n1155) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U828 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
NOR2_X1 U829 ( .A1(n1158), .A2(n1164), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1165), .B(n1166), .ZN(n1164) );
AND2_X1 U831 ( .A1(G478), .A2(n1167), .ZN(n1166) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1168), .ZN(G60) );
XOR2_X1 U833 ( .A(n1169), .B(n1170), .Z(n1168) );
AND2_X1 U834 ( .A1(G475), .A2(n1167), .ZN(n1169) );
XOR2_X1 U835 ( .A(n1171), .B(G104), .Z(G6) );
NAND2_X1 U836 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U837 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U838 ( .A(KEYINPUT38), .ZN(n1175) );
NAND3_X1 U839 ( .A1(n1176), .A2(n1177), .A3(KEYINPUT38), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1178), .A2(n1179), .ZN(G57) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U842 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U843 ( .A(n1184), .B(n1185), .Z(n1180) );
AND2_X1 U844 ( .A1(G472), .A2(n1167), .ZN(n1185) );
NOR2_X1 U845 ( .A1(n1100), .A2(n1186), .ZN(n1178) );
XOR2_X1 U846 ( .A(KEYINPUT14), .B(G952), .Z(n1186) );
NOR2_X1 U847 ( .A1(n1158), .A2(n1187), .ZN(G54) );
NOR2_X1 U848 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U849 ( .A(KEYINPUT36), .B(n1190), .Z(n1189) );
NOR2_X1 U850 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
AND2_X1 U851 ( .A1(n1192), .A2(n1191), .ZN(n1188) );
XOR2_X1 U852 ( .A(n1193), .B(n1194), .Z(n1191) );
NAND2_X1 U853 ( .A1(KEYINPUT45), .A2(n1195), .ZN(n1193) );
NAND2_X1 U854 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U855 ( .A1(n1167), .A2(G469), .ZN(n1192) );
INV_X1 U856 ( .A(n1163), .ZN(n1167) );
NAND2_X1 U857 ( .A1(G902), .A2(n1067), .ZN(n1163) );
NOR2_X1 U858 ( .A1(n1158), .A2(n1198), .ZN(G51) );
XNOR2_X1 U859 ( .A(n1199), .B(n1200), .ZN(n1198) );
XOR2_X1 U860 ( .A(n1201), .B(n1202), .Z(n1199) );
NAND3_X1 U861 ( .A1(n1114), .A2(n1067), .A3(n1203), .ZN(n1201) );
XOR2_X1 U862 ( .A(n1204), .B(KEYINPUT24), .Z(n1203) );
NAND2_X1 U863 ( .A1(n1127), .A2(n1154), .ZN(n1067) );
AND4_X1 U864 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1154) );
AND4_X1 U865 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NOR2_X1 U866 ( .A1(n1174), .A2(n1213), .ZN(n1207) );
NOR2_X1 U867 ( .A1(n1214), .A2(n1061), .ZN(n1213) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1079), .ZN(n1061) );
XOR2_X1 U869 ( .A(n1060), .B(KEYINPUT57), .Z(n1214) );
NOR2_X1 U870 ( .A1(n1177), .A2(n1095), .ZN(n1174) );
INV_X1 U871 ( .A(n1176), .ZN(n1095) );
NAND4_X1 U872 ( .A1(n1080), .A2(n1082), .A3(n1216), .A4(n1217), .ZN(n1177) );
NAND3_X1 U873 ( .A1(n1218), .A2(n1080), .A3(n1219), .ZN(n1206) );
AND4_X1 U874 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1127) );
AND4_X1 U875 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
NOR2_X1 U876 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
NOR4_X1 U877 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1228) );
XOR2_X1 U878 ( .A(KEYINPUT6), .B(n1234), .Z(n1233) );
INV_X1 U879 ( .A(n1079), .ZN(n1230) );
NAND4_X1 U880 ( .A1(n1218), .A2(n1079), .A3(n1235), .A4(n1236), .ZN(n1220) );
OR2_X1 U881 ( .A1(n1237), .A2(KEYINPUT51), .ZN(n1236) );
NAND2_X1 U882 ( .A1(KEYINPUT51), .A2(n1238), .ZN(n1235) );
NAND2_X1 U883 ( .A1(n1234), .A2(n1087), .ZN(n1238) );
NOR2_X1 U884 ( .A1(n1100), .A2(G952), .ZN(n1158) );
XNOR2_X1 U885 ( .A(G146), .B(n1221), .ZN(G48) );
NAND4_X1 U886 ( .A1(n1239), .A2(n1080), .A3(n1240), .A4(n1241), .ZN(n1221) );
XNOR2_X1 U887 ( .A(G143), .B(n1227), .ZN(G45) );
NAND4_X1 U888 ( .A1(n1108), .A2(n1241), .A3(n1176), .A4(n1242), .ZN(n1227) );
AND3_X1 U889 ( .A1(n1218), .A2(n1240), .A3(n1243), .ZN(n1242) );
XOR2_X1 U890 ( .A(n1139), .B(n1226), .Z(G42) );
NAND3_X1 U891 ( .A1(n1080), .A2(n1244), .A3(n1237), .ZN(n1226) );
INV_X1 U892 ( .A(G140), .ZN(n1139) );
XOR2_X1 U893 ( .A(n1147), .B(n1225), .Z(G39) );
NAND3_X1 U894 ( .A1(n1076), .A2(n1245), .A3(n1237), .ZN(n1225) );
INV_X1 U895 ( .A(n1246), .ZN(n1237) );
XOR2_X1 U896 ( .A(G134), .B(n1247), .Z(G36) );
AND2_X1 U897 ( .A1(n1079), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U898 ( .A(G131), .B(n1224), .ZN(G33) );
NAND2_X1 U899 ( .A1(n1248), .A2(n1080), .ZN(n1224) );
NOR2_X1 U900 ( .A1(n1246), .A2(n1093), .ZN(n1248) );
INV_X1 U901 ( .A(n1218), .ZN(n1093) );
NAND2_X1 U902 ( .A1(n1087), .A2(n1241), .ZN(n1246) );
AND2_X1 U903 ( .A1(n1081), .A2(n1240), .ZN(n1087) );
AND2_X1 U904 ( .A1(n1098), .A2(n1249), .ZN(n1081) );
XNOR2_X1 U905 ( .A(G128), .B(n1250), .ZN(G30) );
NAND3_X1 U906 ( .A1(n1239), .A2(n1079), .A3(n1251), .ZN(n1250) );
NOR3_X1 U907 ( .A1(n1231), .A2(KEYINPUT49), .A3(n1234), .ZN(n1251) );
INV_X1 U908 ( .A(n1216), .ZN(n1231) );
INV_X1 U909 ( .A(n1232), .ZN(n1239) );
NAND2_X1 U910 ( .A1(n1176), .A2(n1245), .ZN(n1232) );
XNOR2_X1 U911 ( .A(G101), .B(n1212), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1218), .A2(n1215), .A3(n1076), .ZN(n1212) );
XNOR2_X1 U913 ( .A(G125), .B(n1252), .ZN(G27) );
NAND2_X1 U914 ( .A1(KEYINPUT29), .A2(n1229), .ZN(n1252) );
AND4_X1 U915 ( .A1(n1078), .A2(n1080), .A3(n1253), .A4(n1176), .ZN(n1229) );
NOR2_X1 U916 ( .A1(n1234), .A2(n1092), .ZN(n1253) );
INV_X1 U917 ( .A(n1244), .ZN(n1092) );
INV_X1 U918 ( .A(n1241), .ZN(n1234) );
NAND2_X1 U919 ( .A1(n1099), .A2(n1254), .ZN(n1241) );
NAND4_X1 U920 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1122), .ZN(n1254) );
INV_X1 U921 ( .A(G900), .ZN(n1122) );
NAND3_X1 U922 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(G24) );
NAND2_X1 U923 ( .A1(KEYINPUT44), .A2(n1205), .ZN(n1258) );
OR3_X1 U924 ( .A1(n1205), .A2(KEYINPUT44), .A3(G122), .ZN(n1257) );
NAND2_X1 U925 ( .A1(G122), .A2(n1259), .ZN(n1256) );
NAND2_X1 U926 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U927 ( .A(KEYINPUT44), .ZN(n1261) );
XNOR2_X1 U928 ( .A(KEYINPUT35), .B(n1205), .ZN(n1260) );
NAND4_X1 U929 ( .A1(n1243), .A2(n1219), .A3(n1082), .A4(n1108), .ZN(n1205) );
INV_X1 U930 ( .A(n1060), .ZN(n1082) );
NAND2_X1 U931 ( .A1(n1262), .A2(n1263), .ZN(n1060) );
XOR2_X1 U932 ( .A(n1264), .B(KEYINPUT37), .Z(n1262) );
XOR2_X1 U933 ( .A(n1211), .B(n1265), .Z(G21) );
NAND2_X1 U934 ( .A1(KEYINPUT26), .A2(G119), .ZN(n1265) );
NAND3_X1 U935 ( .A1(n1076), .A2(n1245), .A3(n1219), .ZN(n1211) );
XNOR2_X1 U936 ( .A(G116), .B(n1210), .ZN(G18) );
NAND3_X1 U937 ( .A1(n1218), .A2(n1079), .A3(n1219), .ZN(n1210) );
AND2_X1 U938 ( .A1(n1078), .A2(n1266), .ZN(n1219) );
NOR2_X1 U939 ( .A1(n1267), .A2(n1268), .ZN(n1079) );
XNOR2_X1 U940 ( .A(G113), .B(n1269), .ZN(G15) );
NAND4_X1 U941 ( .A1(n1218), .A2(n1080), .A3(n1266), .A4(n1270), .ZN(n1269) );
XOR2_X1 U942 ( .A(KEYINPUT55), .B(n1078), .Z(n1270) );
NOR2_X1 U943 ( .A1(n1110), .A2(n1077), .ZN(n1078) );
INV_X1 U944 ( .A(n1075), .ZN(n1110) );
AND2_X1 U945 ( .A1(n1243), .A2(n1271), .ZN(n1080) );
XNOR2_X1 U946 ( .A(KEYINPUT22), .B(n1268), .ZN(n1271) );
INV_X1 U947 ( .A(n1108), .ZN(n1268) );
XNOR2_X1 U948 ( .A(n1267), .B(KEYINPUT52), .ZN(n1243) );
XNOR2_X1 U949 ( .A(G110), .B(n1272), .ZN(G12) );
NAND2_X1 U950 ( .A1(KEYINPUT20), .A2(n1273), .ZN(n1272) );
INV_X1 U951 ( .A(n1209), .ZN(n1273) );
NAND3_X1 U952 ( .A1(n1215), .A2(n1244), .A3(n1076), .ZN(n1209) );
NOR2_X1 U953 ( .A1(n1108), .A2(n1267), .ZN(n1076) );
XOR2_X1 U954 ( .A(n1116), .B(G475), .Z(n1267) );
NOR2_X1 U955 ( .A1(n1170), .A2(n1274), .ZN(n1116) );
XNOR2_X1 U956 ( .A(n1275), .B(n1276), .ZN(n1170) );
XOR2_X1 U957 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U958 ( .A(n1279), .B(KEYINPUT19), .ZN(n1278) );
NAND2_X1 U959 ( .A1(n1280), .A2(KEYINPUT3), .ZN(n1279) );
XOR2_X1 U960 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U961 ( .A(G122), .B(G113), .Z(n1282) );
INV_X1 U962 ( .A(G104), .ZN(n1281) );
NOR2_X1 U963 ( .A1(n1283), .A2(n1284), .ZN(n1277) );
XOR2_X1 U964 ( .A(KEYINPUT46), .B(n1285), .Z(n1284) );
NOR2_X1 U965 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U966 ( .A(G143), .B(KEYINPUT56), .ZN(n1286) );
NOR2_X1 U967 ( .A1(G143), .A2(n1288), .ZN(n1283) );
INV_X1 U968 ( .A(n1287), .ZN(n1288) );
NAND2_X1 U969 ( .A1(G214), .A2(n1289), .ZN(n1287) );
XOR2_X1 U970 ( .A(n1290), .B(n1291), .Z(n1275) );
XNOR2_X1 U971 ( .A(n1292), .B(G478), .ZN(n1108) );
NAND2_X1 U972 ( .A1(n1293), .A2(n1165), .ZN(n1292) );
XNOR2_X1 U973 ( .A(n1294), .B(n1295), .ZN(n1165) );
XOR2_X1 U974 ( .A(G134), .B(n1296), .Z(n1295) );
NOR2_X1 U975 ( .A1(KEYINPUT27), .A2(n1297), .ZN(n1296) );
XOR2_X1 U976 ( .A(G122), .B(n1298), .Z(n1297) );
XOR2_X1 U977 ( .A(n1299), .B(n1300), .Z(n1294) );
AND2_X1 U978 ( .A1(G217), .A2(n1301), .ZN(n1300) );
XOR2_X1 U979 ( .A(n1274), .B(KEYINPUT2), .Z(n1293) );
NAND2_X1 U980 ( .A1(n1302), .A2(n1303), .ZN(n1244) );
NAND3_X1 U981 ( .A1(n1304), .A2(n1264), .A3(n1305), .ZN(n1303) );
INV_X1 U982 ( .A(KEYINPUT37), .ZN(n1305) );
XOR2_X1 U983 ( .A(KEYINPUT28), .B(n1107), .Z(n1304) );
NAND2_X1 U984 ( .A1(KEYINPUT37), .A2(n1245), .ZN(n1302) );
NAND2_X1 U985 ( .A1(n1306), .A2(n1307), .ZN(n1245) );
OR3_X1 U986 ( .A1(n1264), .A2(n1263), .A3(KEYINPUT28), .ZN(n1307) );
NAND2_X1 U987 ( .A1(KEYINPUT28), .A2(n1218), .ZN(n1306) );
NOR2_X1 U988 ( .A1(n1107), .A2(n1264), .ZN(n1218) );
XOR2_X1 U989 ( .A(n1308), .B(n1112), .Z(n1264) );
XOR2_X1 U990 ( .A(G472), .B(KEYINPUT58), .Z(n1112) );
NAND2_X1 U991 ( .A1(KEYINPUT8), .A2(n1111), .ZN(n1308) );
NAND2_X1 U992 ( .A1(n1309), .A2(n1310), .ZN(n1111) );
XOR2_X1 U993 ( .A(n1311), .B(n1183), .Z(n1309) );
XNOR2_X1 U994 ( .A(n1312), .B(n1313), .ZN(n1183) );
XNOR2_X1 U995 ( .A(n1314), .B(n1315), .ZN(n1313) );
NAND2_X1 U996 ( .A1(G210), .A2(n1289), .ZN(n1314) );
NOR2_X1 U997 ( .A1(G953), .A2(G237), .ZN(n1289) );
XOR2_X1 U998 ( .A(n1316), .B(G131), .Z(n1312) );
XNOR2_X1 U999 ( .A(n1182), .B(n1317), .ZN(n1311) );
NOR2_X1 U1000 ( .A1(KEYINPUT4), .A2(n1318), .ZN(n1317) );
INV_X1 U1001 ( .A(n1263), .ZN(n1107) );
XNOR2_X1 U1002 ( .A(n1319), .B(n1162), .ZN(n1263) );
NAND2_X1 U1003 ( .A1(G217), .A2(n1320), .ZN(n1162) );
NAND2_X1 U1004 ( .A1(n1161), .A2(n1310), .ZN(n1319) );
NAND2_X1 U1005 ( .A1(n1321), .A2(n1322), .ZN(n1161) );
NAND2_X1 U1006 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1007 ( .A(KEYINPUT21), .B(n1325), .Z(n1323) );
NAND2_X1 U1008 ( .A1(n1326), .A2(n1327), .ZN(n1321) );
INV_X1 U1009 ( .A(n1324), .ZN(n1327) );
XOR2_X1 U1010 ( .A(n1328), .B(n1329), .Z(n1324) );
XOR2_X1 U1011 ( .A(G128), .B(n1330), .Z(n1329) );
XOR2_X1 U1012 ( .A(KEYINPUT32), .B(G146), .Z(n1330) );
XOR2_X1 U1013 ( .A(n1331), .B(n1291), .Z(n1328) );
XOR2_X1 U1014 ( .A(G140), .B(G125), .Z(n1291) );
XOR2_X1 U1015 ( .A(n1332), .B(G110), .Z(n1331) );
NAND2_X1 U1016 ( .A1(KEYINPUT40), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1017 ( .A(KEYINPUT23), .B(n1325), .Z(n1326) );
XOR2_X1 U1018 ( .A(n1334), .B(n1147), .Z(n1325) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1301), .ZN(n1334) );
AND2_X1 U1020 ( .A1(G234), .A2(n1100), .ZN(n1301) );
AND2_X1 U1021 ( .A1(n1266), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U1022 ( .A(n1240), .B(KEYINPUT43), .ZN(n1216) );
NOR2_X1 U1023 ( .A1(n1075), .A2(n1077), .ZN(n1240) );
AND2_X1 U1024 ( .A1(G221), .A2(n1320), .ZN(n1077) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1335), .ZN(n1320) );
XOR2_X1 U1026 ( .A(KEYINPUT15), .B(G902), .Z(n1335) );
XOR2_X1 U1027 ( .A(n1336), .B(G469), .Z(n1075) );
NAND2_X1 U1028 ( .A1(n1337), .A2(n1310), .ZN(n1336) );
XNOR2_X1 U1029 ( .A(n1194), .B(n1338), .ZN(n1337) );
XOR2_X1 U1030 ( .A(KEYINPUT25), .B(n1339), .Z(n1338) );
NOR2_X1 U1031 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1032 ( .A(n1196), .B(KEYINPUT0), .Z(n1341) );
OR3_X1 U1033 ( .A1(n1121), .A2(G953), .A3(n1342), .ZN(n1196) );
INV_X1 U1034 ( .A(G227), .ZN(n1121) );
INV_X1 U1035 ( .A(n1197), .ZN(n1340) );
NAND2_X1 U1036 ( .A1(n1342), .A2(n1343), .ZN(n1197) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1100), .ZN(n1343) );
XOR2_X1 U1038 ( .A(G110), .B(G140), .Z(n1342) );
XNOR2_X1 U1039 ( .A(n1344), .B(n1345), .ZN(n1194) );
XOR2_X1 U1040 ( .A(n1144), .B(n1315), .Z(n1345) );
INV_X1 U1041 ( .A(n1290), .ZN(n1144) );
XNOR2_X1 U1042 ( .A(G131), .B(G146), .ZN(n1290) );
XOR2_X1 U1043 ( .A(n1346), .B(n1347), .Z(n1344) );
INV_X1 U1044 ( .A(n1299), .ZN(n1347) );
XNOR2_X1 U1045 ( .A(G107), .B(n1146), .ZN(n1299) );
XOR2_X1 U1046 ( .A(G128), .B(G143), .Z(n1146) );
XOR2_X1 U1047 ( .A(n1316), .B(G104), .Z(n1346) );
NAND3_X1 U1048 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1316) );
NAND2_X1 U1049 ( .A1(G134), .A2(n1147), .ZN(n1350) );
INV_X1 U1050 ( .A(G137), .ZN(n1147) );
NAND2_X1 U1051 ( .A1(KEYINPUT62), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1052 ( .A1(G137), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1053 ( .A(KEYINPUT5), .B(G134), .Z(n1352) );
NAND2_X1 U1054 ( .A1(n1353), .A2(n1354), .ZN(n1348) );
INV_X1 U1055 ( .A(KEYINPUT62), .ZN(n1354) );
NAND2_X1 U1056 ( .A1(n1355), .A2(n1356), .ZN(n1353) );
OR2_X1 U1057 ( .A1(n1135), .A2(KEYINPUT5), .ZN(n1356) );
NAND3_X1 U1058 ( .A1(G137), .A2(n1135), .A3(KEYINPUT5), .ZN(n1355) );
INV_X1 U1059 ( .A(G134), .ZN(n1135) );
AND2_X1 U1060 ( .A1(n1176), .A2(n1217), .ZN(n1266) );
NAND2_X1 U1061 ( .A1(n1357), .A2(n1099), .ZN(n1217) );
NAND3_X1 U1062 ( .A1(n1255), .A2(n1100), .A3(G952), .ZN(n1099) );
NAND4_X1 U1063 ( .A1(n1358), .A2(G902), .A3(n1255), .A4(n1359), .ZN(n1357) );
INV_X1 U1064 ( .A(G898), .ZN(n1359) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1255) );
XOR2_X1 U1066 ( .A(n1100), .B(KEYINPUT41), .Z(n1358) );
NOR2_X1 U1067 ( .A1(n1098), .A2(n1097), .ZN(n1176) );
INV_X1 U1068 ( .A(n1249), .ZN(n1097) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1360), .ZN(n1249) );
NOR2_X1 U1070 ( .A1(n1113), .A2(n1361), .ZN(n1098) );
AND2_X1 U1071 ( .A1(n1362), .A2(n1115), .ZN(n1361) );
XOR2_X1 U1072 ( .A(KEYINPUT18), .B(n1114), .Z(n1362) );
NOR2_X1 U1073 ( .A1(n1115), .A2(n1114), .ZN(n1113) );
AND2_X1 U1074 ( .A1(G210), .A2(n1360), .ZN(n1114) );
NAND2_X1 U1075 ( .A1(n1363), .A2(n1204), .ZN(n1360) );
XOR2_X1 U1076 ( .A(KEYINPUT48), .B(G237), .Z(n1363) );
NAND2_X1 U1077 ( .A1(n1364), .A2(n1310), .ZN(n1115) );
INV_X1 U1078 ( .A(n1274), .ZN(n1310) );
XOR2_X1 U1079 ( .A(n1204), .B(KEYINPUT1), .Z(n1274) );
INV_X1 U1080 ( .A(G902), .ZN(n1204) );
XOR2_X1 U1081 ( .A(n1365), .B(KEYINPUT9), .Z(n1364) );
NAND3_X1 U1082 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1365) );
NAND2_X1 U1083 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
INV_X1 U1084 ( .A(KEYINPUT53), .ZN(n1370) );
NAND3_X1 U1085 ( .A1(KEYINPUT53), .A2(n1371), .A3(n1200), .ZN(n1367) );
OR2_X1 U1086 ( .A1(n1200), .A2(n1371), .ZN(n1366) );
NOR2_X1 U1087 ( .A1(n1372), .A2(n1369), .ZN(n1371) );
XOR2_X1 U1088 ( .A(n1202), .B(KEYINPUT31), .Z(n1369) );
XNOR2_X1 U1089 ( .A(n1373), .B(n1374), .ZN(n1202) );
XOR2_X1 U1090 ( .A(KEYINPUT59), .B(G125), .Z(n1374) );
XOR2_X1 U1091 ( .A(n1375), .B(n1318), .Z(n1373) );
INV_X1 U1092 ( .A(n1184), .ZN(n1318) );
XOR2_X1 U1093 ( .A(n1376), .B(G128), .Z(n1184) );
NAND2_X1 U1094 ( .A1(KEYINPUT63), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1095 ( .A(G146), .B(G143), .Z(n1377) );
NAND2_X1 U1096 ( .A1(G224), .A2(n1100), .ZN(n1375) );
INV_X1 U1097 ( .A(G953), .ZN(n1100) );
INV_X1 U1098 ( .A(KEYINPUT12), .ZN(n1372) );
NAND2_X1 U1099 ( .A1(n1378), .A2(n1379), .ZN(n1200) );
NAND2_X1 U1100 ( .A1(n1157), .A2(n1156), .ZN(n1379) );
INV_X1 U1101 ( .A(n1380), .ZN(n1157) );
NAND2_X1 U1102 ( .A1(n1381), .A2(n1380), .ZN(n1378) );
NAND3_X1 U1103 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n1380) );
OR2_X1 U1104 ( .A1(n1385), .A2(KEYINPUT10), .ZN(n1384) );
OR3_X1 U1105 ( .A1(n1386), .A2(n1387), .A3(n1315), .ZN(n1383) );
INV_X1 U1106 ( .A(KEYINPUT10), .ZN(n1386) );
NAND2_X1 U1107 ( .A1(n1315), .A2(n1387), .ZN(n1382) );
NAND2_X1 U1108 ( .A1(KEYINPUT34), .A2(n1385), .ZN(n1387) );
XOR2_X1 U1109 ( .A(G107), .B(G104), .Z(n1385) );
XOR2_X1 U1110 ( .A(G101), .B(KEYINPUT33), .Z(n1315) );
XOR2_X1 U1111 ( .A(n1156), .B(KEYINPUT11), .Z(n1381) );
XNOR2_X1 U1112 ( .A(n1182), .B(n1388), .ZN(n1156) );
XOR2_X1 U1113 ( .A(G122), .B(G110), .Z(n1388) );
XOR2_X1 U1114 ( .A(n1389), .B(n1333), .Z(n1182) );
XNOR2_X1 U1115 ( .A(G119), .B(KEYINPUT50), .ZN(n1333) );
XNOR2_X1 U1116 ( .A(G113), .B(n1298), .ZN(n1389) );
XOR2_X1 U1117 ( .A(G116), .B(KEYINPUT42), .Z(n1298) );
endmodule


