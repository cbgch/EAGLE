//Key = 1011111010110011000000110000010011100111011001001110010100110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345;

XOR2_X1 U733 ( .A(n1021), .B(n1022), .Z(G9) );
NOR2_X1 U734 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR4_X1 U735 ( .A1(G953), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1024) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR3_X1 U738 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR2_X1 U739 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U740 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR3_X1 U741 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1035) );
NOR3_X1 U742 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR2_X1 U743 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
NOR4_X1 U744 ( .A1(n1047), .A2(n1042), .A3(n1039), .A4(n1038), .ZN(n1030) );
INV_X1 U745 ( .A(n1045), .ZN(n1038) );
NOR2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U747 ( .A1(n1050), .A2(n1034), .ZN(n1049) );
NOR2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U749 ( .A(KEYINPUT28), .B(n1053), .Z(n1052) );
NOR2_X1 U750 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
NOR2_X1 U751 ( .A1(n1056), .A2(n1032), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR3_X1 U754 ( .A1(n1025), .A2(G953), .A3(G952), .ZN(n1023) );
AND4_X1 U755 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1025) );
XOR2_X1 U756 ( .A(KEYINPUT55), .B(n1059), .Z(n1064) );
AND2_X1 U757 ( .A1(n1060), .A2(n1055), .ZN(n1063) );
XOR2_X1 U758 ( .A(n1065), .B(KEYINPUT23), .Z(n1061) );
NAND4_X1 U759 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1065) );
NOR2_X1 U760 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U761 ( .A(G475), .B(n1072), .Z(n1071) );
XNOR2_X1 U762 ( .A(n1073), .B(n1074), .ZN(n1070) );
NOR2_X1 U763 ( .A1(KEYINPUT26), .A2(n1075), .ZN(n1074) );
XOR2_X1 U764 ( .A(G478), .B(n1076), .Z(n1068) );
NOR2_X1 U765 ( .A1(n1077), .A2(KEYINPUT52), .ZN(n1076) );
XNOR2_X1 U766 ( .A(KEYINPUT32), .B(n1078), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
AND2_X1 U769 ( .A1(G227), .A2(G900), .ZN(n1081) );
NAND2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1079) );
NAND3_X1 U771 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
INV_X1 U772 ( .A(n1088), .ZN(n1086) );
OR2_X1 U773 ( .A1(n1085), .A2(n1087), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1089), .ZN(n1087) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U776 ( .A(KEYINPUT7), .B(n1092), .Z(n1091) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1085) );
XOR2_X1 U778 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U779 ( .A(n1097), .B(n1098), .ZN(n1096) );
NAND2_X1 U780 ( .A1(KEYINPUT41), .A2(n1099), .ZN(n1097) );
XOR2_X1 U781 ( .A(n1100), .B(G134), .Z(n1093) );
XNOR2_X1 U782 ( .A(KEYINPUT6), .B(KEYINPUT29), .ZN(n1100) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(G69) );
XOR2_X1 U784 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U785 ( .A1(n1082), .A2(n1105), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U787 ( .A(n1108), .B(KEYINPUT37), .ZN(n1106) );
NAND2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1103) );
NAND2_X1 U789 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U790 ( .A(n1112), .B(n1113), .Z(n1109) );
XOR2_X1 U791 ( .A(n1114), .B(KEYINPUT30), .Z(n1112) );
NOR2_X1 U792 ( .A1(n1115), .A2(n1082), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1116), .A2(n1111), .ZN(n1115) );
NOR2_X1 U794 ( .A1(n1117), .A2(n1118), .ZN(G66) );
NOR3_X1 U795 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NOR3_X1 U796 ( .A1(n1122), .A2(n1073), .A3(n1123), .ZN(n1121) );
NOR2_X1 U797 ( .A1(n1124), .A2(n1125), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1126), .A2(n1073), .ZN(n1124) );
INV_X1 U799 ( .A(n1027), .ZN(n1126) );
INV_X1 U800 ( .A(n1075), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(G63) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U803 ( .A1(n1131), .A2(G478), .ZN(n1129) );
XNOR2_X1 U804 ( .A(n1117), .B(KEYINPUT58), .ZN(n1127) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1132), .ZN(G60) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U807 ( .A1(n1131), .A2(G475), .ZN(n1133) );
XNOR2_X1 U808 ( .A(G104), .B(n1135), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1117), .A2(n1136), .ZN(G57) );
NOR3_X1 U810 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR2_X1 U811 ( .A1(G101), .A2(n1140), .ZN(n1139) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR3_X1 U813 ( .A1(n1143), .A2(n1144), .A3(n1142), .ZN(n1138) );
INV_X1 U814 ( .A(n1141), .ZN(n1144) );
AND2_X1 U815 ( .A1(n1142), .A2(n1145), .ZN(n1137) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(n1142) );
NAND2_X1 U817 ( .A1(n1131), .A2(G472), .ZN(n1146) );
NOR2_X1 U818 ( .A1(n1117), .A2(n1148), .ZN(G54) );
NOR2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U820 ( .A(KEYINPUT24), .B(n1151), .Z(n1150) );
NOR3_X1 U821 ( .A1(n1152), .A2(n1153), .A3(n1123), .ZN(n1151) );
XOR2_X1 U822 ( .A(KEYINPUT39), .B(n1154), .Z(n1152) );
NOR2_X1 U823 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1153), .A2(n1123), .ZN(n1155) );
INV_X1 U825 ( .A(G469), .ZN(n1153) );
AND2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U828 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U829 ( .A(n1162), .B(n1163), .Z(n1158) );
XOR2_X1 U830 ( .A(n1164), .B(KEYINPUT46), .Z(n1156) );
NAND2_X1 U831 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XNOR2_X1 U832 ( .A(n1162), .B(n1163), .ZN(n1166) );
XOR2_X1 U833 ( .A(G140), .B(n1167), .Z(n1163) );
NOR2_X1 U834 ( .A1(KEYINPUT16), .A2(n1168), .ZN(n1167) );
OR2_X1 U835 ( .A1(n1169), .A2(KEYINPUT20), .ZN(n1162) );
XOR2_X1 U836 ( .A(n1170), .B(n1160), .Z(n1165) );
NOR2_X1 U837 ( .A1(KEYINPUT40), .A2(n1171), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1117), .A2(n1172), .ZN(G51) );
XOR2_X1 U839 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U841 ( .A1(n1131), .A2(n1177), .ZN(n1176) );
INV_X1 U842 ( .A(n1123), .ZN(n1131) );
NAND2_X1 U843 ( .A1(G902), .A2(n1027), .ZN(n1123) );
NAND4_X1 U844 ( .A1(n1092), .A2(n1108), .A3(n1107), .A4(n1090), .ZN(n1027) );
AND4_X1 U845 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1090) );
AND4_X1 U846 ( .A1(n1182), .A2(n1135), .A3(n1183), .A4(n1022), .ZN(n1107) );
NAND2_X1 U847 ( .A1(n1044), .A2(n1184), .ZN(n1022) );
NAND2_X1 U848 ( .A1(n1043), .A2(n1184), .ZN(n1135) );
AND3_X1 U849 ( .A1(n1046), .A2(n1185), .A3(n1186), .ZN(n1184) );
OR2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1182) );
AND4_X1 U851 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1108) );
OR2_X1 U852 ( .A1(n1193), .A2(n1194), .ZN(n1190) );
AND4_X1 U853 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1092) );
NAND3_X1 U854 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
NAND2_X1 U855 ( .A1(n1202), .A2(n1039), .ZN(n1200) );
NAND3_X1 U856 ( .A1(n1044), .A2(n1203), .A3(KEYINPUT57), .ZN(n1202) );
NAND2_X1 U857 ( .A1(n1186), .A2(n1204), .ZN(n1199) );
OR2_X1 U858 ( .A1(n1205), .A2(n1034), .ZN(n1204) );
NAND2_X1 U859 ( .A1(n1206), .A2(n1207), .ZN(n1197) );
NAND2_X1 U860 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND4_X1 U861 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1044), .ZN(n1209) );
NOR2_X1 U862 ( .A1(KEYINPUT34), .A2(n1203), .ZN(n1212) );
NAND3_X1 U863 ( .A1(n1043), .A2(n1213), .A3(n1214), .ZN(n1208) );
XOR2_X1 U864 ( .A(KEYINPUT17), .B(n1210), .Z(n1213) );
NAND2_X1 U865 ( .A1(KEYINPUT34), .A2(n1215), .ZN(n1196) );
NAND2_X1 U866 ( .A1(n1216), .A2(n1217), .ZN(n1195) );
INV_X1 U867 ( .A(KEYINPUT57), .ZN(n1217) );
NAND2_X1 U868 ( .A1(n1218), .A2(n1219), .ZN(n1175) );
NAND2_X1 U869 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XOR2_X1 U870 ( .A(KEYINPUT49), .B(n1222), .Z(n1218) );
NOR2_X1 U871 ( .A1(n1220), .A2(n1221), .ZN(n1222) );
XNOR2_X1 U872 ( .A(KEYINPUT33), .B(G125), .ZN(n1220) );
NOR2_X1 U873 ( .A1(n1082), .A2(G952), .ZN(n1117) );
XNOR2_X1 U874 ( .A(G146), .B(n1178), .ZN(G48) );
NAND3_X1 U875 ( .A1(n1043), .A2(n1053), .A3(n1223), .ZN(n1178) );
XOR2_X1 U876 ( .A(G143), .B(n1224), .Z(G45) );
NOR2_X1 U877 ( .A1(KEYINPUT36), .A2(n1179), .ZN(n1224) );
NAND2_X1 U878 ( .A1(n1225), .A2(n1226), .ZN(n1179) );
XNOR2_X1 U879 ( .A(G140), .B(n1180), .ZN(G42) );
NAND3_X1 U880 ( .A1(n1206), .A2(n1214), .A3(n1227), .ZN(n1180) );
NOR3_X1 U881 ( .A1(n1205), .A2(n1046), .A3(n1039), .ZN(n1227) );
XOR2_X1 U882 ( .A(n1228), .B(n1181), .Z(G39) );
NAND3_X1 U883 ( .A1(n1223), .A2(n1206), .A3(n1045), .ZN(n1181) );
XOR2_X1 U884 ( .A(n1229), .B(n1215), .Z(G36) );
AND3_X1 U885 ( .A1(n1206), .A2(n1044), .A3(n1226), .ZN(n1215) );
INV_X1 U886 ( .A(n1032), .ZN(n1206) );
NAND2_X1 U887 ( .A1(KEYINPUT22), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U888 ( .A(G131), .B(n1231), .ZN(G33) );
NAND3_X1 U889 ( .A1(n1226), .A2(n1043), .A3(n1232), .ZN(n1231) );
XOR2_X1 U890 ( .A(n1032), .B(KEYINPUT0), .Z(n1232) );
NAND2_X1 U891 ( .A1(n1233), .A2(n1055), .ZN(n1032) );
INV_X1 U892 ( .A(n1054), .ZN(n1233) );
AND2_X1 U893 ( .A1(n1214), .A2(n1210), .ZN(n1226) );
XOR2_X1 U894 ( .A(G128), .B(n1216), .Z(G30) );
AND3_X1 U895 ( .A1(n1044), .A2(n1053), .A3(n1223), .ZN(n1216) );
AND3_X1 U896 ( .A1(n1042), .A2(n1039), .A3(n1214), .ZN(n1223) );
NOR2_X1 U897 ( .A1(n1203), .A2(n1211), .ZN(n1214) );
XOR2_X1 U898 ( .A(G101), .B(n1234), .Z(G3) );
NOR2_X1 U899 ( .A1(KEYINPUT9), .A2(n1183), .ZN(n1234) );
NAND3_X1 U900 ( .A1(n1210), .A2(n1185), .A3(n1045), .ZN(n1183) );
NOR3_X1 U901 ( .A1(n1203), .A2(n1235), .A3(n1188), .ZN(n1185) );
XNOR2_X1 U902 ( .A(G125), .B(n1236), .ZN(G27) );
NAND3_X1 U903 ( .A1(KEYINPUT2), .A2(n1201), .A3(n1237), .ZN(n1236) );
NOR3_X1 U904 ( .A1(n1205), .A2(n1039), .A3(n1034), .ZN(n1237) );
NOR3_X1 U905 ( .A1(n1046), .A2(n1211), .A3(n1194), .ZN(n1201) );
AND2_X1 U906 ( .A1(n1238), .A2(n1029), .ZN(n1211) );
NAND3_X1 U907 ( .A1(G902), .A2(n1239), .A3(n1088), .ZN(n1238) );
NOR2_X1 U908 ( .A1(n1082), .A2(G900), .ZN(n1088) );
XOR2_X1 U909 ( .A(n1191), .B(n1240), .Z(G24) );
XOR2_X1 U910 ( .A(KEYINPUT11), .B(G122), .Z(n1240) );
NAND4_X1 U911 ( .A1(n1225), .A2(n1241), .A3(n1046), .A4(n1186), .ZN(n1191) );
AND3_X1 U912 ( .A1(n1242), .A2(n1243), .A3(n1053), .ZN(n1225) );
XOR2_X1 U913 ( .A(G119), .B(n1244), .Z(G21) );
NOR2_X1 U914 ( .A1(n1194), .A2(n1245), .ZN(n1244) );
XOR2_X1 U915 ( .A(n1193), .B(KEYINPUT51), .Z(n1245) );
NAND4_X1 U916 ( .A1(n1045), .A2(n1241), .A3(n1042), .A4(n1039), .ZN(n1193) );
XNOR2_X1 U917 ( .A(G116), .B(n1192), .ZN(G18) );
NAND4_X1 U918 ( .A1(n1241), .A2(n1210), .A3(n1044), .A4(n1053), .ZN(n1192) );
INV_X1 U919 ( .A(n1194), .ZN(n1053) );
XOR2_X1 U920 ( .A(n1188), .B(KEYINPUT44), .Z(n1194) );
NOR2_X1 U921 ( .A1(n1243), .A2(n1246), .ZN(n1044) );
XOR2_X1 U922 ( .A(n1247), .B(n1248), .Z(G15) );
XOR2_X1 U923 ( .A(n1249), .B(KEYINPUT1), .Z(n1248) );
NAND2_X1 U924 ( .A1(KEYINPUT15), .A2(n1250), .ZN(n1247) );
INV_X1 U925 ( .A(n1189), .ZN(n1250) );
NAND4_X1 U926 ( .A1(n1241), .A2(n1210), .A3(n1043), .A4(n1251), .ZN(n1189) );
INV_X1 U927 ( .A(n1205), .ZN(n1043) );
NAND2_X1 U928 ( .A1(n1246), .A2(n1243), .ZN(n1205) );
INV_X1 U929 ( .A(n1037), .ZN(n1210) );
NAND2_X1 U930 ( .A1(n1252), .A2(n1039), .ZN(n1037) );
XOR2_X1 U931 ( .A(KEYINPUT59), .B(n1042), .Z(n1252) );
INV_X1 U932 ( .A(n1046), .ZN(n1042) );
NOR2_X1 U933 ( .A1(n1034), .A2(n1235), .ZN(n1241) );
NAND2_X1 U934 ( .A1(n1253), .A2(n1060), .ZN(n1034) );
XOR2_X1 U935 ( .A(n1168), .B(n1254), .Z(G12) );
NAND2_X1 U936 ( .A1(n1255), .A2(n1251), .ZN(n1254) );
INV_X1 U937 ( .A(n1188), .ZN(n1251) );
NAND2_X1 U938 ( .A1(n1054), .A2(n1055), .ZN(n1188) );
NAND2_X1 U939 ( .A1(G214), .A2(n1256), .ZN(n1055) );
XNOR2_X1 U940 ( .A(n1062), .B(KEYINPUT47), .ZN(n1054) );
XOR2_X1 U941 ( .A(n1257), .B(n1177), .Z(n1062) );
AND2_X1 U942 ( .A1(G210), .A2(n1256), .ZN(n1177) );
NAND2_X1 U943 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
INV_X1 U944 ( .A(G237), .ZN(n1258) );
NAND2_X1 U945 ( .A1(n1260), .A2(n1259), .ZN(n1257) );
XOR2_X1 U946 ( .A(n1173), .B(n1261), .Z(n1260) );
XNOR2_X1 U947 ( .A(n1221), .B(G125), .ZN(n1261) );
XOR2_X1 U948 ( .A(n1262), .B(n1263), .Z(n1173) );
XOR2_X1 U949 ( .A(KEYINPUT54), .B(n1264), .Z(n1263) );
NOR2_X1 U950 ( .A1(n1116), .A2(n1265), .ZN(n1264) );
XOR2_X1 U951 ( .A(KEYINPUT43), .B(G953), .Z(n1265) );
INV_X1 U952 ( .A(G224), .ZN(n1116) );
XOR2_X1 U953 ( .A(n1266), .B(n1113), .Z(n1262) );
XNOR2_X1 U954 ( .A(n1267), .B(n1268), .ZN(n1113) );
XOR2_X1 U955 ( .A(G122), .B(G110), .Z(n1268) );
XOR2_X1 U956 ( .A(n1269), .B(n1270), .Z(n1267) );
NAND2_X1 U957 ( .A1(KEYINPUT48), .A2(G119), .ZN(n1269) );
NAND2_X1 U958 ( .A1(KEYINPUT5), .A2(n1114), .ZN(n1266) );
NAND2_X1 U959 ( .A1(n1271), .A2(n1272), .ZN(n1114) );
NAND2_X1 U960 ( .A1(G101), .A2(n1273), .ZN(n1272) );
XOR2_X1 U961 ( .A(KEYINPUT10), .B(n1274), .Z(n1271) );
NOR2_X1 U962 ( .A1(G101), .A2(n1273), .ZN(n1274) );
XOR2_X1 U963 ( .A(n1187), .B(KEYINPUT61), .Z(n1255) );
NAND4_X1 U964 ( .A1(n1045), .A2(n1186), .A3(n1275), .A4(n1058), .ZN(n1187) );
INV_X1 U965 ( .A(n1203), .ZN(n1058) );
NAND2_X1 U966 ( .A1(n1059), .A2(n1060), .ZN(n1203) );
NAND2_X1 U967 ( .A1(G221), .A2(n1276), .ZN(n1060) );
INV_X1 U968 ( .A(n1253), .ZN(n1059) );
XOR2_X1 U969 ( .A(n1277), .B(n1278), .Z(n1253) );
XOR2_X1 U970 ( .A(KEYINPUT27), .B(G469), .Z(n1278) );
NAND2_X1 U971 ( .A1(n1279), .A2(n1259), .ZN(n1277) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U973 ( .A(n1170), .B(n1171), .Z(n1281) );
XNOR2_X1 U974 ( .A(n1282), .B(n1098), .ZN(n1171) );
XOR2_X1 U975 ( .A(G128), .B(n1283), .Z(n1098) );
NOR2_X1 U976 ( .A1(KEYINPUT35), .A2(n1284), .ZN(n1283) );
XOR2_X1 U977 ( .A(G146), .B(n1285), .Z(n1284) );
NAND3_X1 U978 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1282) );
NAND2_X1 U979 ( .A1(KEYINPUT21), .A2(n1289), .ZN(n1288) );
NAND3_X1 U980 ( .A1(n1290), .A2(n1291), .A3(n1143), .ZN(n1287) );
INV_X1 U981 ( .A(KEYINPUT21), .ZN(n1291) );
OR2_X1 U982 ( .A1(n1143), .A2(n1290), .ZN(n1286) );
NOR2_X1 U983 ( .A1(KEYINPUT25), .A2(n1289), .ZN(n1290) );
INV_X1 U984 ( .A(n1273), .ZN(n1289) );
XOR2_X1 U985 ( .A(G104), .B(G107), .Z(n1273) );
XNOR2_X1 U986 ( .A(n1169), .B(n1292), .ZN(n1280) );
XOR2_X1 U987 ( .A(G140), .B(G110), .Z(n1292) );
AND2_X1 U988 ( .A1(G227), .A2(n1082), .ZN(n1169) );
NOR2_X1 U989 ( .A1(n1235), .A2(n1046), .ZN(n1275) );
XNOR2_X1 U990 ( .A(n1293), .B(n1073), .ZN(n1046) );
NAND2_X1 U991 ( .A1(G217), .A2(n1276), .ZN(n1073) );
NAND2_X1 U992 ( .A1(n1294), .A2(n1259), .ZN(n1276) );
XOR2_X1 U993 ( .A(n1075), .B(KEYINPUT18), .Z(n1293) );
NAND2_X1 U994 ( .A1(n1122), .A2(n1259), .ZN(n1075) );
INV_X1 U995 ( .A(n1125), .ZN(n1122) );
XOR2_X1 U996 ( .A(n1295), .B(n1296), .Z(n1125) );
XOR2_X1 U997 ( .A(n1297), .B(n1298), .Z(n1296) );
NAND2_X1 U998 ( .A1(G221), .A2(n1299), .ZN(n1297) );
XOR2_X1 U999 ( .A(n1300), .B(n1301), .Z(n1295) );
NOR2_X1 U1000 ( .A1(KEYINPUT13), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1001 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1002 ( .A(G128), .B(n1305), .Z(n1304) );
NAND2_X1 U1003 ( .A1(KEYINPUT62), .A2(n1168), .ZN(n1303) );
XOR2_X1 U1004 ( .A(n1228), .B(G146), .Z(n1300) );
INV_X1 U1005 ( .A(G137), .ZN(n1228) );
AND2_X1 U1006 ( .A1(n1029), .A2(n1306), .ZN(n1235) );
NAND4_X1 U1007 ( .A1(G902), .A2(G953), .A3(n1239), .A4(n1111), .ZN(n1306) );
INV_X1 U1008 ( .A(G898), .ZN(n1111) );
NAND3_X1 U1009 ( .A1(n1239), .A2(n1082), .A3(G952), .ZN(n1029) );
NAND2_X1 U1010 ( .A1(G237), .A2(n1294), .ZN(n1239) );
XOR2_X1 U1011 ( .A(G234), .B(KEYINPUT63), .Z(n1294) );
INV_X1 U1012 ( .A(n1039), .ZN(n1186) );
NAND2_X1 U1013 ( .A1(n1078), .A2(n1067), .ZN(n1039) );
NAND3_X1 U1014 ( .A1(n1307), .A2(n1259), .A3(n1308), .ZN(n1067) );
INV_X1 U1015 ( .A(G472), .ZN(n1307) );
NAND2_X1 U1016 ( .A1(G472), .A2(n1309), .ZN(n1078) );
NAND2_X1 U1017 ( .A1(n1308), .A2(n1259), .ZN(n1309) );
XNOR2_X1 U1018 ( .A(n1147), .B(n1310), .ZN(n1308) );
XOR2_X1 U1019 ( .A(KEYINPUT4), .B(n1311), .Z(n1310) );
NOR2_X1 U1020 ( .A1(n1145), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1021 ( .A(n1313), .B(KEYINPUT50), .Z(n1312) );
NAND2_X1 U1022 ( .A1(n1314), .A2(n1143), .ZN(n1313) );
XOR2_X1 U1023 ( .A(n1141), .B(KEYINPUT12), .Z(n1314) );
NOR2_X1 U1024 ( .A1(n1143), .A2(n1141), .ZN(n1145) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1315), .ZN(n1141) );
INV_X1 U1026 ( .A(G101), .ZN(n1143) );
XNOR2_X1 U1027 ( .A(n1316), .B(n1221), .ZN(n1147) );
XOR2_X1 U1028 ( .A(G146), .B(n1317), .Z(n1221) );
XOR2_X1 U1029 ( .A(n1318), .B(n1161), .Z(n1316) );
INV_X1 U1030 ( .A(n1170), .ZN(n1161) );
XNOR2_X1 U1031 ( .A(n1095), .B(n1319), .ZN(n1170) );
NOR2_X1 U1032 ( .A1(G134), .A2(KEYINPUT19), .ZN(n1319) );
XOR2_X1 U1033 ( .A(G131), .B(G137), .Z(n1095) );
NAND3_X1 U1034 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1318) );
NAND3_X1 U1035 ( .A1(G116), .A2(n1305), .A3(G113), .ZN(n1322) );
INV_X1 U1036 ( .A(G119), .ZN(n1305) );
OR3_X1 U1037 ( .A1(G113), .A2(G116), .A3(G119), .ZN(n1321) );
NAND2_X1 U1038 ( .A1(n1270), .A2(G119), .ZN(n1320) );
XOR2_X1 U1039 ( .A(G113), .B(G116), .Z(n1270) );
NOR2_X1 U1040 ( .A1(n1242), .A2(n1243), .ZN(n1045) );
XNOR2_X1 U1041 ( .A(n1323), .B(G475), .ZN(n1243) );
NAND2_X1 U1042 ( .A1(KEYINPUT38), .A2(n1072), .ZN(n1323) );
AND2_X1 U1043 ( .A1(n1324), .A2(n1259), .ZN(n1072) );
XOR2_X1 U1044 ( .A(KEYINPUT60), .B(n1134), .Z(n1324) );
XNOR2_X1 U1045 ( .A(n1325), .B(n1326), .ZN(n1134) );
XOR2_X1 U1046 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1047 ( .A(G122), .B(G104), .Z(n1328) );
XOR2_X1 U1048 ( .A(G146), .B(G131), .Z(n1327) );
XOR2_X1 U1049 ( .A(n1329), .B(n1330), .Z(n1325) );
XOR2_X1 U1050 ( .A(n1331), .B(n1332), .Z(n1330) );
AND2_X1 U1051 ( .A1(n1315), .A2(G214), .ZN(n1332) );
NOR2_X1 U1052 ( .A1(G953), .A2(G237), .ZN(n1315) );
NOR2_X1 U1053 ( .A1(KEYINPUT31), .A2(n1298), .ZN(n1331) );
INV_X1 U1054 ( .A(n1099), .ZN(n1298) );
XOR2_X1 U1055 ( .A(G125), .B(G140), .Z(n1099) );
XNOR2_X1 U1056 ( .A(n1333), .B(n1334), .ZN(n1329) );
NAND2_X1 U1057 ( .A1(KEYINPUT45), .A2(n1285), .ZN(n1334) );
NAND2_X1 U1058 ( .A1(KEYINPUT42), .A2(n1249), .ZN(n1333) );
INV_X1 U1059 ( .A(G113), .ZN(n1249) );
INV_X1 U1060 ( .A(n1246), .ZN(n1242) );
XNOR2_X1 U1061 ( .A(n1077), .B(G478), .ZN(n1246) );
AND2_X1 U1062 ( .A1(n1335), .A2(n1259), .ZN(n1077) );
INV_X1 U1063 ( .A(G902), .ZN(n1259) );
XOR2_X1 U1064 ( .A(KEYINPUT3), .B(n1336), .Z(n1335) );
INV_X1 U1065 ( .A(n1130), .ZN(n1336) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1130) );
XOR2_X1 U1067 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1068 ( .A(n1341), .B(G116), .Z(n1340) );
NAND2_X1 U1069 ( .A1(KEYINPUT8), .A2(n1230), .ZN(n1341) );
INV_X1 U1070 ( .A(G134), .ZN(n1230) );
XOR2_X1 U1071 ( .A(n1342), .B(KEYINPUT56), .Z(n1339) );
INV_X1 U1072 ( .A(G122), .ZN(n1342) );
XNOR2_X1 U1073 ( .A(n1317), .B(n1343), .ZN(n1337) );
XOR2_X1 U1074 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1075 ( .A1(G217), .A2(n1299), .ZN(n1345) );
AND2_X1 U1076 ( .A1(G234), .A2(n1082), .ZN(n1299) );
INV_X1 U1077 ( .A(G953), .ZN(n1082) );
NAND2_X1 U1078 ( .A1(KEYINPUT53), .A2(n1021), .ZN(n1344) );
INV_X1 U1079 ( .A(G107), .ZN(n1021) );
XOR2_X1 U1080 ( .A(G128), .B(n1285), .Z(n1317) );
XOR2_X1 U1081 ( .A(G143), .B(KEYINPUT14), .Z(n1285) );
INV_X1 U1082 ( .A(G110), .ZN(n1168) );
endmodule


