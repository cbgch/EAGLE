//Key = 1010100000000111001011100110100110101001000101001010001011001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358;

XNOR2_X1 U735 ( .A(n1028), .B(n1029), .ZN(G9) );
AND2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1034), .A2(n1035), .A3(G953), .A4(n1036), .ZN(n1033) );
NOR4_X1 U739 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1035) );
AND3_X1 U740 ( .A1(KEYINPUT19), .A2(n1041), .A3(n1042), .ZN(n1038) );
NOR2_X1 U741 ( .A1(KEYINPUT19), .A2(n1043), .ZN(n1037) );
NOR2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U743 ( .A1(n1046), .A2(n1041), .ZN(n1044) );
NAND3_X1 U744 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1034) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1050), .ZN(n1048) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U747 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1045), .ZN(n1054) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U752 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND3_X1 U753 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1060) );
OR2_X1 U754 ( .A1(n1062), .A2(n1064), .ZN(n1066) );
OR3_X1 U755 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1065) );
NAND2_X1 U756 ( .A1(n1042), .A2(n1071), .ZN(n1051) );
INV_X1 U757 ( .A(n1045), .ZN(n1042) );
NAND4_X1 U758 ( .A1(n1058), .A2(n1064), .A3(n1067), .A4(n1062), .ZN(n1045) );
INV_X1 U759 ( .A(n1072), .ZN(n1058) );
NOR3_X1 U760 ( .A1(n1036), .A2(G953), .A3(G952), .ZN(n1032) );
AND4_X1 U761 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1036) );
NOR4_X1 U762 ( .A1(n1070), .A2(n1040), .A3(n1077), .A4(n1078), .ZN(n1076) );
XOR2_X1 U763 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U764 ( .A(G472), .B(KEYINPUT3), .ZN(n1080) );
XNOR2_X1 U765 ( .A(KEYINPUT51), .B(n1081), .ZN(n1077) );
NOR3_X1 U766 ( .A1(n1082), .A2(n1063), .A3(n1039), .ZN(n1075) );
INV_X1 U767 ( .A(n1083), .ZN(n1082) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U770 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U771 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U772 ( .A(n1092), .B(KEYINPUT0), .ZN(n1086) );
INV_X1 U773 ( .A(n1093), .ZN(n1092) );
NAND2_X1 U774 ( .A1(n1094), .A2(n1095), .ZN(n1084) );
NAND2_X1 U775 ( .A1(n1088), .A2(n1091), .ZN(n1094) );
INV_X1 U776 ( .A(KEYINPUT29), .ZN(n1091) );
XNOR2_X1 U777 ( .A(KEYINPUT35), .B(n1093), .ZN(n1088) );
XOR2_X1 U778 ( .A(n1096), .B(n1097), .Z(G72) );
NOR2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1098) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(n1100) );
NOR2_X1 U784 ( .A1(n1047), .A2(G953), .ZN(n1105) );
OR2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U787 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1109), .B(n1110), .Z(n1106) );
XNOR2_X1 U789 ( .A(n1111), .B(n1112), .ZN(n1110) );
INV_X1 U790 ( .A(n1113), .ZN(n1112) );
XOR2_X1 U791 ( .A(KEYINPUT57), .B(n1114), .Z(n1109) );
NOR3_X1 U792 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
AND2_X1 U793 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1117) );
NOR2_X1 U794 ( .A1(KEYINPUT16), .A2(n1118), .ZN(n1116) );
INV_X1 U795 ( .A(KEYINPUT56), .ZN(n1102) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U798 ( .A1(G953), .A2(n1123), .ZN(n1122) );
NAND2_X1 U799 ( .A1(G898), .A2(G224), .ZN(n1123) );
NAND3_X1 U800 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1121) );
NAND2_X1 U801 ( .A1(G953), .A2(n1127), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
XOR2_X1 U803 ( .A(KEYINPUT37), .B(n1130), .Z(n1128) );
NAND2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(n1124) );
XNOR2_X1 U805 ( .A(n1130), .B(KEYINPUT5), .ZN(n1131) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1130) );
NOR2_X1 U807 ( .A1(n1049), .A2(G953), .ZN(n1119) );
NOR2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U810 ( .A(n1139), .B(KEYINPUT60), .Z(n1138) );
OR2_X1 U811 ( .A1(n1140), .A2(n1093), .ZN(n1139) );
NAND2_X1 U812 ( .A1(KEYINPUT34), .A2(n1141), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1142), .ZN(G63) );
XNOR2_X1 U814 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U815 ( .A1(n1145), .A2(n1140), .ZN(n1144) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1146), .ZN(G60) );
XOR2_X1 U817 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1140), .ZN(n1148) );
XOR2_X1 U819 ( .A(G104), .B(n1150), .Z(G6) );
NOR2_X1 U820 ( .A1(n1135), .A2(n1151), .ZN(G57) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U823 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U824 ( .A1(n1158), .A2(n1140), .ZN(n1157) );
INV_X1 U825 ( .A(G472), .ZN(n1158) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
NOR2_X1 U827 ( .A1(n1135), .A2(n1161), .ZN(G54) );
XOR2_X1 U828 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U829 ( .A(n1164), .B(n1113), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1165), .A2(KEYINPUT36), .ZN(n1164) );
XOR2_X1 U831 ( .A(n1166), .B(n1111), .Z(n1165) );
XOR2_X1 U832 ( .A(n1167), .B(n1168), .Z(n1162) );
NOR2_X1 U833 ( .A1(n1169), .A2(n1140), .ZN(n1168) );
NOR3_X1 U834 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1167) );
AND2_X1 U835 ( .A1(n1173), .A2(KEYINPUT1), .ZN(n1172) );
AND3_X1 U836 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1171) );
INV_X1 U837 ( .A(KEYINPUT1), .ZN(n1174) );
NOR2_X1 U838 ( .A1(n1176), .A2(n1175), .ZN(n1170) );
XNOR2_X1 U839 ( .A(G110), .B(n1177), .ZN(n1175) );
NOR2_X1 U840 ( .A1(KEYINPUT44), .A2(n1173), .ZN(n1176) );
NOR2_X1 U841 ( .A1(n1135), .A2(n1178), .ZN(G51) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U843 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U844 ( .A1(n1183), .A2(n1140), .ZN(n1182) );
NAND2_X1 U845 ( .A1(G902), .A2(n1184), .ZN(n1140) );
NAND2_X1 U846 ( .A1(n1049), .A2(n1047), .ZN(n1184) );
AND2_X1 U847 ( .A1(n1185), .A2(n1186), .ZN(n1047) );
NOR4_X1 U848 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
AND4_X1 U849 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1185) );
AND4_X1 U850 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1049) );
NOR4_X1 U851 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1150), .ZN(n1198) );
AND3_X1 U852 ( .A1(n1031), .A2(n1202), .A3(n1069), .ZN(n1150) );
AND2_X1 U853 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
NAND2_X1 U854 ( .A1(n1205), .A2(n1030), .ZN(n1195) );
AND2_X1 U855 ( .A1(n1202), .A2(n1068), .ZN(n1030) );
XNOR2_X1 U856 ( .A(n1031), .B(KEYINPUT22), .ZN(n1205) );
NOR2_X1 U857 ( .A1(n1206), .A2(n1207), .ZN(n1181) );
XOR2_X1 U858 ( .A(KEYINPUT8), .B(n1208), .Z(n1207) );
NOR2_X1 U859 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
AND2_X1 U860 ( .A1(n1210), .A2(n1209), .ZN(n1206) );
XNOR2_X1 U861 ( .A(n1211), .B(n1212), .ZN(n1210) );
NOR2_X1 U862 ( .A1(G125), .A2(KEYINPUT41), .ZN(n1212) );
NOR2_X1 U863 ( .A1(n1099), .A2(G952), .ZN(n1135) );
XNOR2_X1 U864 ( .A(n1213), .B(n1214), .ZN(G48) );
NAND2_X1 U865 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
NAND2_X1 U866 ( .A1(n1190), .A2(n1217), .ZN(n1216) );
INV_X1 U867 ( .A(KEYINPUT27), .ZN(n1217) );
AND4_X1 U868 ( .A1(n1218), .A2(n1069), .A3(n1071), .A4(n1219), .ZN(n1190) );
NAND4_X1 U869 ( .A1(n1220), .A2(n1069), .A3(n1221), .A4(KEYINPUT27), .ZN(n1215) );
AND3_X1 U870 ( .A1(n1222), .A2(n1070), .A3(n1219), .ZN(n1221) );
INV_X1 U871 ( .A(n1223), .ZN(n1220) );
XOR2_X1 U872 ( .A(G143), .B(n1224), .Z(G45) );
NOR3_X1 U873 ( .A1(KEYINPUT11), .A2(n1225), .A3(n1226), .ZN(n1224) );
NOR2_X1 U874 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
INV_X1 U875 ( .A(KEYINPUT55), .ZN(n1228) );
NOR2_X1 U876 ( .A1(n1071), .A2(n1229), .ZN(n1227) );
NOR2_X1 U877 ( .A1(KEYINPUT55), .A2(n1189), .ZN(n1225) );
NOR2_X1 U878 ( .A1(n1229), .A2(n1230), .ZN(n1189) );
NAND4_X1 U879 ( .A1(n1218), .A2(n1046), .A3(n1231), .A4(n1232), .ZN(n1229) );
XOR2_X1 U880 ( .A(n1188), .B(n1233), .Z(G42) );
NOR2_X1 U881 ( .A1(KEYINPUT47), .A2(n1177), .ZN(n1233) );
AND3_X1 U882 ( .A1(n1069), .A2(n1041), .A3(n1234), .ZN(n1188) );
XOR2_X1 U883 ( .A(G137), .B(n1187), .Z(G39) );
AND3_X1 U884 ( .A1(n1064), .A2(n1219), .A3(n1234), .ZN(n1187) );
XNOR2_X1 U885 ( .A(G134), .B(n1193), .ZN(G36) );
NAND3_X1 U886 ( .A1(n1046), .A2(n1068), .A3(n1234), .ZN(n1193) );
XOR2_X1 U887 ( .A(G131), .B(n1235), .Z(G33) );
NOR2_X1 U888 ( .A1(KEYINPUT24), .A2(n1194), .ZN(n1235) );
NAND3_X1 U889 ( .A1(n1069), .A2(n1046), .A3(n1234), .ZN(n1194) );
AND3_X1 U890 ( .A1(n1055), .A2(n1057), .A3(n1218), .ZN(n1234) );
XNOR2_X1 U891 ( .A(G128), .B(n1236), .ZN(G30) );
NOR2_X1 U892 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U893 ( .A1(n1239), .A2(n1192), .ZN(n1238) );
NAND4_X1 U894 ( .A1(n1218), .A2(n1068), .A3(n1071), .A4(n1219), .ZN(n1192) );
INV_X1 U895 ( .A(KEYINPUT28), .ZN(n1239) );
NOR2_X1 U896 ( .A1(KEYINPUT28), .A2(n1240), .ZN(n1237) );
NAND4_X1 U897 ( .A1(n1218), .A2(n1068), .A3(n1219), .A4(n1230), .ZN(n1240) );
INV_X1 U898 ( .A(n1071), .ZN(n1230) );
AND3_X1 U899 ( .A1(n1070), .A2(n1223), .A3(n1067), .ZN(n1218) );
XOR2_X1 U900 ( .A(G101), .B(n1241), .Z(G3) );
NOR2_X1 U901 ( .A1(KEYINPUT12), .A2(n1196), .ZN(n1241) );
NAND3_X1 U902 ( .A1(n1064), .A2(n1202), .A3(n1046), .ZN(n1196) );
XNOR2_X1 U903 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U904 ( .A1(n1041), .A2(n1223), .A3(n1222), .A4(n1242), .ZN(n1191) );
NOR2_X1 U905 ( .A1(n1243), .A2(n1070), .ZN(n1242) );
NAND2_X1 U906 ( .A1(n1072), .A2(n1244), .ZN(n1223) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1108), .ZN(n1244) );
INV_X1 U908 ( .A(G900), .ZN(n1108) );
XOR2_X1 U909 ( .A(n1204), .B(n1246), .Z(G24) );
XOR2_X1 U910 ( .A(KEYINPUT2), .B(G122), .Z(n1246) );
NAND4_X1 U911 ( .A1(n1247), .A2(n1031), .A3(n1231), .A4(n1232), .ZN(n1204) );
XNOR2_X1 U912 ( .A(G119), .B(n1203), .ZN(G21) );
NAND3_X1 U913 ( .A1(n1064), .A2(n1219), .A3(n1247), .ZN(n1203) );
NAND2_X1 U914 ( .A1(n1248), .A2(n1249), .ZN(n1219) );
NAND2_X1 U915 ( .A1(n1046), .A2(n1250), .ZN(n1249) );
NAND3_X1 U916 ( .A1(n1251), .A2(n1252), .A3(KEYINPUT50), .ZN(n1248) );
XOR2_X1 U917 ( .A(G116), .B(n1201), .Z(G18) );
AND3_X1 U918 ( .A1(n1046), .A2(n1068), .A3(n1247), .ZN(n1201) );
NOR2_X1 U919 ( .A1(n1232), .A2(n1253), .ZN(n1068) );
XOR2_X1 U920 ( .A(n1200), .B(n1254), .Z(G15) );
NOR2_X1 U921 ( .A1(KEYINPUT10), .A2(n1255), .ZN(n1254) );
AND3_X1 U922 ( .A1(n1069), .A2(n1046), .A3(n1247), .ZN(n1200) );
AND3_X1 U923 ( .A1(n1222), .A2(n1256), .A3(n1062), .ZN(n1247) );
INV_X1 U924 ( .A(n1070), .ZN(n1062) );
AND2_X1 U925 ( .A1(n1257), .A2(n1251), .ZN(n1046) );
INV_X1 U926 ( .A(n1243), .ZN(n1069) );
NAND2_X1 U927 ( .A1(n1253), .A2(n1232), .ZN(n1243) );
INV_X1 U928 ( .A(n1231), .ZN(n1253) );
XNOR2_X1 U929 ( .A(G110), .B(n1258), .ZN(G12) );
NAND2_X1 U930 ( .A1(KEYINPUT15), .A2(n1199), .ZN(n1258) );
AND3_X1 U931 ( .A1(n1202), .A2(n1041), .A3(n1064), .ZN(n1199) );
NOR2_X1 U932 ( .A1(n1231), .A2(n1232), .ZN(n1064) );
NAND2_X1 U933 ( .A1(n1081), .A2(n1083), .ZN(n1232) );
NAND2_X1 U934 ( .A1(G475), .A2(n1259), .ZN(n1083) );
NAND2_X1 U935 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U936 ( .A1(n1261), .A2(n1149), .A3(n1260), .ZN(n1081) );
XOR2_X1 U937 ( .A(n1147), .B(KEYINPUT39), .Z(n1260) );
XOR2_X1 U938 ( .A(n1262), .B(n1263), .Z(n1147) );
XOR2_X1 U939 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U940 ( .A(n1255), .B(G104), .ZN(n1265) );
INV_X1 U941 ( .A(G113), .ZN(n1255) );
XNOR2_X1 U942 ( .A(n1214), .B(G131), .ZN(n1264) );
XOR2_X1 U943 ( .A(n1266), .B(n1267), .Z(n1262) );
XOR2_X1 U944 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR3_X1 U945 ( .A1(n1115), .A2(n1270), .A3(n1271), .ZN(n1269) );
NOR2_X1 U946 ( .A1(n1272), .A2(n1118), .ZN(n1271) );
INV_X1 U947 ( .A(KEYINPUT13), .ZN(n1272) );
NOR2_X1 U948 ( .A1(KEYINPUT13), .A2(n1273), .ZN(n1270) );
NOR2_X1 U949 ( .A1(KEYINPUT38), .A2(n1274), .ZN(n1268) );
XOR2_X1 U950 ( .A(G143), .B(n1275), .Z(n1274) );
NOR3_X1 U951 ( .A1(n1276), .A2(G237), .A3(n1277), .ZN(n1275) );
INV_X1 U952 ( .A(G214), .ZN(n1277) );
XNOR2_X1 U953 ( .A(KEYINPUT52), .B(n1099), .ZN(n1276) );
INV_X1 U954 ( .A(G475), .ZN(n1149) );
XNOR2_X1 U955 ( .A(n1073), .B(KEYINPUT63), .ZN(n1231) );
XNOR2_X1 U956 ( .A(n1278), .B(n1145), .ZN(n1073) );
INV_X1 U957 ( .A(G478), .ZN(n1145) );
NAND2_X1 U958 ( .A1(n1143), .A2(n1261), .ZN(n1278) );
XNOR2_X1 U959 ( .A(n1279), .B(n1280), .ZN(n1143) );
XOR2_X1 U960 ( .A(n1281), .B(n1266), .Z(n1280) );
NAND2_X1 U961 ( .A1(n1282), .A2(G217), .ZN(n1281) );
XOR2_X1 U962 ( .A(n1283), .B(n1284), .Z(n1279) );
NOR2_X1 U963 ( .A1(KEYINPUT6), .A2(n1285), .ZN(n1284) );
XOR2_X1 U964 ( .A(G128), .B(n1286), .Z(n1285) );
XOR2_X1 U965 ( .A(G143), .B(G134), .Z(n1286) );
XNOR2_X1 U966 ( .A(G107), .B(G116), .ZN(n1283) );
NAND2_X1 U967 ( .A1(n1287), .A2(n1288), .ZN(n1041) );
NAND2_X1 U968 ( .A1(n1031), .A2(n1250), .ZN(n1288) );
NOR2_X1 U969 ( .A1(n1252), .A2(n1251), .ZN(n1031) );
OR3_X1 U970 ( .A1(n1257), .A2(n1251), .A3(n1250), .ZN(n1287) );
INV_X1 U971 ( .A(KEYINPUT50), .ZN(n1250) );
XOR2_X1 U972 ( .A(G472), .B(n1289), .Z(n1251) );
NOR2_X1 U973 ( .A1(KEYINPUT42), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U974 ( .A(KEYINPUT31), .B(n1079), .ZN(n1290) );
NAND2_X1 U975 ( .A1(n1261), .A2(n1291), .ZN(n1079) );
NAND2_X1 U976 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U977 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U978 ( .A1(n1296), .A2(n1160), .ZN(n1295) );
XNOR2_X1 U979 ( .A(n1297), .B(n1154), .ZN(n1294) );
XOR2_X1 U980 ( .A(n1298), .B(KEYINPUT9), .Z(n1292) );
NAND3_X1 U981 ( .A1(n1296), .A2(n1160), .A3(n1299), .ZN(n1298) );
XOR2_X1 U982 ( .A(n1297), .B(n1154), .Z(n1299) );
XNOR2_X1 U983 ( .A(n1300), .B(n1113), .ZN(n1154) );
XOR2_X1 U984 ( .A(n1211), .B(KEYINPUT62), .Z(n1300) );
NAND2_X1 U985 ( .A1(KEYINPUT18), .A2(n1155), .ZN(n1297) );
XNOR2_X1 U986 ( .A(n1301), .B(n1302), .ZN(n1155) );
XNOR2_X1 U987 ( .A(G116), .B(KEYINPUT53), .ZN(n1301) );
NAND4_X1 U988 ( .A1(G210), .A2(G101), .A3(n1303), .A4(n1099), .ZN(n1160) );
XOR2_X1 U989 ( .A(KEYINPUT7), .B(n1159), .Z(n1296) );
OR2_X1 U990 ( .A1(G101), .A2(n1304), .ZN(n1159) );
AND3_X1 U991 ( .A1(n1303), .A2(n1099), .A3(G210), .ZN(n1304) );
INV_X1 U992 ( .A(n1252), .ZN(n1257) );
XOR2_X1 U993 ( .A(n1305), .B(n1093), .Z(n1252) );
NAND2_X1 U994 ( .A1(G217), .A2(n1306), .ZN(n1093) );
XNOR2_X1 U995 ( .A(KEYINPUT54), .B(n1307), .ZN(n1305) );
NOR2_X1 U996 ( .A1(n1090), .A2(KEYINPUT40), .ZN(n1307) );
INV_X1 U997 ( .A(n1095), .ZN(n1090) );
NAND2_X1 U998 ( .A1(n1141), .A2(n1261), .ZN(n1095) );
XNOR2_X1 U999 ( .A(n1308), .B(n1309), .ZN(n1141) );
XOR2_X1 U1000 ( .A(G137), .B(n1310), .Z(n1309) );
NOR2_X1 U1001 ( .A1(KEYINPUT46), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1002 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1003 ( .A(n1314), .B(n1315), .Z(n1313) );
NAND2_X1 U1004 ( .A1(n1316), .A2(n1118), .ZN(n1315) );
NAND2_X1 U1005 ( .A1(n1177), .A2(n1273), .ZN(n1118) );
INV_X1 U1006 ( .A(n1115), .ZN(n1316) );
NOR2_X1 U1007 ( .A1(n1177), .A2(n1273), .ZN(n1115) );
NAND2_X1 U1008 ( .A1(n1317), .A2(KEYINPUT21), .ZN(n1314) );
XNOR2_X1 U1009 ( .A(G119), .B(n1318), .ZN(n1317) );
XOR2_X1 U1010 ( .A(KEYINPUT45), .B(G128), .Z(n1318) );
XNOR2_X1 U1011 ( .A(G146), .B(G110), .ZN(n1312) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1282), .ZN(n1308) );
AND2_X1 U1013 ( .A1(G234), .A2(n1099), .ZN(n1282) );
AND3_X1 U1014 ( .A1(n1070), .A2(n1256), .A3(n1222), .ZN(n1202) );
AND2_X1 U1015 ( .A1(n1071), .A2(n1067), .ZN(n1222) );
XNOR2_X1 U1016 ( .A(n1063), .B(KEYINPUT33), .ZN(n1067) );
AND2_X1 U1017 ( .A1(G221), .A2(n1306), .ZN(n1063) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1319), .ZN(n1306) );
NOR2_X1 U1019 ( .A1(n1055), .A2(n1039), .ZN(n1071) );
INV_X1 U1020 ( .A(n1057), .ZN(n1039) );
NAND2_X1 U1021 ( .A1(n1320), .A2(G214), .ZN(n1057) );
XOR2_X1 U1022 ( .A(n1321), .B(KEYINPUT59), .Z(n1320) );
INV_X1 U1023 ( .A(n1040), .ZN(n1055) );
XOR2_X1 U1024 ( .A(n1322), .B(n1183), .Z(n1040) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1321), .ZN(n1183) );
NAND2_X1 U1026 ( .A1(n1319), .A2(n1303), .ZN(n1321) );
INV_X1 U1027 ( .A(G237), .ZN(n1303) );
NAND2_X1 U1028 ( .A1(n1323), .A2(n1261), .ZN(n1322) );
XOR2_X1 U1029 ( .A(n1324), .B(n1179), .Z(n1323) );
XNOR2_X1 U1030 ( .A(n1134), .B(n1325), .ZN(n1179) );
XNOR2_X1 U1031 ( .A(n1326), .B(n1129), .ZN(n1325) );
INV_X1 U1032 ( .A(n1132), .ZN(n1129) );
XOR2_X1 U1033 ( .A(n1327), .B(n1328), .Z(n1132) );
NOR2_X1 U1034 ( .A1(KEYINPUT49), .A2(n1329), .ZN(n1328) );
NOR2_X1 U1035 ( .A1(KEYINPUT23), .A2(n1133), .ZN(n1326) );
AND2_X1 U1036 ( .A1(n1330), .A2(n1331), .ZN(n1133) );
OR2_X1 U1037 ( .A1(n1302), .A2(G116), .ZN(n1331) );
NAND2_X1 U1038 ( .A1(n1332), .A2(G116), .ZN(n1330) );
XOR2_X1 U1039 ( .A(KEYINPUT30), .B(n1302), .Z(n1332) );
XOR2_X1 U1040 ( .A(G113), .B(G119), .Z(n1302) );
XNOR2_X1 U1041 ( .A(G110), .B(n1266), .ZN(n1134) );
XNOR2_X1 U1042 ( .A(G122), .B(KEYINPUT20), .ZN(n1266) );
NAND3_X1 U1043 ( .A1(n1333), .A2(n1334), .A3(KEYINPUT32), .ZN(n1324) );
NAND2_X1 U1044 ( .A1(n1209), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1045 ( .A(KEYINPUT4), .B(n1336), .Z(n1333) );
NOR2_X1 U1046 ( .A1(n1209), .A2(n1335), .ZN(n1336) );
XNOR2_X1 U1047 ( .A(n1211), .B(n1273), .ZN(n1335) );
INV_X1 U1048 ( .A(G125), .ZN(n1273) );
NAND2_X1 U1049 ( .A1(n1337), .A2(n1338), .ZN(n1211) );
NAND2_X1 U1050 ( .A1(G128), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1051 ( .A(n1340), .B(KEYINPUT58), .Z(n1337) );
OR2_X1 U1052 ( .A1(n1339), .A2(G128), .ZN(n1340) );
AND2_X1 U1053 ( .A1(G224), .A2(n1099), .ZN(n1209) );
NAND2_X1 U1054 ( .A1(n1072), .A2(n1341), .ZN(n1256) );
NAND4_X1 U1055 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1127), .ZN(n1341) );
INV_X1 U1056 ( .A(G898), .ZN(n1127) );
NAND3_X1 U1057 ( .A1(n1245), .A2(n1099), .A3(G952), .ZN(n1072) );
NAND2_X1 U1058 ( .A1(G237), .A2(G234), .ZN(n1245) );
XOR2_X1 U1059 ( .A(n1342), .B(n1169), .Z(n1070) );
INV_X1 U1060 ( .A(G469), .ZN(n1169) );
NAND2_X1 U1061 ( .A1(n1343), .A2(n1261), .ZN(n1342) );
XNOR2_X1 U1062 ( .A(n1319), .B(KEYINPUT25), .ZN(n1261) );
INV_X1 U1063 ( .A(G902), .ZN(n1319) );
XOR2_X1 U1064 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1065 ( .A(n1166), .B(n1113), .ZN(n1345) );
XOR2_X1 U1066 ( .A(G131), .B(n1346), .Z(n1113) );
XOR2_X1 U1067 ( .A(G137), .B(G134), .Z(n1346) );
XOR2_X1 U1068 ( .A(n1329), .B(n1347), .Z(n1166) );
XOR2_X1 U1069 ( .A(KEYINPUT43), .B(n1327), .Z(n1347) );
XNOR2_X1 U1070 ( .A(G104), .B(n1028), .ZN(n1327) );
INV_X1 U1071 ( .A(G107), .ZN(n1028) );
XNOR2_X1 U1072 ( .A(G101), .B(KEYINPUT61), .ZN(n1329) );
XOR2_X1 U1073 ( .A(n1348), .B(n1349), .Z(n1344) );
XNOR2_X1 U1074 ( .A(n1350), .B(n1173), .ZN(n1349) );
NAND2_X1 U1075 ( .A1(G227), .A2(n1099), .ZN(n1173) );
INV_X1 U1076 ( .A(G953), .ZN(n1099) );
NAND2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND4_X1 U1078 ( .A1(KEYINPUT14), .A2(n1353), .A3(n1177), .A4(n1354), .ZN(n1352) );
INV_X1 U1079 ( .A(KEYINPUT17), .ZN(n1354) );
NAND2_X1 U1080 ( .A1(n1355), .A2(n1356), .ZN(n1351) );
NAND2_X1 U1081 ( .A1(n1357), .A2(n1177), .ZN(n1356) );
INV_X1 U1082 ( .A(G140), .ZN(n1177) );
NAND2_X1 U1083 ( .A1(KEYINPUT17), .A2(G110), .ZN(n1357) );
NAND2_X1 U1084 ( .A1(KEYINPUT14), .A2(n1353), .ZN(n1355) );
INV_X1 U1085 ( .A(G110), .ZN(n1353) );
NAND2_X1 U1086 ( .A1(KEYINPUT48), .A2(n1111), .ZN(n1348) );
XNOR2_X1 U1087 ( .A(n1358), .B(G128), .ZN(n1111) );
NAND2_X1 U1088 ( .A1(KEYINPUT26), .A2(n1339), .ZN(n1358) );
XNOR2_X1 U1089 ( .A(G143), .B(n1214), .ZN(n1339) );
INV_X1 U1090 ( .A(G146), .ZN(n1214) );
endmodule


