//Key = 0011001100011110110101101001011010010001111110100100110110100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370;

XNOR2_X1 U752 ( .A(G107), .B(n1037), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR2_X1 U754 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND4_X1 U755 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NAND4_X1 U756 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
NOR2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND3_X1 U758 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NAND3_X1 U760 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1066), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
OR3_X1 U766 ( .A1(n1069), .A2(n1051), .A3(n1047), .ZN(n1068) );
INV_X1 U767 ( .A(KEYINPUT19), .ZN(n1047) );
NAND2_X1 U768 ( .A1(n1059), .A2(n1070), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1040) );
NAND3_X1 U771 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1074) );
XNOR2_X1 U772 ( .A(n1080), .B(KEYINPUT2), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1073) );
NOR2_X1 U774 ( .A1(n1050), .A2(n1082), .ZN(n1080) );
NAND3_X1 U775 ( .A1(n1062), .A2(n1057), .A3(n1052), .ZN(n1050) );
INV_X1 U776 ( .A(n1083), .ZN(n1052) );
NOR3_X1 U777 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1038) );
INV_X1 U778 ( .A(n1075), .ZN(n1084) );
NAND4_X1 U779 ( .A1(n1085), .A2(n1059), .A3(n1086), .A4(n1087), .ZN(n1075) );
NOR4_X1 U780 ( .A1(n1077), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1087) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
INV_X1 U782 ( .A(n1093), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1086) );
XNOR2_X1 U784 ( .A(G475), .B(n1096), .ZN(n1085) );
XOR2_X1 U785 ( .A(n1097), .B(n1098), .Z(G72) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U787 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1101) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NAND2_X1 U790 ( .A1(G953), .A2(n1104), .ZN(n1103) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(n1102) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(n1106) );
XNOR2_X1 U793 ( .A(n1109), .B(n1110), .ZN(n1105) );
NAND2_X1 U794 ( .A1(KEYINPUT42), .A2(n1111), .ZN(n1109) );
NOR2_X1 U795 ( .A1(n1043), .A2(G953), .ZN(n1097) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U798 ( .A1(n1042), .A2(G953), .ZN(n1115) );
NAND3_X1 U799 ( .A1(KEYINPUT58), .A2(n1116), .A3(n1117), .ZN(n1114) );
XOR2_X1 U800 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U801 ( .A(n1120), .B(n1121), .Z(n1118) );
NAND2_X1 U802 ( .A1(KEYINPUT16), .A2(n1122), .ZN(n1120) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1116) );
XNOR2_X1 U804 ( .A(G953), .B(KEYINPUT14), .ZN(n1123) );
NAND2_X1 U805 ( .A1(G953), .A2(n1125), .ZN(n1112) );
NAND2_X1 U806 ( .A1(G898), .A2(G224), .ZN(n1125) );
NOR2_X1 U807 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U808 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U809 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
XNOR2_X1 U810 ( .A(n1132), .B(KEYINPUT12), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(G63) );
XNOR2_X1 U812 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1131), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1132), .A2(n1137), .ZN(G60) );
NOR3_X1 U815 ( .A1(n1096), .A2(n1138), .A3(n1139), .ZN(n1137) );
NOR3_X1 U816 ( .A1(n1140), .A2(n1141), .A3(n1131), .ZN(n1139) );
INV_X1 U817 ( .A(n1142), .ZN(n1140) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1142), .ZN(n1138) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1141), .ZN(n1143) );
INV_X1 U820 ( .A(G475), .ZN(n1141) );
NOR2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U822 ( .A(G104), .B(n1147), .Z(G6) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U824 ( .A1(n1132), .A2(n1150), .ZN(G57) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U826 ( .A(n1153), .B(n1154), .ZN(n1152) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1151) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1131), .ZN(n1156) );
NAND2_X1 U829 ( .A1(KEYINPUT24), .A2(n1158), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n1132), .A2(n1159), .ZN(G54) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U832 ( .A1(n1162), .A2(KEYINPUT20), .ZN(n1161) );
NOR2_X1 U833 ( .A1(n1163), .A2(n1131), .ZN(n1162) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NAND3_X1 U835 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
INV_X1 U836 ( .A(n1169), .ZN(n1168) );
XOR2_X1 U837 ( .A(n1170), .B(KEYINPUT37), .Z(n1164) );
NAND2_X1 U838 ( .A1(n1169), .A2(n1171), .ZN(n1170) );
NAND2_X1 U839 ( .A1(n1166), .A2(n1167), .ZN(n1171) );
NAND2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1167) );
XOR2_X1 U841 ( .A(n1108), .B(n1174), .Z(n1172) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1166) );
INV_X1 U843 ( .A(n1173), .ZN(n1176) );
XNOR2_X1 U844 ( .A(n1174), .B(n1108), .ZN(n1175) );
XNOR2_X1 U845 ( .A(n1177), .B(n1178), .ZN(n1169) );
XNOR2_X1 U846 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U847 ( .A1(n1132), .A2(n1181), .ZN(G51) );
XOR2_X1 U848 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR2_X1 U849 ( .A1(n1184), .A2(n1131), .ZN(n1183) );
NAND2_X1 U850 ( .A1(G902), .A2(n1185), .ZN(n1131) );
NAND2_X1 U851 ( .A1(n1042), .A2(n1043), .ZN(n1185) );
INV_X1 U852 ( .A(n1145), .ZN(n1043) );
NAND4_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1145) );
NOR4_X1 U854 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
NOR2_X1 U855 ( .A1(KEYINPUT23), .A2(n1194), .ZN(n1193) );
NOR4_X1 U856 ( .A1(n1195), .A2(n1196), .A3(n1061), .A4(n1197), .ZN(n1190) );
XNOR2_X1 U857 ( .A(n1198), .B(KEYINPUT34), .ZN(n1195) );
NOR2_X1 U858 ( .A1(n1199), .A2(n1200), .ZN(n1188) );
NAND3_X1 U859 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1186) );
NAND2_X1 U860 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
NAND4_X1 U861 ( .A1(KEYINPUT23), .A2(n1059), .A3(n1206), .A4(n1196), .ZN(n1205) );
INV_X1 U862 ( .A(n1146), .ZN(n1042) );
NAND4_X1 U863 ( .A1(n1207), .A2(n1037), .A3(n1208), .A4(n1209), .ZN(n1146) );
NOR4_X1 U864 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
INV_X1 U865 ( .A(n1214), .ZN(n1213) );
NOR2_X1 U866 ( .A1(n1215), .A2(n1216), .ZN(n1208) );
NOR3_X1 U867 ( .A1(n1149), .A2(n1217), .A3(n1218), .ZN(n1216) );
NOR2_X1 U868 ( .A1(KEYINPUT46), .A2(n1219), .ZN(n1218) );
NOR3_X1 U869 ( .A1(n1220), .A2(n1196), .A3(n1067), .ZN(n1219) );
AND2_X1 U870 ( .A1(n1148), .A2(KEYINPUT46), .ZN(n1217) );
INV_X1 U871 ( .A(n1221), .ZN(n1148) );
NAND2_X1 U872 ( .A1(n1203), .A2(n1057), .ZN(n1149) );
INV_X1 U873 ( .A(n1222), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1221), .A2(n1057), .A3(n1223), .ZN(n1037) );
XOR2_X1 U875 ( .A(n1092), .B(KEYINPUT50), .Z(n1184) );
NOR2_X1 U876 ( .A1(n1224), .A2(n1225), .ZN(n1182) );
XOR2_X1 U877 ( .A(KEYINPUT1), .B(n1226), .Z(n1225) );
AND2_X1 U878 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U879 ( .A1(n1227), .A2(n1228), .ZN(n1224) );
XNOR2_X1 U880 ( .A(n1229), .B(n1230), .ZN(n1228) );
XOR2_X1 U881 ( .A(n1231), .B(n1232), .Z(n1229) );
NOR2_X1 U882 ( .A1(KEYINPUT9), .A2(n1233), .ZN(n1232) );
NOR2_X1 U883 ( .A1(n1076), .A2(G952), .ZN(n1132) );
XNOR2_X1 U884 ( .A(G146), .B(n1187), .ZN(G48) );
NAND4_X1 U885 ( .A1(n1234), .A2(n1203), .A3(n1198), .A4(n1081), .ZN(n1187) );
XNOR2_X1 U886 ( .A(n1235), .B(n1192), .ZN(G45) );
AND4_X1 U887 ( .A1(n1236), .A2(n1095), .A3(n1237), .A4(n1238), .ZN(n1192) );
NOR2_X1 U888 ( .A1(n1196), .A2(n1197), .ZN(n1238) );
XNOR2_X1 U889 ( .A(n1179), .B(n1239), .ZN(G42) );
NOR4_X1 U890 ( .A1(KEYINPUT54), .A2(n1072), .A3(n1060), .A4(n1204), .ZN(n1239) );
INV_X1 U891 ( .A(n1201), .ZN(n1072) );
XOR2_X1 U892 ( .A(n1191), .B(n1240), .Z(G39) );
XNOR2_X1 U893 ( .A(KEYINPUT26), .B(n1110), .ZN(n1240) );
AND3_X1 U894 ( .A1(n1198), .A2(n1062), .A3(n1241), .ZN(n1191) );
NAND2_X1 U895 ( .A1(n1242), .A2(n1243), .ZN(G36) );
NAND2_X1 U896 ( .A1(n1200), .A2(n1244), .ZN(n1243) );
NAND2_X1 U897 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U898 ( .A1(KEYINPUT38), .A2(n1247), .ZN(n1246) );
XOR2_X1 U899 ( .A(n1248), .B(KEYINPUT8), .Z(n1245) );
OR3_X1 U900 ( .A1(n1249), .A2(KEYINPUT38), .A3(n1200), .ZN(n1242) );
NOR3_X1 U901 ( .A1(n1061), .A2(n1071), .A3(n1204), .ZN(n1200) );
INV_X1 U902 ( .A(n1223), .ZN(n1061) );
INV_X1 U903 ( .A(n1247), .ZN(n1249) );
XNOR2_X1 U904 ( .A(n1248), .B(KEYINPUT3), .ZN(n1247) );
XNOR2_X1 U905 ( .A(G134), .B(KEYINPUT7), .ZN(n1248) );
XOR2_X1 U906 ( .A(n1250), .B(n1199), .Z(G33) );
NOR3_X1 U907 ( .A1(n1060), .A2(n1071), .A3(n1204), .ZN(n1199) );
INV_X1 U908 ( .A(n1241), .ZN(n1204) );
NOR2_X1 U909 ( .A1(n1049), .A2(n1197), .ZN(n1241) );
INV_X1 U910 ( .A(n1234), .ZN(n1197) );
INV_X1 U911 ( .A(n1054), .ZN(n1049) );
NOR2_X1 U912 ( .A1(n1251), .A2(n1077), .ZN(n1054) );
INV_X1 U913 ( .A(n1237), .ZN(n1071) );
NAND2_X1 U914 ( .A1(KEYINPUT49), .A2(n1252), .ZN(n1250) );
INV_X1 U915 ( .A(G131), .ZN(n1252) );
XNOR2_X1 U916 ( .A(G128), .B(n1253), .ZN(G30) );
NAND2_X1 U917 ( .A1(n1254), .A2(n1081), .ZN(n1253) );
XOR2_X1 U918 ( .A(n1255), .B(KEYINPUT63), .Z(n1254) );
NAND3_X1 U919 ( .A1(n1198), .A2(n1223), .A3(n1234), .ZN(n1255) );
NOR2_X1 U920 ( .A1(n1067), .A2(n1256), .ZN(n1234) );
XNOR2_X1 U921 ( .A(G101), .B(n1222), .ZN(G3) );
NAND3_X1 U922 ( .A1(n1221), .A2(n1237), .A3(n1062), .ZN(n1222) );
XOR2_X1 U923 ( .A(n1194), .B(n1257), .Z(G27) );
NAND2_X1 U924 ( .A1(KEYINPUT43), .A2(G125), .ZN(n1257) );
NAND4_X1 U925 ( .A1(n1203), .A2(n1059), .A3(n1258), .A4(n1201), .ZN(n1194) );
NOR2_X1 U926 ( .A1(n1256), .A2(n1196), .ZN(n1258) );
INV_X1 U927 ( .A(n1206), .ZN(n1256) );
NAND2_X1 U928 ( .A1(n1083), .A2(n1259), .ZN(n1206) );
NAND4_X1 U929 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1104), .ZN(n1259) );
INV_X1 U930 ( .A(G900), .ZN(n1104) );
INV_X1 U931 ( .A(n1082), .ZN(n1059) );
XNOR2_X1 U932 ( .A(G122), .B(n1207), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1261), .A2(n1236), .A3(n1057), .A4(n1095), .ZN(n1207) );
NAND2_X1 U934 ( .A1(n1262), .A2(n1263), .ZN(n1057) );
OR3_X1 U935 ( .A1(n1090), .A2(n1094), .A3(KEYINPUT45), .ZN(n1263) );
NAND2_X1 U936 ( .A1(KEYINPUT45), .A2(n1201), .ZN(n1262) );
XOR2_X1 U937 ( .A(G119), .B(n1212), .Z(G21) );
AND3_X1 U938 ( .A1(n1198), .A2(n1062), .A3(n1261), .ZN(n1212) );
XOR2_X1 U939 ( .A(G116), .B(n1264), .Z(G18) );
NOR2_X1 U940 ( .A1(KEYINPUT0), .A2(n1214), .ZN(n1264) );
NAND3_X1 U941 ( .A1(n1223), .A2(n1237), .A3(n1261), .ZN(n1214) );
NOR2_X1 U942 ( .A1(n1265), .A2(n1266), .ZN(n1223) );
XOR2_X1 U943 ( .A(n1211), .B(n1267), .Z(G15) );
NOR2_X1 U944 ( .A1(KEYINPUT28), .A2(n1268), .ZN(n1267) );
AND3_X1 U945 ( .A1(n1261), .A2(n1237), .A3(n1203), .ZN(n1211) );
INV_X1 U946 ( .A(n1060), .ZN(n1203) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1236), .ZN(n1060) );
XNOR2_X1 U948 ( .A(n1266), .B(KEYINPUT41), .ZN(n1236) );
INV_X1 U949 ( .A(n1095), .ZN(n1265) );
NAND2_X1 U950 ( .A1(n1269), .A2(n1270), .ZN(n1237) );
NAND3_X1 U951 ( .A1(n1090), .A2(n1271), .A3(n1272), .ZN(n1270) );
INV_X1 U952 ( .A(KEYINPUT45), .ZN(n1272) );
NAND2_X1 U953 ( .A1(KEYINPUT45), .A2(n1198), .ZN(n1269) );
AND2_X1 U954 ( .A1(n1094), .A2(n1090), .ZN(n1198) );
NOR3_X1 U955 ( .A1(n1196), .A2(n1273), .A3(n1082), .ZN(n1261) );
NAND2_X1 U956 ( .A1(n1046), .A2(n1051), .ZN(n1082) );
INV_X1 U957 ( .A(n1069), .ZN(n1046) );
XOR2_X1 U958 ( .A(n1210), .B(n1274), .Z(G12) );
NOR2_X1 U959 ( .A1(KEYINPUT48), .A2(n1275), .ZN(n1274) );
INV_X1 U960 ( .A(G110), .ZN(n1275) );
AND3_X1 U961 ( .A1(n1221), .A2(n1201), .A3(n1062), .ZN(n1210) );
NOR2_X1 U962 ( .A1(n1095), .A2(n1266), .ZN(n1062) );
XNOR2_X1 U963 ( .A(n1096), .B(n1276), .ZN(n1266) );
NOR2_X1 U964 ( .A1(KEYINPUT18), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U965 ( .A(G475), .B(KEYINPUT62), .ZN(n1277) );
NOR2_X1 U966 ( .A1(n1142), .A2(G902), .ZN(n1096) );
XNOR2_X1 U967 ( .A(n1278), .B(n1279), .ZN(n1142) );
XOR2_X1 U968 ( .A(n1107), .B(n1280), .Z(n1279) );
XOR2_X1 U969 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR3_X1 U970 ( .A1(n1283), .A2(KEYINPUT51), .A3(n1284), .ZN(n1282) );
NOR2_X1 U971 ( .A1(G104), .A2(n1285), .ZN(n1284) );
XOR2_X1 U972 ( .A(n1286), .B(KEYINPUT29), .Z(n1283) );
NAND2_X1 U973 ( .A1(G104), .A2(n1285), .ZN(n1286) );
XNOR2_X1 U974 ( .A(n1268), .B(G122), .ZN(n1285) );
INV_X1 U975 ( .A(G113), .ZN(n1268) );
NAND2_X1 U976 ( .A1(G214), .A2(n1287), .ZN(n1281) );
XNOR2_X1 U977 ( .A(n1288), .B(n1233), .ZN(n1107) );
XNOR2_X1 U978 ( .A(G131), .B(G140), .ZN(n1288) );
XNOR2_X1 U979 ( .A(G143), .B(n1289), .ZN(n1278) );
XOR2_X1 U980 ( .A(KEYINPUT60), .B(G146), .Z(n1289) );
XOR2_X1 U981 ( .A(n1290), .B(n1136), .Z(n1095) );
INV_X1 U982 ( .A(G478), .ZN(n1136) );
NAND2_X1 U983 ( .A1(n1134), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U984 ( .A(n1292), .B(n1293), .ZN(n1134) );
XOR2_X1 U985 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U986 ( .A(n1296), .B(n1297), .Z(n1295) );
AND3_X1 U987 ( .A1(G234), .A2(n1076), .A3(G217), .ZN(n1297) );
NAND2_X1 U988 ( .A1(KEYINPUT21), .A2(n1111), .ZN(n1296) );
XNOR2_X1 U989 ( .A(G116), .B(G107), .ZN(n1294) );
XOR2_X1 U990 ( .A(n1298), .B(n1299), .Z(n1292) );
XNOR2_X1 U991 ( .A(KEYINPUT53), .B(n1235), .ZN(n1299) );
INV_X1 U992 ( .A(G143), .ZN(n1235) );
XNOR2_X1 U993 ( .A(G128), .B(G122), .ZN(n1298) );
NOR2_X1 U994 ( .A1(n1090), .A2(n1271), .ZN(n1201) );
INV_X1 U995 ( .A(n1094), .ZN(n1271) );
XOR2_X1 U996 ( .A(n1300), .B(n1130), .Z(n1094) );
NAND2_X1 U997 ( .A1(G217), .A2(n1301), .ZN(n1130) );
NAND2_X1 U998 ( .A1(n1302), .A2(n1291), .ZN(n1300) );
XOR2_X1 U999 ( .A(KEYINPUT6), .B(n1129), .Z(n1302) );
XNOR2_X1 U1000 ( .A(n1303), .B(n1304), .ZN(n1129) );
XOR2_X1 U1001 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1002 ( .A(n1307), .B(n1308), .Z(n1306) );
AND3_X1 U1003 ( .A1(G221), .A2(n1076), .A3(G234), .ZN(n1308) );
NAND2_X1 U1004 ( .A1(KEYINPUT55), .A2(n1177), .ZN(n1307) );
NAND2_X1 U1005 ( .A1(KEYINPUT30), .A2(n1309), .ZN(n1305) );
XNOR2_X1 U1006 ( .A(n1233), .B(n1310), .ZN(n1309) );
XNOR2_X1 U1007 ( .A(n1311), .B(KEYINPUT59), .ZN(n1310) );
NAND2_X1 U1008 ( .A1(KEYINPUT32), .A2(n1179), .ZN(n1311) );
INV_X1 U1009 ( .A(n1312), .ZN(n1233) );
XNOR2_X1 U1010 ( .A(n1313), .B(n1314), .ZN(n1303) );
XNOR2_X1 U1011 ( .A(n1315), .B(n1316), .ZN(n1314) );
NOR2_X1 U1012 ( .A1(KEYINPUT15), .A2(n1110), .ZN(n1316) );
NAND2_X1 U1013 ( .A1(KEYINPUT11), .A2(G119), .ZN(n1315) );
XOR2_X1 U1014 ( .A(n1317), .B(n1157), .Z(n1090) );
INV_X1 U1015 ( .A(G472), .ZN(n1157) );
NAND3_X1 U1016 ( .A1(n1318), .A2(n1291), .A3(n1319), .ZN(n1317) );
NAND3_X1 U1017 ( .A1(n1320), .A2(n1321), .A3(n1153), .ZN(n1319) );
XOR2_X1 U1018 ( .A(n1322), .B(n1323), .Z(n1320) );
NOR2_X1 U1019 ( .A1(n1154), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1020 ( .A1(n1325), .A2(n1326), .ZN(n1318) );
NAND2_X1 U1021 ( .A1(n1153), .A2(n1321), .ZN(n1326) );
INV_X1 U1022 ( .A(KEYINPUT4), .ZN(n1321) );
XNOR2_X1 U1023 ( .A(n1230), .B(n1173), .ZN(n1153) );
XOR2_X1 U1024 ( .A(n1327), .B(n1323), .Z(n1325) );
XNOR2_X1 U1025 ( .A(n1158), .B(n1328), .ZN(n1323) );
XOR2_X1 U1026 ( .A(KEYINPUT36), .B(KEYINPUT27), .Z(n1328) );
XNOR2_X1 U1027 ( .A(n1329), .B(n1330), .ZN(n1158) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1287), .ZN(n1329) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1287) );
NOR2_X1 U1030 ( .A1(n1122), .A2(n1324), .ZN(n1327) );
INV_X1 U1031 ( .A(KEYINPUT17), .ZN(n1324) );
NOR3_X1 U1032 ( .A1(n1196), .A2(n1273), .A3(n1067), .ZN(n1221) );
NAND2_X1 U1033 ( .A1(n1069), .A2(n1051), .ZN(n1067) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1301), .ZN(n1051) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1291), .ZN(n1301) );
XOR2_X1 U1036 ( .A(n1331), .B(n1163), .Z(n1069) );
INV_X1 U1037 ( .A(G469), .ZN(n1163) );
NAND2_X1 U1038 ( .A1(n1332), .A2(n1291), .ZN(n1331) );
XOR2_X1 U1039 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1040 ( .A(n1108), .B(n1335), .Z(n1334) );
XNOR2_X1 U1041 ( .A(n1336), .B(n1173), .ZN(n1335) );
XOR2_X1 U1042 ( .A(G131), .B(n1337), .Z(n1173) );
NOR2_X1 U1043 ( .A1(KEYINPUT10), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1044 ( .A(n1111), .B(n1339), .ZN(n1338) );
XNOR2_X1 U1045 ( .A(KEYINPUT44), .B(n1110), .ZN(n1339) );
INV_X1 U1046 ( .A(G137), .ZN(n1110) );
INV_X1 U1047 ( .A(G134), .ZN(n1111) );
NAND2_X1 U1048 ( .A1(KEYINPUT35), .A2(n1174), .ZN(n1336) );
XNOR2_X1 U1049 ( .A(n1340), .B(n1341), .ZN(n1174) );
NOR2_X1 U1050 ( .A1(KEYINPUT25), .A2(G104), .ZN(n1341) );
XNOR2_X1 U1051 ( .A(G101), .B(G107), .ZN(n1340) );
XOR2_X1 U1052 ( .A(n1230), .B(KEYINPUT22), .Z(n1108) );
XOR2_X1 U1053 ( .A(n1342), .B(n1343), .Z(n1333) );
XNOR2_X1 U1054 ( .A(KEYINPUT5), .B(n1179), .ZN(n1343) );
INV_X1 U1055 ( .A(G140), .ZN(n1179) );
XOR2_X1 U1056 ( .A(n1344), .B(n1180), .Z(n1342) );
AND2_X1 U1057 ( .A1(G227), .A2(n1076), .ZN(n1180) );
NAND2_X1 U1058 ( .A1(KEYINPUT39), .A2(n1177), .ZN(n1344) );
INV_X1 U1059 ( .A(n1220), .ZN(n1273) );
NAND2_X1 U1060 ( .A1(n1083), .A2(n1345), .ZN(n1220) );
NAND4_X1 U1061 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1124), .ZN(n1345) );
INV_X1 U1062 ( .A(G898), .ZN(n1124) );
NAND3_X1 U1063 ( .A1(n1260), .A2(n1076), .A3(G952), .ZN(n1083) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1260) );
INV_X1 U1065 ( .A(n1081), .ZN(n1196) );
NOR2_X1 U1066 ( .A1(n1077), .A2(n1078), .ZN(n1081) );
INV_X1 U1067 ( .A(n1251), .ZN(n1078) );
NAND2_X1 U1068 ( .A1(n1346), .A2(n1093), .ZN(n1251) );
NAND2_X1 U1069 ( .A1(n1091), .A2(n1092), .ZN(n1093) );
XOR2_X1 U1070 ( .A(n1347), .B(KEYINPUT57), .Z(n1346) );
OR2_X1 U1071 ( .A1(n1092), .A2(n1091), .ZN(n1347) );
AND2_X1 U1072 ( .A1(n1348), .A2(n1291), .ZN(n1091) );
XOR2_X1 U1073 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1074 ( .A(n1227), .B(n1231), .ZN(n1350) );
NAND2_X1 U1075 ( .A1(G224), .A2(n1076), .ZN(n1231) );
INV_X1 U1076 ( .A(G953), .ZN(n1076) );
NAND2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1227) );
OR2_X1 U1078 ( .A1(n1119), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1079 ( .A(n1354), .B(KEYINPUT33), .Z(n1351) );
NAND2_X1 U1080 ( .A1(n1353), .A2(n1119), .ZN(n1354) );
XNOR2_X1 U1081 ( .A(n1355), .B(G122), .ZN(n1119) );
NAND2_X1 U1082 ( .A1(KEYINPUT13), .A2(n1177), .ZN(n1355) );
XNOR2_X1 U1083 ( .A(G110), .B(KEYINPUT47), .ZN(n1177) );
XNOR2_X1 U1084 ( .A(n1121), .B(n1122), .ZN(n1353) );
INV_X1 U1085 ( .A(n1154), .ZN(n1122) );
XNOR2_X1 U1086 ( .A(n1356), .B(n1357), .ZN(n1154) );
XOR2_X1 U1087 ( .A(KEYINPUT40), .B(G119), .Z(n1357) );
XNOR2_X1 U1088 ( .A(G113), .B(G116), .ZN(n1356) );
XNOR2_X1 U1089 ( .A(n1358), .B(n1359), .ZN(n1121) );
XOR2_X1 U1090 ( .A(G107), .B(G104), .Z(n1359) );
NAND2_X1 U1091 ( .A1(KEYINPUT56), .A2(n1330), .ZN(n1358) );
INV_X1 U1092 ( .A(G101), .ZN(n1330) );
NAND3_X1 U1093 ( .A1(n1360), .A2(n1361), .A3(n1362), .ZN(n1349) );
OR2_X1 U1094 ( .A1(n1230), .A2(n1312), .ZN(n1362) );
NAND2_X1 U1095 ( .A1(KEYINPUT31), .A2(n1363), .ZN(n1361) );
NAND2_X1 U1096 ( .A1(n1364), .A2(n1312), .ZN(n1363) );
XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1230), .ZN(n1364) );
NAND2_X1 U1098 ( .A1(n1365), .A2(n1366), .ZN(n1360) );
INV_X1 U1099 ( .A(KEYINPUT31), .ZN(n1366) );
NAND2_X1 U1100 ( .A1(n1367), .A2(n1368), .ZN(n1365) );
OR2_X1 U1101 ( .A1(n1230), .A2(KEYINPUT52), .ZN(n1368) );
NAND3_X1 U1102 ( .A1(n1230), .A2(n1312), .A3(KEYINPUT52), .ZN(n1367) );
XOR2_X1 U1103 ( .A(G125), .B(KEYINPUT61), .Z(n1312) );
XOR2_X1 U1104 ( .A(G143), .B(n1313), .Z(n1230) );
XOR2_X1 U1105 ( .A(G128), .B(G146), .Z(n1313) );
NAND2_X1 U1106 ( .A1(G210), .A2(n1369), .ZN(n1092) );
AND2_X1 U1107 ( .A1(G214), .A2(n1369), .ZN(n1077) );
NAND2_X1 U1108 ( .A1(n1370), .A2(n1291), .ZN(n1369) );
INV_X1 U1109 ( .A(G902), .ZN(n1291) );
INV_X1 U1110 ( .A(G237), .ZN(n1370) );
endmodule


