//Key = 0011110010100011100001010110101001100001010001100101110011010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319;

XOR2_X1 U718 ( .A(G107), .B(n999), .Z(G9) );
NAND4_X1 U719 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(G75) );
NAND4_X1 U720 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1002) );
NOR3_X1 U721 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NOR2_X1 U722 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND3_X1 U723 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1008) );
NOR3_X1 U724 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1006) );
NOR2_X1 U725 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
XNOR2_X1 U726 ( .A(KEYINPUT42), .B(n1021), .ZN(n1020) );
NOR2_X1 U727 ( .A1(G469), .A2(n1022), .ZN(n1017) );
XOR2_X1 U728 ( .A(n1021), .B(KEYINPUT58), .Z(n1022) );
XNOR2_X1 U729 ( .A(G475), .B(n1023), .ZN(n1016) );
XOR2_X1 U730 ( .A(n1024), .B(n1025), .Z(n1004) );
NAND3_X1 U731 ( .A1(n1026), .A2(n1027), .A3(G952), .ZN(n1001) );
NAND2_X1 U732 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND3_X1 U733 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U734 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U735 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
OR2_X1 U736 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U737 ( .A1(n1039), .A2(n1040), .ZN(n1033) );
NAND2_X1 U738 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U739 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XOR2_X1 U740 ( .A(n1045), .B(KEYINPUT19), .Z(n1043) );
NAND4_X1 U741 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1028) );
AND2_X1 U742 ( .A1(n1039), .A2(n1035), .ZN(n1049) );
OR2_X1 U743 ( .A1(n1030), .A2(n1032), .ZN(n1048) );
NAND3_X1 U744 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1053), .ZN(n1052) );
NAND2_X1 U746 ( .A1(n1030), .A2(n1054), .ZN(n1053) );
NAND2_X1 U747 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
NAND2_X1 U748 ( .A1(n1057), .A2(n1054), .ZN(n1056) );
INV_X1 U749 ( .A(KEYINPUT31), .ZN(n1054) );
XOR2_X1 U750 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U751 ( .A(n1060), .B(n1061), .Z(n1059) );
NAND2_X1 U752 ( .A1(G953), .A2(n1062), .ZN(n1061) );
NAND2_X1 U753 ( .A1(G900), .A2(G227), .ZN(n1062) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U755 ( .A1(G953), .A2(n1065), .ZN(n1064) );
XOR2_X1 U756 ( .A(n1066), .B(n1067), .Z(n1063) );
XOR2_X1 U757 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U758 ( .A1(KEYINPUT39), .A2(n1070), .ZN(n1068) );
XOR2_X1 U759 ( .A(n1071), .B(n1072), .Z(n1066) );
NOR2_X1 U760 ( .A1(KEYINPUT32), .A2(n1073), .ZN(n1072) );
XOR2_X1 U761 ( .A(n1074), .B(n1075), .Z(n1071) );
NOR2_X1 U762 ( .A1(G134), .A2(KEYINPUT9), .ZN(n1075) );
AND2_X1 U763 ( .A1(n1076), .A2(n1003), .ZN(n1058) );
XOR2_X1 U764 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U765 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U767 ( .A(n1003), .B(KEYINPUT7), .Z(n1081) );
NAND4_X1 U768 ( .A1(n1083), .A2(n1084), .A3(KEYINPUT49), .A4(n1085), .ZN(n1079) );
NOR2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U770 ( .A1(G898), .A2(n1003), .ZN(n1087) );
INV_X1 U771 ( .A(n1088), .ZN(n1086) );
NAND2_X1 U772 ( .A1(KEYINPUT30), .A2(n1089), .ZN(n1084) );
NAND2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U774 ( .A1(n1092), .A2(n1093), .ZN(n1083) );
INV_X1 U775 ( .A(KEYINPUT30), .ZN(n1093) );
XOR2_X1 U776 ( .A(n1094), .B(n1095), .Z(n1092) );
NOR3_X1 U777 ( .A1(n1003), .A2(KEYINPUT43), .A3(n1096), .ZN(n1077) );
NOR2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U779 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XOR2_X1 U780 ( .A(n1101), .B(n1102), .Z(n1100) );
OR2_X1 U781 ( .A1(n1103), .A2(n1012), .ZN(n1101) );
NOR2_X1 U782 ( .A1(n1099), .A2(n1104), .ZN(G63) );
XOR2_X1 U783 ( .A(n1105), .B(n1106), .Z(n1104) );
AND2_X1 U784 ( .A1(G478), .A2(n1107), .ZN(n1106) );
NAND2_X1 U785 ( .A1(KEYINPUT52), .A2(n1108), .ZN(n1105) );
NOR3_X1 U786 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G60) );
NOR3_X1 U787 ( .A1(n1112), .A2(G953), .A3(G952), .ZN(n1111) );
AND2_X1 U788 ( .A1(n1112), .A2(n1099), .ZN(n1110) );
INV_X1 U789 ( .A(KEYINPUT47), .ZN(n1112) );
XOR2_X1 U790 ( .A(n1113), .B(n1114), .Z(n1109) );
NAND2_X1 U791 ( .A1(n1107), .A2(G475), .ZN(n1113) );
XOR2_X1 U792 ( .A(G104), .B(n1115), .Z(G6) );
NOR2_X1 U793 ( .A1(n1099), .A2(n1116), .ZN(G57) );
XOR2_X1 U794 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U795 ( .A(G101), .B(n1119), .ZN(n1118) );
NOR2_X1 U796 ( .A1(KEYINPUT40), .A2(n1120), .ZN(n1119) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U799 ( .A1(KEYINPUT13), .A2(n1125), .ZN(n1124) );
XOR2_X1 U800 ( .A(KEYINPUT51), .B(n1126), .Z(n1125) );
INV_X1 U801 ( .A(n1127), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1107), .A2(G472), .ZN(n1123) );
NAND2_X1 U803 ( .A1(KEYINPUT59), .A2(n1128), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1099), .A2(n1129), .ZN(G54) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U806 ( .A(n1127), .B(n1132), .Z(n1131) );
XOR2_X1 U807 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U808 ( .A(n1135), .B(n1136), .Z(n1130) );
XNOR2_X1 U809 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U810 ( .A1(G140), .A2(KEYINPUT44), .ZN(n1138) );
NOR3_X1 U811 ( .A1(n1103), .A2(KEYINPUT17), .A3(n1019), .ZN(n1137) );
INV_X1 U812 ( .A(G469), .ZN(n1019) );
INV_X1 U813 ( .A(n1107), .ZN(n1103) );
XOR2_X1 U814 ( .A(n1139), .B(KEYINPUT12), .Z(n1135) );
NOR2_X1 U815 ( .A1(n1140), .A2(n1141), .ZN(G51) );
XOR2_X1 U816 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U817 ( .A(n1144), .B(n1073), .Z(n1143) );
XOR2_X1 U818 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U819 ( .A1(n1107), .A2(n1025), .ZN(n1145) );
NOR2_X1 U820 ( .A1(n1147), .A2(n1000), .ZN(n1107) );
NOR2_X1 U821 ( .A1(n1076), .A2(n1082), .ZN(n1000) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1082) );
NOR4_X1 U823 ( .A1(n1150), .A2(n1151), .A3(n1115), .A4(n999), .ZN(n1149) );
AND3_X1 U824 ( .A1(n1039), .A2(n1152), .A3(n1153), .ZN(n999) );
AND3_X1 U825 ( .A1(n1039), .A2(n1152), .A3(n1154), .ZN(n1115) );
NOR4_X1 U826 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
INV_X1 U828 ( .A(n1161), .ZN(n1157) );
NAND4_X1 U829 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1076) );
AND4_X1 U830 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND3_X1 U831 ( .A1(n1170), .A2(n1153), .A3(n1035), .ZN(n1169) );
AND2_X1 U832 ( .A1(n1171), .A2(n1172), .ZN(n1164) );
XOR2_X1 U833 ( .A(n1173), .B(n1174), .Z(n1142) );
XOR2_X1 U834 ( .A(KEYINPUT5), .B(KEYINPUT36), .Z(n1174) );
XOR2_X1 U835 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U836 ( .A1(KEYINPUT6), .A2(n1177), .ZN(n1176) );
XOR2_X1 U837 ( .A(KEYINPUT25), .B(n1074), .Z(n1177) );
INV_X1 U838 ( .A(G125), .ZN(n1074) );
XNOR2_X1 U839 ( .A(n1099), .B(KEYINPUT10), .ZN(n1140) );
NOR2_X1 U840 ( .A1(n1003), .A2(G952), .ZN(n1099) );
XOR2_X1 U841 ( .A(n1178), .B(n1171), .Z(G48) );
NAND3_X1 U842 ( .A1(n1154), .A2(n1179), .A3(n1180), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1162), .B(n1181), .Z(G45) );
NOR2_X1 U844 ( .A1(G143), .A2(KEYINPUT62), .ZN(n1181) );
NAND4_X1 U845 ( .A1(n1170), .A2(n1179), .A3(n1182), .A4(n1183), .ZN(n1162) );
XNOR2_X1 U846 ( .A(n1163), .B(n1184), .ZN(G42) );
NOR2_X1 U847 ( .A1(KEYINPUT37), .A2(n1185), .ZN(n1184) );
XOR2_X1 U848 ( .A(KEYINPUT61), .B(G140), .Z(n1185) );
NAND4_X1 U849 ( .A1(n1154), .A2(n1035), .A3(n1038), .A4(n1186), .ZN(n1163) );
XOR2_X1 U850 ( .A(n1187), .B(n1168), .Z(G39) );
NAND3_X1 U851 ( .A1(n1180), .A2(n1035), .A3(n1032), .ZN(n1168) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(G36) );
NAND3_X1 U853 ( .A1(KEYINPUT3), .A2(n1190), .A3(n1191), .ZN(n1189) );
NAND2_X1 U854 ( .A1(G134), .A2(n1192), .ZN(n1188) );
NAND2_X1 U855 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U856 ( .A1(n1190), .A2(n1195), .ZN(n1194) );
INV_X1 U857 ( .A(KEYINPUT41), .ZN(n1195) );
NAND2_X1 U858 ( .A1(KEYINPUT41), .A2(n1196), .ZN(n1193) );
NAND2_X1 U859 ( .A1(KEYINPUT3), .A2(n1190), .ZN(n1196) );
AND3_X1 U860 ( .A1(n1153), .A2(n1197), .A3(n1170), .ZN(n1190) );
XOR2_X1 U861 ( .A(KEYINPUT0), .B(n1035), .Z(n1197) );
XOR2_X1 U862 ( .A(n1198), .B(n1167), .Z(G33) );
NAND3_X1 U863 ( .A1(n1154), .A2(n1035), .A3(n1170), .ZN(n1167) );
AND2_X1 U864 ( .A1(n1037), .A2(n1186), .ZN(n1170) );
NOR2_X1 U865 ( .A1(n1199), .A2(n1044), .ZN(n1035) );
INV_X1 U866 ( .A(n1013), .ZN(n1044) );
XOR2_X1 U867 ( .A(n1166), .B(n1200), .Z(G30) );
XNOR2_X1 U868 ( .A(G128), .B(KEYINPUT60), .ZN(n1200) );
NAND3_X1 U869 ( .A1(n1153), .A2(n1179), .A3(n1180), .ZN(n1166) );
AND3_X1 U870 ( .A1(n1010), .A2(n1201), .A3(n1186), .ZN(n1180) );
AND2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1186) );
INV_X1 U872 ( .A(n1050), .ZN(n1153) );
XOR2_X1 U873 ( .A(G101), .B(n1151), .Z(G3) );
AND3_X1 U874 ( .A1(n1037), .A2(n1152), .A3(n1032), .ZN(n1151) );
AND3_X1 U875 ( .A1(n1204), .A2(n1205), .A3(n1202), .ZN(n1152) );
INV_X1 U876 ( .A(n1206), .ZN(n1037) );
XOR2_X1 U877 ( .A(G125), .B(n1207), .Z(G27) );
NOR2_X1 U878 ( .A1(KEYINPUT55), .A2(n1172), .ZN(n1207) );
NAND4_X1 U879 ( .A1(n1030), .A2(n1154), .A3(n1208), .A4(n1038), .ZN(n1172) );
AND2_X1 U880 ( .A1(n1203), .A2(n1179), .ZN(n1208) );
NAND2_X1 U881 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NAND2_X1 U882 ( .A1(n1211), .A2(n1065), .ZN(n1210) );
INV_X1 U883 ( .A(G900), .ZN(n1065) );
INV_X1 U884 ( .A(n1051), .ZN(n1154) );
XOR2_X1 U885 ( .A(G122), .B(n1212), .Z(G24) );
NOR2_X1 U886 ( .A1(KEYINPUT38), .A2(n1161), .ZN(n1212) );
NAND4_X1 U887 ( .A1(n1182), .A2(n1183), .A3(n1179), .A4(n1213), .ZN(n1161) );
NOR2_X1 U888 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
INV_X1 U889 ( .A(n1039), .ZN(n1214) );
NOR2_X1 U890 ( .A1(n1201), .A2(n1010), .ZN(n1039) );
XOR2_X1 U891 ( .A(G119), .B(n1150), .Z(G21) );
NOR3_X1 U892 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1150) );
NAND3_X1 U893 ( .A1(n1179), .A2(n1201), .A3(n1010), .ZN(n1217) );
INV_X1 U894 ( .A(n1041), .ZN(n1179) );
XOR2_X1 U895 ( .A(G116), .B(n1156), .Z(G18) );
NOR4_X1 U896 ( .A1(n1215), .A2(n1206), .A3(n1050), .A4(n1041), .ZN(n1156) );
NAND2_X1 U897 ( .A1(n1218), .A2(n1182), .ZN(n1050) );
INV_X1 U898 ( .A(n1005), .ZN(n1182) );
XOR2_X1 U899 ( .A(G113), .B(n1155), .Z(G15) );
NOR4_X1 U900 ( .A1(n1215), .A2(n1206), .A3(n1159), .A4(n1051), .ZN(n1155) );
NAND2_X1 U901 ( .A1(n1005), .A2(n1183), .ZN(n1051) );
INV_X1 U902 ( .A(n1204), .ZN(n1159) );
NAND2_X1 U903 ( .A1(n1219), .A2(n1010), .ZN(n1206) );
NAND2_X1 U904 ( .A1(n1030), .A2(n1205), .ZN(n1215) );
AND2_X1 U905 ( .A1(n1057), .A2(n1015), .ZN(n1030) );
XNOR2_X1 U906 ( .A(G110), .B(n1220), .ZN(G12) );
NAND2_X1 U907 ( .A1(n1221), .A2(n1204), .ZN(n1220) );
XOR2_X1 U908 ( .A(n1041), .B(KEYINPUT15), .Z(n1204) );
NAND2_X1 U909 ( .A1(n1199), .A2(n1013), .ZN(n1041) );
NAND2_X1 U910 ( .A1(G214), .A2(n1222), .ZN(n1013) );
INV_X1 U911 ( .A(n1045), .ZN(n1199) );
XOR2_X1 U912 ( .A(n1223), .B(n1025), .Z(n1045) );
AND2_X1 U913 ( .A1(G210), .A2(n1222), .ZN(n1025) );
NAND2_X1 U914 ( .A1(n1224), .A2(n1147), .ZN(n1222) );
XOR2_X1 U915 ( .A(KEYINPUT23), .B(G237), .Z(n1224) );
XNOR2_X1 U916 ( .A(KEYINPUT20), .B(n1225), .ZN(n1223) );
NOR2_X1 U917 ( .A1(KEYINPUT54), .A2(n1024), .ZN(n1225) );
NAND3_X1 U918 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1024) );
OR2_X1 U919 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U920 ( .A1(n1229), .A2(n1231), .ZN(n1226) );
NAND2_X1 U921 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U922 ( .A1(KEYINPUT53), .A2(n1230), .ZN(n1233) );
OR2_X1 U923 ( .A1(KEYINPUT35), .A2(n1234), .ZN(n1230) );
OR2_X1 U924 ( .A1(n1234), .A2(KEYINPUT53), .ZN(n1232) );
XOR2_X1 U925 ( .A(n1175), .B(KEYINPUT21), .Z(n1234) );
NAND3_X1 U926 ( .A1(n1088), .A2(n1090), .A3(n1091), .ZN(n1175) );
NAND2_X1 U927 ( .A1(n1235), .A2(n1236), .ZN(n1091) );
INV_X1 U928 ( .A(n1094), .ZN(n1235) );
NAND3_X1 U929 ( .A1(n1237), .A2(n1094), .A3(n1095), .ZN(n1090) );
NAND2_X1 U930 ( .A1(n1238), .A2(n1239), .ZN(n1094) );
NAND2_X1 U931 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
NAND3_X1 U932 ( .A1(n1240), .A2(n1241), .A3(n1236), .ZN(n1088) );
INV_X1 U933 ( .A(n1095), .ZN(n1236) );
XOR2_X1 U934 ( .A(n1242), .B(n1134), .Z(n1095) );
XNOR2_X1 U935 ( .A(G122), .B(KEYINPUT11), .ZN(n1242) );
INV_X1 U936 ( .A(n1238), .ZN(n1241) );
XNOR2_X1 U937 ( .A(n1243), .B(n1244), .ZN(n1238) );
NOR2_X1 U938 ( .A1(G101), .A2(KEYINPUT1), .ZN(n1244) );
INV_X1 U939 ( .A(n1239), .ZN(n1240) );
XOR2_X1 U940 ( .A(n1245), .B(G113), .Z(n1239) );
NAND2_X1 U941 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U942 ( .A1(G116), .A2(n1248), .ZN(n1247) );
XOR2_X1 U943 ( .A(KEYINPUT26), .B(n1249), .Z(n1246) );
NOR2_X1 U944 ( .A1(G116), .A2(n1248), .ZN(n1249) );
XOR2_X1 U945 ( .A(n1073), .B(n1250), .Z(n1229) );
XNOR2_X1 U946 ( .A(n1251), .B(n1146), .ZN(n1250) );
NOR2_X1 U947 ( .A1(n1097), .A2(G953), .ZN(n1146) );
INV_X1 U948 ( .A(G224), .ZN(n1097) );
NAND2_X1 U949 ( .A1(KEYINPUT2), .A2(n1252), .ZN(n1251) );
XOR2_X1 U950 ( .A(KEYINPUT25), .B(G125), .Z(n1252) );
XOR2_X1 U951 ( .A(n1160), .B(KEYINPUT57), .Z(n1221) );
NAND4_X1 U952 ( .A1(n1032), .A2(n1038), .A3(n1202), .A4(n1205), .ZN(n1160) );
NAND2_X1 U953 ( .A1(n1209), .A2(n1253), .ZN(n1205) );
NAND2_X1 U954 ( .A1(n1211), .A2(n1098), .ZN(n1253) );
INV_X1 U955 ( .A(G898), .ZN(n1098) );
AND3_X1 U956 ( .A1(G902), .A2(n1027), .A3(G953), .ZN(n1211) );
NAND3_X1 U957 ( .A1(n1027), .A2(n1003), .A3(G952), .ZN(n1209) );
NAND2_X1 U958 ( .A1(n1254), .A2(G234), .ZN(n1027) );
XOR2_X1 U959 ( .A(n1255), .B(KEYINPUT4), .Z(n1254) );
NOR2_X1 U960 ( .A1(n1057), .A2(n1055), .ZN(n1202) );
INV_X1 U961 ( .A(n1015), .ZN(n1055) );
NAND2_X1 U962 ( .A1(G221), .A2(n1256), .ZN(n1015) );
XOR2_X1 U963 ( .A(n1021), .B(G469), .Z(n1057) );
NAND2_X1 U964 ( .A1(n1257), .A2(n1228), .ZN(n1021) );
XOR2_X1 U965 ( .A(n1133), .B(n1258), .Z(n1257) );
XNOR2_X1 U966 ( .A(n1259), .B(n1260), .ZN(n1258) );
NOR2_X1 U967 ( .A1(KEYINPUT50), .A2(n1127), .ZN(n1260) );
NOR2_X1 U968 ( .A1(KEYINPUT27), .A2(n1261), .ZN(n1259) );
XOR2_X1 U969 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U970 ( .A(n1070), .B(n1139), .Z(n1263) );
NAND2_X1 U971 ( .A1(G227), .A2(n1003), .ZN(n1139) );
INV_X1 U972 ( .A(G140), .ZN(n1070) );
XOR2_X1 U973 ( .A(n1264), .B(n1073), .Z(n1133) );
XNOR2_X1 U974 ( .A(G101), .B(n1243), .ZN(n1264) );
XOR2_X1 U975 ( .A(G104), .B(G107), .Z(n1243) );
NOR2_X1 U976 ( .A1(n1010), .A2(n1219), .ZN(n1038) );
INV_X1 U977 ( .A(n1201), .ZN(n1219) );
NAND3_X1 U978 ( .A1(n1265), .A2(n1266), .A3(n1014), .ZN(n1201) );
NAND2_X1 U979 ( .A1(n1011), .A2(n1012), .ZN(n1014) );
NAND2_X1 U980 ( .A1(KEYINPUT22), .A2(n1012), .ZN(n1266) );
OR3_X1 U981 ( .A1(n1011), .A2(KEYINPUT22), .A3(n1012), .ZN(n1265) );
NAND2_X1 U982 ( .A1(G217), .A2(n1256), .ZN(n1012) );
NAND2_X1 U983 ( .A1(G234), .A2(n1147), .ZN(n1256) );
INV_X1 U984 ( .A(G902), .ZN(n1147) );
AND2_X1 U985 ( .A1(n1102), .A2(n1228), .ZN(n1011) );
XNOR2_X1 U986 ( .A(n1267), .B(n1268), .ZN(n1102) );
XOR2_X1 U987 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U988 ( .A(G125), .B(n1271), .Z(n1270) );
NOR2_X1 U989 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U990 ( .A(n1274), .B(KEYINPUT33), .Z(n1273) );
NAND2_X1 U991 ( .A1(n1134), .A2(n1275), .ZN(n1274) );
NOR2_X1 U992 ( .A1(n1134), .A2(n1275), .ZN(n1272) );
NAND2_X1 U993 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
OR2_X1 U994 ( .A1(n1248), .A2(G128), .ZN(n1277) );
XOR2_X1 U995 ( .A(n1278), .B(KEYINPUT24), .Z(n1276) );
NAND2_X1 U996 ( .A1(G128), .A2(n1248), .ZN(n1278) );
INV_X1 U997 ( .A(n1262), .ZN(n1134) );
XNOR2_X1 U998 ( .A(G110), .B(KEYINPUT48), .ZN(n1262) );
AND2_X1 U999 ( .A1(n1279), .A2(G221), .ZN(n1269) );
XOR2_X1 U1000 ( .A(n1187), .B(n1280), .Z(n1267) );
XOR2_X1 U1001 ( .A(G146), .B(G140), .Z(n1280) );
INV_X1 U1002 ( .A(G137), .ZN(n1187) );
XNOR2_X1 U1003 ( .A(n1281), .B(G472), .ZN(n1010) );
NAND2_X1 U1004 ( .A1(n1282), .A2(n1228), .ZN(n1281) );
XOR2_X1 U1005 ( .A(n1121), .B(n1283), .Z(n1282) );
XOR2_X1 U1006 ( .A(n1284), .B(n1127), .Z(n1283) );
XOR2_X1 U1007 ( .A(n1191), .B(n1069), .Z(n1127) );
XOR2_X1 U1008 ( .A(G137), .B(G131), .Z(n1069) );
NAND2_X1 U1009 ( .A1(n1285), .A2(KEYINPUT46), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(n1128), .B(G101), .ZN(n1285) );
AND3_X1 U1011 ( .A1(n1255), .A2(n1003), .A3(G210), .ZN(n1128) );
XOR2_X1 U1012 ( .A(n1286), .B(n1287), .Z(n1121) );
XNOR2_X1 U1013 ( .A(G113), .B(n1288), .ZN(n1287) );
NAND2_X1 U1014 ( .A1(KEYINPUT56), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U1015 ( .A(n1073), .B(n1248), .ZN(n1286) );
XOR2_X1 U1016 ( .A(G119), .B(KEYINPUT8), .Z(n1248) );
XNOR2_X1 U1017 ( .A(n1178), .B(n1290), .ZN(n1073) );
INV_X1 U1018 ( .A(G146), .ZN(n1178) );
INV_X1 U1019 ( .A(n1216), .ZN(n1032) );
NAND2_X1 U1020 ( .A1(n1005), .A2(n1218), .ZN(n1216) );
INV_X1 U1021 ( .A(n1183), .ZN(n1218) );
NAND2_X1 U1022 ( .A1(n1291), .A2(n1292), .ZN(n1183) );
NAND2_X1 U1023 ( .A1(n1293), .A2(G475), .ZN(n1292) );
XOR2_X1 U1024 ( .A(KEYINPUT63), .B(n1294), .Z(n1291) );
NOR2_X1 U1025 ( .A1(G475), .A2(n1293), .ZN(n1294) );
XOR2_X1 U1026 ( .A(n1023), .B(KEYINPUT29), .Z(n1293) );
NAND2_X1 U1027 ( .A1(n1295), .A2(n1228), .ZN(n1023) );
XOR2_X1 U1028 ( .A(KEYINPUT16), .B(n1296), .Z(n1295) );
INV_X1 U1029 ( .A(n1114), .ZN(n1296) );
XOR2_X1 U1030 ( .A(n1297), .B(n1298), .Z(n1114) );
XOR2_X1 U1031 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1032 ( .A(G122), .B(G113), .Z(n1300) );
XOR2_X1 U1033 ( .A(G146), .B(G125), .Z(n1299) );
XOR2_X1 U1034 ( .A(n1301), .B(n1302), .Z(n1297) );
XNOR2_X1 U1035 ( .A(G104), .B(n1303), .ZN(n1302) );
NAND3_X1 U1036 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1303) );
OR2_X1 U1037 ( .A1(n1307), .A2(KEYINPUT34), .ZN(n1306) );
NAND3_X1 U1038 ( .A1(KEYINPUT34), .A2(n1307), .A3(G131), .ZN(n1305) );
NAND2_X1 U1039 ( .A1(n1308), .A2(n1198), .ZN(n1304) );
INV_X1 U1040 ( .A(G131), .ZN(n1198) );
NAND2_X1 U1041 ( .A1(KEYINPUT34), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1042 ( .A(KEYINPUT28), .B(n1307), .ZN(n1309) );
XOR2_X1 U1043 ( .A(n1310), .B(G143), .Z(n1307) );
NAND3_X1 U1044 ( .A1(n1255), .A2(n1003), .A3(G214), .ZN(n1310) );
INV_X1 U1045 ( .A(G237), .ZN(n1255) );
NAND2_X1 U1046 ( .A1(KEYINPUT45), .A2(G140), .ZN(n1301) );
XOR2_X1 U1047 ( .A(n1311), .B(G478), .Z(n1005) );
NAND2_X1 U1048 ( .A1(n1108), .A2(n1228), .ZN(n1311) );
XOR2_X1 U1049 ( .A(G902), .B(KEYINPUT14), .Z(n1228) );
XNOR2_X1 U1050 ( .A(n1312), .B(n1313), .ZN(n1108) );
XOR2_X1 U1051 ( .A(n1191), .B(n1314), .Z(n1313) );
NAND2_X1 U1052 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1053 ( .A1(G107), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1054 ( .A(n1318), .B(KEYINPUT18), .Z(n1315) );
OR2_X1 U1055 ( .A1(n1317), .A2(G107), .ZN(n1318) );
XNOR2_X1 U1056 ( .A(n1289), .B(G122), .ZN(n1317) );
INV_X1 U1057 ( .A(G116), .ZN(n1289) );
INV_X1 U1058 ( .A(G134), .ZN(n1191) );
XOR2_X1 U1059 ( .A(n1319), .B(n1290), .Z(n1312) );
XOR2_X1 U1060 ( .A(G143), .B(G128), .Z(n1290) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1279), .ZN(n1319) );
AND2_X1 U1062 ( .A1(G234), .A2(n1003), .ZN(n1279) );
INV_X1 U1063 ( .A(G953), .ZN(n1003) );
endmodule


