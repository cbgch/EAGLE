//Key = 0010110100100001010111101001000110110110000111000010000011001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405;

XNOR2_X1 U762 ( .A(G107), .B(n1055), .ZN(G9) );
NOR2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR4_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
INV_X1 U765 ( .A(G952), .ZN(n1060) );
NAND4_X1 U766 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1058) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1070) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1068) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U778 ( .A1(n1089), .A2(n1090), .A3(KEYINPUT10), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1072), .A2(n1091), .ZN(n1063) );
NAND2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1085), .A2(n1094), .ZN(n1093) );
XOR2_X1 U782 ( .A(n1095), .B(KEYINPUT12), .Z(n1092) );
NAND3_X1 U783 ( .A1(n1096), .A2(n1097), .A3(n1085), .ZN(n1095) );
XNOR2_X1 U784 ( .A(KEYINPUT39), .B(n1098), .ZN(n1097) );
NAND2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1062) );
INV_X1 U786 ( .A(KEYINPUT10), .ZN(n1100) );
NAND4_X1 U787 ( .A1(n1085), .A2(n1089), .A3(n1066), .A4(n1090), .ZN(n1099) );
AND3_X1 U788 ( .A1(n1079), .A2(n1071), .A3(n1075), .ZN(n1085) );
NOR3_X1 U789 ( .A1(n1061), .A2(n1101), .A3(n1102), .ZN(n1056) );
XNOR2_X1 U790 ( .A(G952), .B(KEYINPUT35), .ZN(n1102) );
INV_X1 U791 ( .A(n1065), .ZN(n1101) );
NAND4_X1 U792 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1065) );
NOR4_X1 U793 ( .A1(n1107), .A2(n1089), .A3(n1108), .A4(n1109), .ZN(n1106) );
XOR2_X1 U794 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U795 ( .A1(KEYINPUT60), .A2(n1112), .ZN(n1110) );
INV_X1 U796 ( .A(n1113), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1108) );
XOR2_X1 U798 ( .A(KEYINPUT49), .B(G475), .Z(n1115) );
NAND2_X1 U799 ( .A1(KEYINPUT50), .A2(n1116), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1117), .A2(n1084), .ZN(n1105) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U802 ( .A(KEYINPUT22), .B(n1120), .ZN(n1119) );
XNOR2_X1 U803 ( .A(G469), .B(n1121), .ZN(n1104) );
NAND2_X1 U804 ( .A1(KEYINPUT34), .A2(n1122), .ZN(n1121) );
XOR2_X1 U805 ( .A(G472), .B(n1123), .Z(n1103) );
NOR2_X1 U806 ( .A1(n1124), .A2(KEYINPUT59), .ZN(n1123) );
XOR2_X1 U807 ( .A(n1125), .B(n1126), .Z(G72) );
XOR2_X1 U808 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
AND2_X1 U810 ( .A1(G227), .A2(G900), .ZN(n1129) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
NAND2_X1 U812 ( .A1(G953), .A2(n1133), .ZN(n1132) );
XOR2_X1 U813 ( .A(n1134), .B(n1135), .Z(n1131) );
XNOR2_X1 U814 ( .A(n1136), .B(n1137), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1138), .ZN(n1125) );
NAND2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(G69) );
NAND3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
XOR2_X1 U818 ( .A(n1144), .B(KEYINPUT6), .Z(n1143) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1141) );
NAND2_X1 U820 ( .A1(n1147), .A2(n1148), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1149), .A2(n1144), .ZN(n1148) );
NAND2_X1 U822 ( .A1(G953), .A2(n1150), .ZN(n1144) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1150) );
OR2_X1 U824 ( .A1(n1142), .A2(KEYINPUT6), .ZN(n1149) );
INV_X1 U825 ( .A(KEYINPUT1), .ZN(n1142) );
XNOR2_X1 U826 ( .A(n1145), .B(n1146), .ZN(n1147) );
AND2_X1 U827 ( .A1(n1130), .A2(n1151), .ZN(n1146) );
NOR2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1145) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1152) );
NOR2_X1 U830 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XOR2_X1 U831 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U832 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1156), .A2(n1162), .ZN(G63) );
NOR3_X1 U834 ( .A1(n1113), .A2(n1163), .A3(n1164), .ZN(n1162) );
AND3_X1 U835 ( .A1(n1165), .A2(G478), .A3(n1166), .ZN(n1164) );
NOR2_X1 U836 ( .A1(n1167), .A2(n1165), .ZN(n1163) );
AND2_X1 U837 ( .A1(n1059), .A2(G478), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1156), .A2(n1168), .ZN(G60) );
XNOR2_X1 U839 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U840 ( .A(KEYINPUT8), .B(n1171), .Z(n1170) );
AND2_X1 U841 ( .A1(G475), .A2(n1166), .ZN(n1171) );
XOR2_X1 U842 ( .A(n1172), .B(n1173), .Z(G6) );
NAND2_X1 U843 ( .A1(KEYINPUT61), .A2(G104), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1156), .A2(n1174), .ZN(G57) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U846 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NAND2_X1 U847 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
INV_X1 U848 ( .A(n1181), .ZN(n1180) );
XOR2_X1 U849 ( .A(KEYINPUT63), .B(n1182), .Z(n1179) );
NAND2_X1 U850 ( .A1(n1182), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U851 ( .A(n1183), .B(n1184), .ZN(n1181) );
NOR2_X1 U852 ( .A1(KEYINPUT51), .A2(n1185), .ZN(n1184) );
NAND3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1183) );
NAND2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U855 ( .A1(KEYINPUT29), .A2(n1191), .ZN(n1187) );
NAND2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U857 ( .A(KEYINPUT32), .B(n1137), .ZN(n1192) );
NAND2_X1 U858 ( .A1(n1194), .A2(n1195), .ZN(n1186) );
INV_X1 U859 ( .A(KEYINPUT29), .ZN(n1195) );
NAND2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NAND3_X1 U861 ( .A1(KEYINPUT32), .A2(n1193), .A3(n1137), .ZN(n1197) );
OR2_X1 U862 ( .A1(n1137), .A2(KEYINPUT32), .ZN(n1196) );
AND2_X1 U863 ( .A1(n1166), .A2(G472), .ZN(n1182) );
INV_X1 U864 ( .A(n1161), .ZN(n1166) );
NOR2_X1 U865 ( .A1(n1156), .A2(n1198), .ZN(G54) );
NOR2_X1 U866 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U867 ( .A(n1201), .B(KEYINPUT19), .Z(n1200) );
NAND2_X1 U868 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U869 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
XNOR2_X1 U870 ( .A(n1204), .B(n1205), .ZN(n1203) );
NAND2_X1 U871 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
NAND2_X1 U872 ( .A1(n1208), .A2(n1137), .ZN(n1207) );
XOR2_X1 U873 ( .A(KEYINPUT17), .B(n1209), .Z(n1206) );
NOR2_X1 U874 ( .A1(n1137), .A2(n1208), .ZN(n1209) );
INV_X1 U875 ( .A(n1190), .ZN(n1137) );
NOR2_X1 U876 ( .A1(n1161), .A2(n1210), .ZN(n1202) );
NOR2_X1 U877 ( .A1(n1130), .A2(G952), .ZN(n1156) );
NOR2_X1 U878 ( .A1(n1211), .A2(n1212), .ZN(G51) );
XOR2_X1 U879 ( .A(n1213), .B(n1214), .Z(n1212) );
XNOR2_X1 U880 ( .A(n1193), .B(n1215), .ZN(n1214) );
XOR2_X1 U881 ( .A(n1216), .B(n1217), .Z(n1213) );
XOR2_X1 U882 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U883 ( .A1(n1120), .A2(n1161), .ZN(n1219) );
NAND2_X1 U884 ( .A1(G902), .A2(n1059), .ZN(n1161) );
OR2_X1 U885 ( .A1(n1151), .A2(n1138), .ZN(n1059) );
NAND4_X1 U886 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1138) );
NOR4_X1 U887 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
INV_X1 U888 ( .A(n1228), .ZN(n1226) );
NAND2_X1 U889 ( .A1(n1072), .A2(n1229), .ZN(n1222) );
NAND2_X1 U890 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U891 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XNOR2_X1 U892 ( .A(KEYINPUT53), .B(n1077), .ZN(n1233) );
NAND2_X1 U893 ( .A1(n1234), .A2(n1079), .ZN(n1230) );
NAND3_X1 U894 ( .A1(n1235), .A2(n1236), .A3(n1232), .ZN(n1220) );
NAND4_X1 U895 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1151) );
AND4_X1 U896 ( .A1(n1241), .A2(n1172), .A3(n1055), .A4(n1242), .ZN(n1240) );
NAND3_X1 U897 ( .A1(n1075), .A2(n1243), .A3(n1244), .ZN(n1055) );
NAND3_X1 U898 ( .A1(n1244), .A2(n1075), .A3(n1245), .ZN(n1172) );
NOR3_X1 U899 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1239) );
NOR2_X1 U900 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
AND4_X1 U901 ( .A1(n1249), .A2(n1251), .A3(n1066), .A4(n1235), .ZN(n1247) );
AND3_X1 U902 ( .A1(n1252), .A2(n1087), .A3(n1075), .ZN(n1251) );
INV_X1 U903 ( .A(KEYINPUT20), .ZN(n1249) );
NAND2_X1 U904 ( .A1(KEYINPUT37), .A2(n1253), .ZN(n1216) );
NOR2_X1 U905 ( .A1(n1254), .A2(n1130), .ZN(n1211) );
XNOR2_X1 U906 ( .A(G952), .B(KEYINPUT45), .ZN(n1254) );
XOR2_X1 U907 ( .A(G146), .B(n1225), .Z(G48) );
AND3_X1 U908 ( .A1(n1245), .A2(n1236), .A3(n1234), .ZN(n1225) );
XNOR2_X1 U909 ( .A(G143), .B(n1255), .ZN(G45) );
NAND3_X1 U910 ( .A1(n1235), .A2(n1256), .A3(n1232), .ZN(n1255) );
XNOR2_X1 U911 ( .A(KEYINPUT26), .B(n1087), .ZN(n1256) );
INV_X1 U912 ( .A(n1236), .ZN(n1087) );
XNOR2_X1 U913 ( .A(G140), .B(n1221), .ZN(G42) );
NAND3_X1 U914 ( .A1(n1257), .A2(n1094), .A3(n1072), .ZN(n1221) );
XNOR2_X1 U915 ( .A(G137), .B(n1258), .ZN(G39) );
NAND3_X1 U916 ( .A1(n1259), .A2(n1079), .A3(n1234), .ZN(n1258) );
XOR2_X1 U917 ( .A(KEYINPUT14), .B(n1072), .Z(n1259) );
NAND3_X1 U918 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(G36) );
NAND2_X1 U919 ( .A1(n1227), .A2(n1263), .ZN(n1262) );
NAND2_X1 U920 ( .A1(KEYINPUT28), .A2(n1264), .ZN(n1261) );
NAND2_X1 U921 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XNOR2_X1 U922 ( .A(KEYINPUT54), .B(n1263), .ZN(n1265) );
NAND2_X1 U923 ( .A1(n1267), .A2(n1268), .ZN(n1260) );
INV_X1 U924 ( .A(KEYINPUT28), .ZN(n1268) );
NAND2_X1 U925 ( .A1(n1269), .A2(n1270), .ZN(n1267) );
OR3_X1 U926 ( .A1(n1263), .A2(n1227), .A3(KEYINPUT54), .ZN(n1270) );
INV_X1 U927 ( .A(n1266), .ZN(n1227) );
NAND3_X1 U928 ( .A1(n1232), .A2(n1243), .A3(n1072), .ZN(n1266) );
NOR3_X1 U929 ( .A1(n1081), .A2(n1271), .A3(n1272), .ZN(n1232) );
INV_X1 U930 ( .A(n1273), .ZN(n1081) );
NAND2_X1 U931 ( .A1(KEYINPUT54), .A2(n1263), .ZN(n1269) );
XNOR2_X1 U932 ( .A(G131), .B(n1274), .ZN(G33) );
NAND3_X1 U933 ( .A1(n1072), .A2(n1273), .A3(n1275), .ZN(n1274) );
NOR3_X1 U934 ( .A1(n1077), .A2(n1276), .A3(n1271), .ZN(n1275) );
INV_X1 U935 ( .A(n1094), .ZN(n1271) );
XNOR2_X1 U936 ( .A(n1277), .B(KEYINPUT33), .ZN(n1276) );
AND2_X1 U937 ( .A1(n1090), .A2(n1278), .ZN(n1072) );
XNOR2_X1 U938 ( .A(n1279), .B(n1224), .ZN(G30) );
AND3_X1 U939 ( .A1(n1243), .A2(n1236), .A3(n1234), .ZN(n1224) );
AND4_X1 U940 ( .A1(n1277), .A2(n1094), .A3(n1280), .A4(n1084), .ZN(n1234) );
XNOR2_X1 U941 ( .A(G101), .B(n1241), .ZN(G3) );
NAND3_X1 U942 ( .A1(n1244), .A2(n1079), .A3(n1273), .ZN(n1241) );
XNOR2_X1 U943 ( .A(n1253), .B(n1281), .ZN(G27) );
NOR2_X1 U944 ( .A1(KEYINPUT47), .A2(n1228), .ZN(n1281) );
NAND3_X1 U945 ( .A1(n1066), .A2(n1236), .A3(n1257), .ZN(n1228) );
AND4_X1 U946 ( .A1(n1277), .A2(n1245), .A3(n1083), .A4(n1084), .ZN(n1257) );
INV_X1 U947 ( .A(n1272), .ZN(n1277) );
NAND2_X1 U948 ( .A1(n1071), .A2(n1282), .ZN(n1272) );
NAND2_X1 U949 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND3_X1 U950 ( .A1(G953), .A2(n1133), .A3(G902), .ZN(n1283) );
INV_X1 U951 ( .A(G900), .ZN(n1133) );
NAND3_X1 U952 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(G24) );
NAND2_X1 U953 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U954 ( .A1(KEYINPUT31), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U955 ( .A(KEYINPUT4), .B(n1250), .ZN(n1290) );
NAND3_X1 U956 ( .A1(KEYINPUT31), .A2(G122), .A3(n1250), .ZN(n1286) );
OR2_X1 U957 ( .A1(n1250), .A2(KEYINPUT31), .ZN(n1285) );
NAND3_X1 U958 ( .A1(n1291), .A2(n1075), .A3(n1235), .ZN(n1250) );
NOR2_X1 U959 ( .A1(n1292), .A2(n1293), .ZN(n1235) );
NOR2_X1 U960 ( .A1(n1084), .A2(n1280), .ZN(n1075) );
XOR2_X1 U961 ( .A(G119), .B(n1246), .Z(G21) );
AND4_X1 U962 ( .A1(n1291), .A2(n1079), .A3(n1280), .A4(n1084), .ZN(n1246) );
XNOR2_X1 U963 ( .A(G116), .B(n1237), .ZN(G18) );
NAND3_X1 U964 ( .A1(n1273), .A2(n1243), .A3(n1291), .ZN(n1237) );
INV_X1 U965 ( .A(n1078), .ZN(n1243) );
NAND2_X1 U966 ( .A1(n1294), .A2(n1295), .ZN(n1078) );
XNOR2_X1 U967 ( .A(KEYINPUT27), .B(n1293), .ZN(n1294) );
XNOR2_X1 U968 ( .A(G113), .B(n1238), .ZN(G15) );
NAND3_X1 U969 ( .A1(n1273), .A2(n1245), .A3(n1291), .ZN(n1238) );
AND3_X1 U970 ( .A1(n1252), .A2(n1236), .A3(n1066), .ZN(n1291) );
NOR2_X1 U971 ( .A1(n1296), .A2(n1107), .ZN(n1066) );
NOR2_X1 U972 ( .A1(n1084), .A2(n1083), .ZN(n1273) );
XNOR2_X1 U973 ( .A(G110), .B(n1242), .ZN(G12) );
NAND4_X1 U974 ( .A1(n1083), .A2(n1244), .A3(n1079), .A4(n1084), .ZN(n1242) );
XOR2_X1 U975 ( .A(n1297), .B(n1160), .Z(n1084) );
NAND2_X1 U976 ( .A1(G217), .A2(n1298), .ZN(n1160) );
OR2_X1 U977 ( .A1(n1159), .A2(G902), .ZN(n1297) );
XNOR2_X1 U978 ( .A(n1299), .B(n1300), .ZN(n1159) );
AND2_X1 U979 ( .A1(G221), .A2(n1301), .ZN(n1300) );
XOR2_X1 U980 ( .A(n1302), .B(G137), .Z(n1299) );
NAND2_X1 U981 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U982 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U983 ( .A(n1307), .B(KEYINPUT46), .Z(n1303) );
OR2_X1 U984 ( .A1(n1306), .A2(n1305), .ZN(n1307) );
XNOR2_X1 U985 ( .A(G146), .B(n1308), .ZN(n1305) );
NOR2_X1 U986 ( .A1(KEYINPUT48), .A2(n1136), .ZN(n1308) );
NAND2_X1 U987 ( .A1(n1309), .A2(n1310), .ZN(n1136) );
NAND2_X1 U988 ( .A1(n1253), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U989 ( .A(n1312), .B(n1313), .ZN(n1306) );
XNOR2_X1 U990 ( .A(G110), .B(G128), .ZN(n1312) );
NAND2_X1 U991 ( .A1(n1314), .A2(n1315), .ZN(n1079) );
OR2_X1 U992 ( .A1(n1077), .A2(KEYINPUT27), .ZN(n1315) );
INV_X1 U993 ( .A(n1245), .ZN(n1077) );
NOR2_X1 U994 ( .A1(n1293), .A2(n1295), .ZN(n1245) );
INV_X1 U995 ( .A(n1292), .ZN(n1295) );
NAND3_X1 U996 ( .A1(n1293), .A2(n1292), .A3(KEYINPUT27), .ZN(n1314) );
XOR2_X1 U997 ( .A(n1113), .B(n1316), .Z(n1292) );
NOR2_X1 U998 ( .A1(KEYINPUT9), .A2(n1111), .ZN(n1316) );
XOR2_X1 U999 ( .A(G478), .B(KEYINPUT41), .Z(n1111) );
NOR2_X1 U1000 ( .A1(n1165), .A2(G902), .ZN(n1113) );
XNOR2_X1 U1001 ( .A(n1317), .B(n1318), .ZN(n1165) );
XNOR2_X1 U1002 ( .A(n1279), .B(n1319), .ZN(n1318) );
XNOR2_X1 U1003 ( .A(n1320), .B(G134), .ZN(n1319) );
INV_X1 U1004 ( .A(G128), .ZN(n1279) );
XOR2_X1 U1005 ( .A(n1321), .B(n1322), .Z(n1317) );
NOR2_X1 U1006 ( .A1(KEYINPUT0), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1007 ( .A(n1324), .B(n1325), .ZN(n1323) );
XNOR2_X1 U1008 ( .A(n1289), .B(G116), .ZN(n1325) );
NAND2_X1 U1009 ( .A1(n1301), .A2(G217), .ZN(n1321) );
AND2_X1 U1010 ( .A1(G234), .A2(n1130), .ZN(n1301) );
XNOR2_X1 U1011 ( .A(n1116), .B(n1326), .ZN(n1293) );
XOR2_X1 U1012 ( .A(KEYINPUT44), .B(G475), .Z(n1326) );
NAND2_X1 U1013 ( .A1(n1169), .A2(n1327), .ZN(n1116) );
XNOR2_X1 U1014 ( .A(n1328), .B(n1329), .ZN(n1169) );
XOR2_X1 U1015 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1016 ( .A(n1332), .B(n1333), .ZN(n1331) );
NOR2_X1 U1017 ( .A1(KEYINPUT13), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1018 ( .A(n1335), .B(G146), .Z(n1334) );
NAND2_X1 U1019 ( .A1(n1336), .A2(n1309), .ZN(n1335) );
NAND2_X1 U1020 ( .A1(G125), .A2(G140), .ZN(n1309) );
NAND2_X1 U1021 ( .A1(n1337), .A2(n1311), .ZN(n1336) );
XNOR2_X1 U1022 ( .A(G125), .B(KEYINPUT18), .ZN(n1337) );
NAND2_X1 U1023 ( .A1(KEYINPUT7), .A2(n1338), .ZN(n1332) );
XNOR2_X1 U1024 ( .A(n1289), .B(G113), .ZN(n1338) );
INV_X1 U1025 ( .A(G122), .ZN(n1289) );
AND2_X1 U1026 ( .A1(G214), .A2(n1339), .ZN(n1330) );
XNOR2_X1 U1027 ( .A(G104), .B(n1340), .ZN(n1328) );
XNOR2_X1 U1028 ( .A(n1320), .B(G131), .ZN(n1340) );
AND3_X1 U1029 ( .A1(n1094), .A2(n1236), .A3(n1252), .ZN(n1244) );
AND2_X1 U1030 ( .A1(n1341), .A2(n1071), .ZN(n1252) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1071) );
NAND2_X1 U1032 ( .A1(n1284), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1033 ( .A1(G902), .A2(n1153), .ZN(n1342) );
NOR2_X1 U1034 ( .A1(n1130), .A2(G898), .ZN(n1153) );
NAND2_X1 U1035 ( .A1(n1343), .A2(G952), .ZN(n1284) );
XNOR2_X1 U1036 ( .A(n1061), .B(KEYINPUT42), .ZN(n1343) );
XOR2_X1 U1037 ( .A(G953), .B(KEYINPUT58), .Z(n1061) );
NOR2_X1 U1038 ( .A1(n1090), .A2(n1089), .ZN(n1236) );
INV_X1 U1039 ( .A(n1278), .ZN(n1089) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1344), .ZN(n1278) );
XOR2_X1 U1041 ( .A(n1345), .B(n1120), .Z(n1090) );
NAND2_X1 U1042 ( .A1(G210), .A2(n1344), .ZN(n1120) );
NAND2_X1 U1043 ( .A1(n1346), .A2(n1327), .ZN(n1344) );
INV_X1 U1044 ( .A(G237), .ZN(n1346) );
NAND2_X1 U1045 ( .A1(KEYINPUT21), .A2(n1118), .ZN(n1345) );
NAND3_X1 U1046 ( .A1(n1347), .A2(n1327), .A3(n1348), .ZN(n1118) );
XOR2_X1 U1047 ( .A(n1349), .B(KEYINPUT36), .Z(n1348) );
OR2_X1 U1048 ( .A1(n1350), .A2(n1215), .ZN(n1349) );
NAND2_X1 U1049 ( .A1(n1215), .A2(n1350), .ZN(n1347) );
XNOR2_X1 U1050 ( .A(n1351), .B(n1218), .ZN(n1350) );
AND2_X1 U1051 ( .A1(G224), .A2(n1130), .ZN(n1218) );
NAND3_X1 U1052 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
NAND2_X1 U1053 ( .A1(G125), .A2(n1193), .ZN(n1354) );
NAND2_X1 U1054 ( .A1(KEYINPUT23), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1055 ( .A1(n1356), .A2(n1253), .ZN(n1355) );
INV_X1 U1056 ( .A(G125), .ZN(n1253) );
XNOR2_X1 U1057 ( .A(KEYINPUT11), .B(n1193), .ZN(n1356) );
NAND2_X1 U1058 ( .A1(n1357), .A2(n1358), .ZN(n1352) );
INV_X1 U1059 ( .A(KEYINPUT23), .ZN(n1358) );
NAND2_X1 U1060 ( .A1(n1359), .A2(n1360), .ZN(n1357) );
OR3_X1 U1061 ( .A1(G125), .A2(KEYINPUT11), .A3(n1193), .ZN(n1360) );
NAND2_X1 U1062 ( .A1(KEYINPUT11), .A2(n1193), .ZN(n1359) );
INV_X1 U1063 ( .A(n1189), .ZN(n1193) );
XOR2_X1 U1064 ( .A(n1361), .B(n1155), .Z(n1215) );
XOR2_X1 U1065 ( .A(n1362), .B(n1363), .Z(n1155) );
XNOR2_X1 U1066 ( .A(G101), .B(n1364), .ZN(n1363) );
NAND3_X1 U1067 ( .A1(n1365), .A2(n1366), .A3(KEYINPUT24), .ZN(n1364) );
NAND2_X1 U1068 ( .A1(KEYINPUT43), .A2(n1367), .ZN(n1366) );
XNOR2_X1 U1069 ( .A(G104), .B(G107), .ZN(n1367) );
OR3_X1 U1070 ( .A1(n1324), .A2(G104), .A3(KEYINPUT43), .ZN(n1365) );
XNOR2_X1 U1071 ( .A(G110), .B(G122), .ZN(n1362) );
NAND2_X1 U1072 ( .A1(n1154), .A2(n1368), .ZN(n1361) );
XOR2_X1 U1073 ( .A(KEYINPUT62), .B(KEYINPUT16), .Z(n1368) );
AND2_X1 U1074 ( .A1(n1369), .A2(n1370), .ZN(n1154) );
OR2_X1 U1075 ( .A1(n1185), .A2(KEYINPUT55), .ZN(n1370) );
NAND3_X1 U1076 ( .A1(G113), .A2(n1371), .A3(KEYINPUT55), .ZN(n1369) );
NOR2_X1 U1077 ( .A1(n1096), .A2(n1107), .ZN(n1094) );
INV_X1 U1078 ( .A(n1098), .ZN(n1107) );
NAND2_X1 U1079 ( .A1(G221), .A2(n1298), .ZN(n1098) );
NAND2_X1 U1080 ( .A1(G234), .A2(n1327), .ZN(n1298) );
INV_X1 U1081 ( .A(n1296), .ZN(n1096) );
XOR2_X1 U1082 ( .A(n1122), .B(n1210), .Z(n1296) );
INV_X1 U1083 ( .A(G469), .ZN(n1210) );
NAND2_X1 U1084 ( .A1(n1372), .A2(n1327), .ZN(n1122) );
XNOR2_X1 U1085 ( .A(n1190), .B(n1373), .ZN(n1372) );
XNOR2_X1 U1086 ( .A(n1374), .B(n1375), .ZN(n1373) );
NOR2_X1 U1087 ( .A1(KEYINPUT52), .A2(n1208), .ZN(n1375) );
XNOR2_X1 U1088 ( .A(n1376), .B(n1377), .ZN(n1208) );
NOR2_X1 U1089 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
NOR2_X1 U1090 ( .A1(KEYINPUT3), .A2(n1380), .ZN(n1379) );
INV_X1 U1091 ( .A(n1381), .ZN(n1380) );
NOR2_X1 U1092 ( .A1(KEYINPUT57), .A2(n1381), .ZN(n1378) );
NAND2_X1 U1093 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
NAND2_X1 U1094 ( .A1(G104), .A2(n1324), .ZN(n1383) );
XOR2_X1 U1095 ( .A(KEYINPUT56), .B(n1384), .Z(n1382) );
NOR2_X1 U1096 ( .A1(n1385), .A2(n1324), .ZN(n1384) );
INV_X1 U1097 ( .A(G107), .ZN(n1324) );
XNOR2_X1 U1098 ( .A(G104), .B(KEYINPUT15), .ZN(n1385) );
XNOR2_X1 U1099 ( .A(n1135), .B(G101), .ZN(n1376) );
XOR2_X1 U1100 ( .A(G128), .B(n1386), .Z(n1135) );
NOR2_X1 U1101 ( .A1(n1205), .A2(KEYINPUT25), .ZN(n1374) );
AND2_X1 U1102 ( .A1(n1387), .A2(n1388), .ZN(n1205) );
NAND3_X1 U1103 ( .A1(G227), .A2(n1130), .A3(n1389), .ZN(n1388) );
XNOR2_X1 U1104 ( .A(G110), .B(G140), .ZN(n1389) );
NAND2_X1 U1105 ( .A1(n1390), .A2(n1391), .ZN(n1387) );
NAND2_X1 U1106 ( .A1(G227), .A2(n1130), .ZN(n1391) );
INV_X1 U1107 ( .A(G953), .ZN(n1130) );
XNOR2_X1 U1108 ( .A(n1311), .B(G110), .ZN(n1390) );
INV_X1 U1109 ( .A(G140), .ZN(n1311) );
INV_X1 U1110 ( .A(n1280), .ZN(n1083) );
XOR2_X1 U1111 ( .A(n1124), .B(G472), .Z(n1280) );
AND3_X1 U1112 ( .A1(n1392), .A2(n1393), .A3(n1327), .ZN(n1124) );
INV_X1 U1113 ( .A(G902), .ZN(n1327) );
NAND2_X1 U1114 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
INV_X1 U1115 ( .A(KEYINPUT30), .ZN(n1395) );
XOR2_X1 U1116 ( .A(n1396), .B(n1397), .Z(n1394) );
NAND3_X1 U1117 ( .A1(n1397), .A2(n1396), .A3(KEYINPUT30), .ZN(n1392) );
XOR2_X1 U1118 ( .A(n1398), .B(n1399), .Z(n1396) );
XNOR2_X1 U1119 ( .A(n1185), .B(n1189), .ZN(n1399) );
XOR2_X1 U1120 ( .A(G128), .B(n1400), .Z(n1189) );
NOR2_X1 U1121 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
NOR3_X1 U1122 ( .A1(KEYINPUT38), .A2(G146), .A3(n1320), .ZN(n1402) );
NOR2_X1 U1123 ( .A1(n1386), .A2(n1403), .ZN(n1401) );
INV_X1 U1124 ( .A(KEYINPUT38), .ZN(n1403) );
XNOR2_X1 U1125 ( .A(n1320), .B(G146), .ZN(n1386) );
INV_X1 U1126 ( .A(G143), .ZN(n1320) );
XNOR2_X1 U1127 ( .A(n1371), .B(G113), .ZN(n1185) );
XOR2_X1 U1128 ( .A(G116), .B(n1313), .Z(n1371) );
XOR2_X1 U1129 ( .A(G119), .B(KEYINPUT40), .Z(n1313) );
XNOR2_X1 U1130 ( .A(n1190), .B(KEYINPUT2), .ZN(n1398) );
XOR2_X1 U1131 ( .A(G131), .B(n1404), .Z(n1190) );
XNOR2_X1 U1132 ( .A(G137), .B(n1263), .ZN(n1404) );
INV_X1 U1133 ( .A(G134), .ZN(n1263) );
XOR2_X1 U1134 ( .A(n1176), .B(KEYINPUT5), .Z(n1397) );
XNOR2_X1 U1135 ( .A(n1405), .B(G101), .ZN(n1176) );
NAND2_X1 U1136 ( .A1(n1339), .A2(G210), .ZN(n1405) );
NOR2_X1 U1137 ( .A1(G953), .A2(G237), .ZN(n1339) );
endmodule


