//Key = 1110000111100001100010100110111000101001110111110111100010011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330;

XNOR2_X1 U744 ( .A(G107), .B(n1016), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1018) );
NOR2_X1 U747 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U748 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U749 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR2_X1 U750 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR3_X1 U751 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR3_X1 U752 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NOR3_X1 U753 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1032) );
NOR2_X1 U754 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(n1038) );
XNOR2_X1 U756 ( .A(n1044), .B(KEYINPUT4), .ZN(n1043) );
NOR3_X1 U757 ( .A1(n1034), .A2(n1045), .A3(n1040), .ZN(n1029) );
NOR2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR4_X1 U759 ( .A1(n1048), .A2(n1040), .A3(n1031), .A4(n1034), .ZN(n1024) );
INV_X1 U760 ( .A(n1049), .ZN(n1031) );
NOR2_X1 U761 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1052), .A2(n1026), .ZN(n1050) );
NOR3_X1 U763 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n1017) );
AND2_X1 U764 ( .A1(n1053), .A2(n1054), .ZN(n1019) );
NOR4_X1 U765 ( .A1(n1042), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1054) );
XNOR2_X1 U766 ( .A(n1058), .B(KEYINPUT36), .ZN(n1057) );
XNOR2_X1 U767 ( .A(n1027), .B(KEYINPUT56), .ZN(n1056) );
XOR2_X1 U768 ( .A(n1059), .B(n1060), .Z(n1055) );
XOR2_X1 U769 ( .A(KEYINPUT10), .B(G472), .Z(n1060) );
NOR4_X1 U770 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1053) );
XOR2_X1 U771 ( .A(KEYINPUT14), .B(n1026), .Z(n1064) );
NAND2_X1 U772 ( .A1(n1065), .A2(n1066), .ZN(G72) );
NAND2_X1 U773 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U774 ( .A(n1069), .B(n1070), .Z(n1067) );
NAND2_X1 U775 ( .A1(KEYINPUT63), .A2(n1071), .ZN(n1070) );
NAND2_X1 U776 ( .A1(n1072), .A2(G953), .ZN(n1065) );
XOR2_X1 U777 ( .A(n1069), .B(n1073), .Z(n1072) );
AND2_X1 U778 ( .A1(G227), .A2(G900), .ZN(n1073) );
NAND2_X1 U779 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND2_X1 U780 ( .A1(G953), .A2(n1076), .ZN(n1075) );
XOR2_X1 U781 ( .A(n1077), .B(n1078), .Z(n1074) );
XNOR2_X1 U782 ( .A(n1079), .B(n1080), .ZN(n1078) );
XOR2_X1 U783 ( .A(n1081), .B(n1082), .Z(n1077) );
NOR2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U785 ( .A(n1085), .B(KEYINPUT30), .Z(n1084) );
NAND2_X1 U786 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U787 ( .A1(n1087), .A2(n1086), .ZN(n1083) );
XNOR2_X1 U788 ( .A(KEYINPUT35), .B(n1088), .ZN(n1086) );
XNOR2_X1 U789 ( .A(G131), .B(KEYINPUT60), .ZN(n1081) );
XOR2_X1 U790 ( .A(n1089), .B(n1090), .Z(G69) );
XOR2_X1 U791 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U792 ( .A1(n1093), .A2(n1068), .ZN(n1092) );
AND2_X1 U793 ( .A1(G224), .A2(G898), .ZN(n1093) );
NOR2_X1 U794 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
XNOR2_X1 U795 ( .A(G953), .B(KEYINPUT20), .ZN(n1095) );
NOR2_X1 U796 ( .A1(n1096), .A2(n1097), .ZN(n1089) );
NOR2_X1 U797 ( .A1(n1098), .A2(n1099), .ZN(G66) );
XOR2_X1 U798 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U799 ( .A1(n1102), .A2(G217), .ZN(n1100) );
NOR2_X1 U800 ( .A1(n1098), .A2(n1103), .ZN(G63) );
XOR2_X1 U801 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U802 ( .A1(n1102), .A2(G478), .ZN(n1104) );
NOR2_X1 U803 ( .A1(n1098), .A2(n1106), .ZN(G60) );
XOR2_X1 U804 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U805 ( .A1(n1102), .A2(G475), .ZN(n1107) );
NAND2_X1 U806 ( .A1(n1109), .A2(n1110), .ZN(G6) );
NAND2_X1 U807 ( .A1(G104), .A2(n1111), .ZN(n1110) );
XOR2_X1 U808 ( .A(KEYINPUT46), .B(n1112), .Z(n1109) );
NOR2_X1 U809 ( .A1(G104), .A2(n1111), .ZN(n1112) );
NOR2_X1 U810 ( .A1(n1098), .A2(n1113), .ZN(G57) );
XOR2_X1 U811 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U812 ( .A(n1116), .B(n1117), .ZN(n1115) );
XNOR2_X1 U813 ( .A(G101), .B(KEYINPUT42), .ZN(n1117) );
XOR2_X1 U814 ( .A(n1118), .B(n1119), .Z(n1114) );
NOR3_X1 U815 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NOR2_X1 U816 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR3_X1 U817 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1121) );
INV_X1 U818 ( .A(n1124), .ZN(n1125) );
NAND2_X1 U819 ( .A1(n1128), .A2(n1129), .ZN(n1124) );
XNOR2_X1 U820 ( .A(n1130), .B(KEYINPUT8), .ZN(n1128) );
INV_X1 U821 ( .A(n1131), .ZN(n1120) );
NAND2_X1 U822 ( .A1(n1102), .A2(G472), .ZN(n1118) );
NOR2_X1 U823 ( .A1(n1132), .A2(n1133), .ZN(G54) );
XOR2_X1 U824 ( .A(KEYINPUT54), .B(n1098), .Z(n1133) );
XOR2_X1 U825 ( .A(n1134), .B(n1135), .Z(n1132) );
XOR2_X1 U826 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U827 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U828 ( .A1(KEYINPUT6), .A2(n1140), .ZN(n1139) );
XOR2_X1 U829 ( .A(n1141), .B(n1142), .Z(n1134) );
XNOR2_X1 U830 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U831 ( .A1(KEYINPUT33), .A2(n1145), .ZN(n1144) );
AND2_X1 U832 ( .A1(G469), .A2(n1102), .ZN(n1145) );
XNOR2_X1 U833 ( .A(G140), .B(KEYINPUT59), .ZN(n1141) );
NOR2_X1 U834 ( .A1(n1098), .A2(n1146), .ZN(G51) );
XOR2_X1 U835 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U836 ( .A1(n1102), .A2(n1149), .ZN(n1148) );
AND2_X1 U837 ( .A1(G902), .A2(n1021), .ZN(n1102) );
NAND2_X1 U838 ( .A1(n1094), .A2(n1150), .ZN(n1021) );
INV_X1 U839 ( .A(n1071), .ZN(n1150) );
NAND4_X1 U840 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1071) );
AND4_X1 U841 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
NAND2_X1 U842 ( .A1(n1159), .A2(n1051), .ZN(n1153) );
XOR2_X1 U843 ( .A(n1160), .B(KEYINPUT9), .Z(n1159) );
NAND2_X1 U844 ( .A1(n1161), .A2(n1162), .ZN(n1151) );
NAND2_X1 U845 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U846 ( .A1(n1049), .A2(n1165), .ZN(n1164) );
XOR2_X1 U847 ( .A(KEYINPUT48), .B(n1166), .Z(n1165) );
NAND2_X1 U848 ( .A1(n1036), .A2(n1046), .ZN(n1163) );
AND4_X1 U849 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1094) );
AND4_X1 U850 ( .A1(n1016), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1170) );
NAND3_X1 U851 ( .A1(n1046), .A2(n1044), .A3(n1174), .ZN(n1016) );
NOR2_X1 U852 ( .A1(n1175), .A2(n1176), .ZN(n1169) );
INV_X1 U853 ( .A(n1111), .ZN(n1176) );
NAND3_X1 U854 ( .A1(n1174), .A2(n1044), .A3(n1047), .ZN(n1111) );
NAND2_X1 U855 ( .A1(KEYINPUT7), .A2(n1177), .ZN(n1147) );
XOR2_X1 U856 ( .A(n1178), .B(n1097), .Z(n1177) );
NOR4_X1 U857 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT11), .A4(n1181), .ZN(n1178) );
AND3_X1 U858 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1180) );
OR2_X1 U859 ( .A1(G125), .A2(n1185), .ZN(n1184) );
NOR2_X1 U860 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
NAND2_X1 U861 ( .A1(n1186), .A2(n1185), .ZN(n1183) );
XNOR2_X1 U862 ( .A(KEYINPUT61), .B(n1187), .ZN(n1186) );
NOR2_X1 U863 ( .A1(n1068), .A2(G952), .ZN(n1098) );
XOR2_X1 U864 ( .A(G146), .B(n1188), .Z(G48) );
NOR2_X1 U865 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U866 ( .A(n1160), .B(KEYINPUT5), .Z(n1189) );
NAND3_X1 U867 ( .A1(n1166), .A2(n1047), .A3(n1191), .ZN(n1160) );
XNOR2_X1 U868 ( .A(G143), .B(n1152), .ZN(G45) );
NAND4_X1 U869 ( .A1(n1058), .A2(n1061), .A3(n1051), .A4(n1192), .ZN(n1152) );
NOR2_X1 U870 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U871 ( .A1(n1195), .A2(n1196), .ZN(G42) );
NAND2_X1 U872 ( .A1(G140), .A2(n1158), .ZN(n1196) );
XOR2_X1 U873 ( .A(n1197), .B(KEYINPUT53), .Z(n1195) );
OR2_X1 U874 ( .A1(n1158), .A2(G140), .ZN(n1197) );
NAND3_X1 U875 ( .A1(n1047), .A2(n1035), .A3(n1161), .ZN(n1158) );
XNOR2_X1 U876 ( .A(G137), .B(n1198), .ZN(G39) );
NAND4_X1 U877 ( .A1(KEYINPUT41), .A2(n1161), .A3(n1166), .A4(n1049), .ZN(n1198) );
XNOR2_X1 U878 ( .A(G134), .B(n1199), .ZN(G36) );
NAND4_X1 U879 ( .A1(KEYINPUT29), .A2(n1161), .A3(n1036), .A4(n1046), .ZN(n1199) );
XNOR2_X1 U880 ( .A(G131), .B(n1157), .ZN(G33) );
NAND3_X1 U881 ( .A1(n1047), .A2(n1036), .A3(n1161), .ZN(n1157) );
NOR3_X1 U882 ( .A1(n1026), .A2(n1027), .A3(n1194), .ZN(n1161) );
INV_X1 U883 ( .A(n1052), .ZN(n1027) );
XNOR2_X1 U884 ( .A(n1200), .B(n1201), .ZN(G30) );
NOR2_X1 U885 ( .A1(KEYINPUT21), .A2(n1156), .ZN(n1201) );
NAND4_X1 U886 ( .A1(n1191), .A2(n1166), .A3(n1046), .A4(n1051), .ZN(n1156) );
INV_X1 U887 ( .A(n1194), .ZN(n1191) );
NAND3_X1 U888 ( .A1(n1202), .A2(n1203), .A3(n1041), .ZN(n1194) );
XOR2_X1 U889 ( .A(n1175), .B(n1204), .Z(G3) );
NOR2_X1 U890 ( .A1(KEYINPUT13), .A2(n1205), .ZN(n1204) );
AND3_X1 U891 ( .A1(n1049), .A2(n1174), .A3(n1036), .ZN(n1175) );
XOR2_X1 U892 ( .A(n1155), .B(n1206), .Z(G27) );
NAND2_X1 U893 ( .A1(KEYINPUT50), .A2(G125), .ZN(n1206) );
NAND4_X1 U894 ( .A1(n1051), .A2(n1202), .A3(n1035), .A4(n1207), .ZN(n1155) );
NOR2_X1 U895 ( .A1(n1034), .A2(n1208), .ZN(n1207) );
INV_X1 U896 ( .A(n1037), .ZN(n1034) );
NAND2_X1 U897 ( .A1(n1023), .A2(n1209), .ZN(n1202) );
NAND4_X1 U898 ( .A1(n1210), .A2(G953), .A3(n1211), .A4(n1076), .ZN(n1209) );
INV_X1 U899 ( .A(G900), .ZN(n1076) );
XOR2_X1 U900 ( .A(n1167), .B(n1212), .Z(G24) );
XNOR2_X1 U901 ( .A(G122), .B(KEYINPUT23), .ZN(n1212) );
NAND4_X1 U902 ( .A1(n1213), .A2(n1044), .A3(n1058), .A4(n1061), .ZN(n1167) );
INV_X1 U903 ( .A(n1040), .ZN(n1044) );
NAND2_X1 U904 ( .A1(n1214), .A2(n1215), .ZN(n1040) );
XNOR2_X1 U905 ( .A(G119), .B(n1168), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1213), .A2(n1049), .A3(n1166), .ZN(n1168) );
AND2_X1 U907 ( .A1(n1216), .A2(n1063), .ZN(n1166) );
XNOR2_X1 U908 ( .A(G116), .B(n1173), .ZN(G18) );
NAND3_X1 U909 ( .A1(n1213), .A2(n1046), .A3(n1036), .ZN(n1173) );
NOR2_X1 U910 ( .A1(n1061), .A2(n1217), .ZN(n1046) );
XNOR2_X1 U911 ( .A(G113), .B(n1172), .ZN(G15) );
NAND3_X1 U912 ( .A1(n1036), .A2(n1213), .A3(n1047), .ZN(n1172) );
INV_X1 U913 ( .A(n1208), .ZN(n1047) );
NAND2_X1 U914 ( .A1(n1217), .A2(n1061), .ZN(n1208) );
INV_X1 U915 ( .A(n1058), .ZN(n1217) );
AND2_X1 U916 ( .A1(n1037), .A2(n1218), .ZN(n1213) );
NOR2_X1 U917 ( .A1(n1041), .A2(n1042), .ZN(n1037) );
INV_X1 U918 ( .A(n1203), .ZN(n1042) );
INV_X1 U919 ( .A(n1193), .ZN(n1036) );
NAND2_X1 U920 ( .A1(n1216), .A2(n1214), .ZN(n1193) );
INV_X1 U921 ( .A(n1063), .ZN(n1214) );
XOR2_X1 U922 ( .A(n1219), .B(KEYINPUT27), .Z(n1216) );
XNOR2_X1 U923 ( .A(G110), .B(n1171), .ZN(G12) );
NAND3_X1 U924 ( .A1(n1035), .A2(n1174), .A3(n1049), .ZN(n1171) );
NOR2_X1 U925 ( .A1(n1058), .A2(n1061), .ZN(n1049) );
XNOR2_X1 U926 ( .A(n1220), .B(G475), .ZN(n1061) );
NAND2_X1 U927 ( .A1(n1108), .A2(n1221), .ZN(n1220) );
XOR2_X1 U928 ( .A(n1222), .B(n1223), .Z(n1108) );
XNOR2_X1 U929 ( .A(n1224), .B(n1225), .ZN(n1223) );
NOR2_X1 U930 ( .A1(KEYINPUT17), .A2(n1226), .ZN(n1225) );
NAND2_X1 U931 ( .A1(n1227), .A2(KEYINPUT34), .ZN(n1224) );
XOR2_X1 U932 ( .A(n1228), .B(G131), .Z(n1227) );
NAND2_X1 U933 ( .A1(n1229), .A2(KEYINPUT39), .ZN(n1228) );
XNOR2_X1 U934 ( .A(n1230), .B(n1231), .ZN(n1229) );
NAND3_X1 U935 ( .A1(n1232), .A2(n1068), .A3(G214), .ZN(n1230) );
XOR2_X1 U936 ( .A(n1233), .B(n1234), .Z(n1222) );
NOR2_X1 U937 ( .A1(KEYINPUT58), .A2(n1235), .ZN(n1234) );
XOR2_X1 U938 ( .A(G104), .B(n1236), .Z(n1235) );
XNOR2_X1 U939 ( .A(G146), .B(G125), .ZN(n1233) );
XNOR2_X1 U940 ( .A(n1237), .B(G478), .ZN(n1058) );
NAND2_X1 U941 ( .A1(n1105), .A2(n1221), .ZN(n1237) );
XOR2_X1 U942 ( .A(n1238), .B(n1239), .Z(n1105) );
XOR2_X1 U943 ( .A(n1240), .B(n1241), .Z(n1239) );
NAND2_X1 U944 ( .A1(G217), .A2(n1242), .ZN(n1241) );
NAND2_X1 U945 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
NAND2_X1 U946 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U947 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U948 ( .A1(KEYINPUT22), .A2(n1087), .ZN(n1248) );
INV_X1 U949 ( .A(KEYINPUT62), .ZN(n1247) );
NAND2_X1 U950 ( .A1(G134), .A2(n1249), .ZN(n1243) );
NAND2_X1 U951 ( .A1(KEYINPUT22), .A2(n1250), .ZN(n1249) );
OR2_X1 U952 ( .A1(n1245), .A2(KEYINPUT62), .ZN(n1250) );
XNOR2_X1 U953 ( .A(G128), .B(n1231), .ZN(n1245) );
XNOR2_X1 U954 ( .A(G107), .B(n1251), .ZN(n1238) );
XOR2_X1 U955 ( .A(G122), .B(G116), .Z(n1251) );
AND3_X1 U956 ( .A1(n1041), .A2(n1203), .A3(n1218), .ZN(n1174) );
AND2_X1 U957 ( .A1(n1051), .A2(n1252), .ZN(n1218) );
NAND2_X1 U958 ( .A1(n1023), .A2(n1253), .ZN(n1252) );
NAND3_X1 U959 ( .A1(n1210), .A2(n1211), .A3(n1096), .ZN(n1253) );
NOR2_X1 U960 ( .A1(n1068), .A2(G898), .ZN(n1096) );
XNOR2_X1 U961 ( .A(G902), .B(KEYINPUT16), .ZN(n1210) );
NAND3_X1 U962 ( .A1(n1211), .A2(n1068), .A3(G952), .ZN(n1023) );
NAND2_X1 U963 ( .A1(G234), .A2(G237), .ZN(n1211) );
INV_X1 U964 ( .A(n1190), .ZN(n1051) );
NAND2_X1 U965 ( .A1(n1026), .A2(n1052), .ZN(n1190) );
NAND2_X1 U966 ( .A1(G214), .A2(n1254), .ZN(n1052) );
XNOR2_X1 U967 ( .A(n1255), .B(n1149), .ZN(n1026) );
AND2_X1 U968 ( .A1(G210), .A2(n1254), .ZN(n1149) );
NAND2_X1 U969 ( .A1(n1256), .A2(n1221), .ZN(n1254) );
XOR2_X1 U970 ( .A(KEYINPUT15), .B(G237), .Z(n1256) );
NAND2_X1 U971 ( .A1(n1257), .A2(n1221), .ZN(n1255) );
XOR2_X1 U972 ( .A(n1258), .B(n1097), .Z(n1257) );
XNOR2_X1 U973 ( .A(n1259), .B(n1260), .ZN(n1097) );
XOR2_X1 U974 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U975 ( .A(n1263), .B(n1264), .ZN(n1262) );
INV_X1 U976 ( .A(G119), .ZN(n1264) );
NAND2_X1 U977 ( .A1(KEYINPUT2), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U978 ( .A(KEYINPUT47), .B(KEYINPUT0), .ZN(n1261) );
XOR2_X1 U979 ( .A(n1136), .B(n1266), .Z(n1259) );
XOR2_X1 U980 ( .A(n1267), .B(n1236), .Z(n1266) );
XOR2_X1 U981 ( .A(G113), .B(G122), .Z(n1236) );
NOR2_X1 U982 ( .A1(G116), .A2(KEYINPUT32), .ZN(n1267) );
XNOR2_X1 U983 ( .A(G110), .B(n1268), .ZN(n1136) );
NAND3_X1 U984 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1258) );
INV_X1 U985 ( .A(n1181), .ZN(n1271) );
NOR3_X1 U986 ( .A1(n1182), .A2(G125), .A3(n1185), .ZN(n1181) );
NAND2_X1 U987 ( .A1(n1272), .A2(G125), .ZN(n1270) );
XOR2_X1 U988 ( .A(n1185), .B(n1182), .Z(n1272) );
NAND3_X1 U989 ( .A1(n1182), .A2(n1185), .A3(n1187), .ZN(n1269) );
INV_X1 U990 ( .A(G125), .ZN(n1187) );
AND2_X1 U991 ( .A1(G224), .A2(n1068), .ZN(n1182) );
NAND2_X1 U992 ( .A1(G221), .A2(n1273), .ZN(n1203) );
NAND2_X1 U993 ( .A1(G234), .A2(n1221), .ZN(n1273) );
XOR2_X1 U994 ( .A(n1062), .B(KEYINPUT38), .Z(n1041) );
XNOR2_X1 U995 ( .A(n1274), .B(G469), .ZN(n1062) );
NAND3_X1 U996 ( .A1(n1275), .A2(n1221), .A3(n1276), .ZN(n1274) );
NAND2_X1 U997 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U998 ( .A1(KEYINPUT43), .A2(n1279), .ZN(n1278) );
XOR2_X1 U999 ( .A(n1280), .B(n1281), .Z(n1277) );
NOR2_X1 U1000 ( .A1(KEYINPUT12), .A2(n1282), .ZN(n1280) );
NAND3_X1 U1001 ( .A1(n1283), .A2(n1279), .A3(KEYINPUT43), .ZN(n1275) );
XNOR2_X1 U1002 ( .A(n1226), .B(G110), .ZN(n1279) );
INV_X1 U1003 ( .A(G140), .ZN(n1226) );
XOR2_X1 U1004 ( .A(n1284), .B(n1281), .Z(n1283) );
XNOR2_X1 U1005 ( .A(n1285), .B(n1286), .ZN(n1281) );
XNOR2_X1 U1006 ( .A(n1140), .B(n1268), .ZN(n1286) );
XNOR2_X1 U1007 ( .A(n1205), .B(G104), .ZN(n1268) );
INV_X1 U1008 ( .A(G101), .ZN(n1205) );
INV_X1 U1009 ( .A(n1080), .ZN(n1140) );
XNOR2_X1 U1010 ( .A(n1287), .B(n1288), .ZN(n1080) );
XNOR2_X1 U1011 ( .A(G143), .B(KEYINPUT49), .ZN(n1287) );
XOR2_X1 U1012 ( .A(n1138), .B(KEYINPUT24), .Z(n1285) );
XNOR2_X1 U1013 ( .A(n1289), .B(n1290), .ZN(n1138) );
XNOR2_X1 U1014 ( .A(KEYINPUT40), .B(n1265), .ZN(n1290) );
INV_X1 U1015 ( .A(G107), .ZN(n1265) );
NOR2_X1 U1016 ( .A1(n1143), .A2(KEYINPUT12), .ZN(n1284) );
INV_X1 U1017 ( .A(n1282), .ZN(n1143) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1068), .ZN(n1282) );
AND2_X1 U1019 ( .A1(n1215), .A2(n1063), .ZN(n1035) );
NAND3_X1 U1020 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1063) );
OR2_X1 U1021 ( .A1(n1294), .A2(n1101), .ZN(n1293) );
NAND3_X1 U1022 ( .A1(n1101), .A2(n1294), .A3(n1221), .ZN(n1292) );
NAND2_X1 U1023 ( .A1(G217), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1024 ( .A(n1296), .B(n1297), .Z(n1101) );
XOR2_X1 U1025 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U1026 ( .A(G119), .B(n1300), .ZN(n1299) );
NOR2_X1 U1027 ( .A1(G110), .A2(KEYINPUT18), .ZN(n1300) );
XNOR2_X1 U1028 ( .A(G137), .B(KEYINPUT37), .ZN(n1298) );
XOR2_X1 U1029 ( .A(n1301), .B(n1079), .Z(n1296) );
XOR2_X1 U1030 ( .A(G140), .B(G125), .Z(n1079) );
XOR2_X1 U1031 ( .A(n1302), .B(n1288), .Z(n1301) );
XNOR2_X1 U1032 ( .A(n1200), .B(G146), .ZN(n1288) );
NAND2_X1 U1033 ( .A1(n1242), .A2(G221), .ZN(n1302) );
NOR2_X1 U1034 ( .A1(n1295), .A2(G953), .ZN(n1242) );
INV_X1 U1035 ( .A(G234), .ZN(n1295) );
NAND2_X1 U1036 ( .A1(G217), .A2(G902), .ZN(n1291) );
XOR2_X1 U1037 ( .A(n1219), .B(KEYINPUT44), .Z(n1215) );
XOR2_X1 U1038 ( .A(n1059), .B(n1303), .Z(n1219) );
NOR2_X1 U1039 ( .A1(KEYINPUT31), .A2(n1304), .ZN(n1303) );
XOR2_X1 U1040 ( .A(KEYINPUT3), .B(G472), .Z(n1304) );
NAND2_X1 U1041 ( .A1(n1305), .A2(n1221), .ZN(n1059) );
INV_X1 U1042 ( .A(G902), .ZN(n1221) );
XOR2_X1 U1043 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1044 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U1045 ( .A1(KEYINPUT26), .A2(n1116), .ZN(n1309) );
AND3_X1 U1046 ( .A1(n1232), .A2(n1068), .A3(G210), .ZN(n1116) );
INV_X1 U1047 ( .A(G953), .ZN(n1068) );
XOR2_X1 U1048 ( .A(G237), .B(KEYINPUT52), .Z(n1232) );
NAND3_X1 U1049 ( .A1(n1310), .A2(n1311), .A3(n1131), .ZN(n1308) );
NAND2_X1 U1050 ( .A1(n1126), .A2(n1127), .ZN(n1131) );
NOR2_X1 U1051 ( .A1(n1130), .A2(n1129), .ZN(n1126) );
NAND2_X1 U1052 ( .A1(n1312), .A2(n1129), .ZN(n1311) );
INV_X1 U1053 ( .A(n1289), .ZN(n1129) );
XNOR2_X1 U1054 ( .A(n1130), .B(n1127), .ZN(n1312) );
NAND3_X1 U1055 ( .A1(n1130), .A2(n1123), .A3(n1289), .ZN(n1310) );
XNOR2_X1 U1056 ( .A(n1313), .B(G131), .ZN(n1289) );
NAND3_X1 U1057 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1313) );
NAND2_X1 U1058 ( .A1(G137), .A2(n1087), .ZN(n1316) );
INV_X1 U1059 ( .A(G134), .ZN(n1087) );
NAND2_X1 U1060 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
INV_X1 U1061 ( .A(KEYINPUT1), .ZN(n1318) );
NAND2_X1 U1062 ( .A1(n1319), .A2(n1088), .ZN(n1317) );
XNOR2_X1 U1063 ( .A(KEYINPUT28), .B(G134), .ZN(n1319) );
NAND2_X1 U1064 ( .A1(KEYINPUT1), .A2(n1320), .ZN(n1314) );
NAND2_X1 U1065 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR2_X1 U1066 ( .A1(G134), .A2(KEYINPUT28), .ZN(n1322) );
NAND3_X1 U1067 ( .A1(G134), .A2(n1088), .A3(KEYINPUT28), .ZN(n1321) );
INV_X1 U1068 ( .A(G137), .ZN(n1088) );
INV_X1 U1069 ( .A(n1127), .ZN(n1123) );
XNOR2_X1 U1070 ( .A(n1323), .B(n1324), .ZN(n1127) );
NOR2_X1 U1071 ( .A1(KEYINPUT57), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1072 ( .A(G113), .B(KEYINPUT25), .ZN(n1325) );
XNOR2_X1 U1073 ( .A(G116), .B(G119), .ZN(n1323) );
XNOR2_X1 U1074 ( .A(n1185), .B(KEYINPUT19), .ZN(n1130) );
NAND2_X1 U1075 ( .A1(n1326), .A2(n1327), .ZN(n1185) );
NAND2_X1 U1076 ( .A1(n1328), .A2(n1200), .ZN(n1327) );
XOR2_X1 U1077 ( .A(n1329), .B(KEYINPUT55), .Z(n1326) );
OR2_X1 U1078 ( .A1(n1200), .A2(n1328), .ZN(n1329) );
XNOR2_X1 U1079 ( .A(n1330), .B(G146), .ZN(n1328) );
NAND2_X1 U1080 ( .A1(KEYINPUT51), .A2(n1231), .ZN(n1330) );
INV_X1 U1081 ( .A(G143), .ZN(n1231) );
INV_X1 U1082 ( .A(G128), .ZN(n1200) );
XNOR2_X1 U1083 ( .A(G101), .B(KEYINPUT45), .ZN(n1306) );
endmodule


