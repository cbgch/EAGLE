//Key = 0010100001010110010001011001010010101010010011000011110100010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339;

XNOR2_X1 U735 ( .A(G107), .B(n1017), .ZN(G9) );
NOR2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR4_X1 U737 ( .A1(G953), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1019) );
NOR2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U739 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR3_X1 U740 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NOR3_X1 U741 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NOR2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
XNOR2_X1 U745 ( .A(KEYINPUT45), .B(n1039), .ZN(n1038) );
XNOR2_X1 U746 ( .A(n1040), .B(KEYINPUT60), .ZN(n1037) );
NOR2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1028) );
NOR3_X1 U750 ( .A1(n1042), .A2(n1047), .A3(n1048), .ZN(n1046) );
AND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U752 ( .A(n1051), .ZN(n1027) );
NOR3_X1 U753 ( .A1(n1042), .A2(n1047), .A3(n1052), .ZN(n1025) );
NOR2_X1 U754 ( .A1(n1053), .A2(n1034), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1030), .ZN(n1053) );
INV_X1 U756 ( .A(n1045), .ZN(n1030) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U758 ( .A1(KEYINPUT57), .A2(n1057), .ZN(n1055) );
AND2_X1 U759 ( .A1(n1058), .A2(n1034), .ZN(n1047) );
INV_X1 U760 ( .A(n1059), .ZN(n1034) );
NAND3_X1 U761 ( .A1(n1045), .A2(n1060), .A3(KEYINPUT57), .ZN(n1058) );
NOR3_X1 U762 ( .A1(n1020), .A2(G953), .A3(G952), .ZN(n1018) );
AND4_X1 U763 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1020) );
NOR4_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
XNOR2_X1 U765 ( .A(n1069), .B(n1070), .ZN(n1068) );
XNOR2_X1 U766 ( .A(n1071), .B(n1072), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1073), .B(KEYINPUT58), .Z(n1072) );
NAND3_X1 U768 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1065) );
XOR2_X1 U769 ( .A(n1077), .B(KEYINPUT26), .Z(n1076) );
OR2_X1 U770 ( .A1(n1078), .A2(KEYINPUT9), .ZN(n1075) );
NAND3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(KEYINPUT9), .ZN(n1074) );
NOR3_X1 U772 ( .A1(n1050), .A2(n1080), .A3(n1081), .ZN(n1063) );
XOR2_X1 U773 ( .A(n1082), .B(n1083), .Z(G72) );
NOR2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
OR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U779 ( .A(KEYINPUT44), .B(n1094), .Z(n1088) );
NOR3_X1 U780 ( .A1(n1095), .A2(n1093), .A3(n1092), .ZN(n1094) );
XNOR2_X1 U781 ( .A(n1096), .B(n1097), .ZN(n1092) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(n1097) );
XNOR2_X1 U783 ( .A(G140), .B(n1100), .ZN(n1099) );
NAND2_X1 U784 ( .A1(KEYINPUT38), .A2(G131), .ZN(n1098) );
XNOR2_X1 U785 ( .A(n1101), .B(n1102), .ZN(n1096) );
XOR2_X1 U786 ( .A(KEYINPUT15), .B(n1090), .Z(n1095) );
AND2_X1 U787 ( .A1(n1085), .A2(n1103), .ZN(n1090) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(G69) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U791 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR3_X1 U792 ( .A1(n1112), .A2(KEYINPUT47), .A3(G953), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1115), .A2(n1085), .ZN(n1104) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XNOR2_X1 U797 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR2_X1 U798 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U799 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U801 ( .A1(n1069), .A2(n1123), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1127), .ZN(G60) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U804 ( .A1(n1130), .A2(n1123), .ZN(n1129) );
NOR2_X1 U805 ( .A1(KEYINPUT8), .A2(n1131), .ZN(n1128) );
XNOR2_X1 U806 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U807 ( .A1(n1118), .A2(n1133), .ZN(G57) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U809 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U810 ( .A1(KEYINPUT10), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U811 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR2_X1 U812 ( .A1(n1141), .A2(n1123), .ZN(n1140) );
NOR2_X1 U813 ( .A1(G101), .A2(KEYINPUT20), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1118), .A2(n1142), .ZN(G54) );
XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U816 ( .A(n1145), .B(n1146), .ZN(n1144) );
XNOR2_X1 U817 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1143) );
XOR2_X1 U819 ( .A(KEYINPUT0), .B(n1151), .Z(n1150) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1123), .ZN(n1149) );
INV_X1 U821 ( .A(G469), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1118), .A2(n1153), .ZN(G51) );
XOR2_X1 U823 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1123), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1157), .A2(n1022), .ZN(n1123) );
OR3_X1 U826 ( .A1(n1103), .A2(n1114), .A3(n1158), .ZN(n1022) );
XOR2_X1 U827 ( .A(n1113), .B(KEYINPUT12), .Z(n1158) );
AND2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(n1113) );
XNOR2_X1 U829 ( .A(n1161), .B(KEYINPUT52), .ZN(n1159) );
NAND4_X1 U830 ( .A1(n1132), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1114) );
AND4_X1 U831 ( .A1(n1165), .A2(n1017), .A3(n1166), .A4(n1167), .ZN(n1164) );
NAND4_X1 U832 ( .A1(n1168), .A2(n1060), .A3(n1160), .A4(n1059), .ZN(n1017) );
NAND2_X1 U833 ( .A1(n1169), .A2(n1160), .ZN(n1163) );
NAND4_X1 U834 ( .A1(n1056), .A2(n1168), .A3(n1160), .A4(n1059), .ZN(n1132) );
NAND4_X1 U835 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1103) );
NOR4_X1 U836 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NOR2_X1 U837 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
NAND2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1171) );
NAND2_X1 U839 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND4_X1 U840 ( .A1(KEYINPUT39), .A2(n1184), .A3(n1044), .A4(n1185), .ZN(n1183) );
INV_X1 U841 ( .A(n1056), .ZN(n1185) );
XNOR2_X1 U842 ( .A(KEYINPUT50), .B(n1186), .ZN(n1182) );
OR2_X1 U843 ( .A1(n1187), .A2(KEYINPUT39), .ZN(n1170) );
XNOR2_X1 U844 ( .A(KEYINPUT37), .B(n1188), .ZN(n1157) );
NOR2_X1 U845 ( .A1(n1085), .A2(G952), .ZN(n1118) );
XOR2_X1 U846 ( .A(G146), .B(n1179), .Z(G48) );
AND3_X1 U847 ( .A1(n1184), .A2(n1056), .A3(n1189), .ZN(n1179) );
XOR2_X1 U848 ( .A(n1190), .B(n1177), .Z(G45) );
AND3_X1 U849 ( .A1(n1043), .A2(n1184), .A3(n1191), .ZN(n1177) );
NAND2_X1 U850 ( .A1(KEYINPUT27), .A2(n1192), .ZN(n1190) );
XOR2_X1 U851 ( .A(n1187), .B(n1193), .Z(G42) );
XNOR2_X1 U852 ( .A(KEYINPUT55), .B(n1194), .ZN(n1193) );
NAND4_X1 U853 ( .A1(n1184), .A2(n1044), .A3(n1056), .A4(n1180), .ZN(n1187) );
XOR2_X1 U854 ( .A(G137), .B(n1195), .Z(G39) );
NOR2_X1 U855 ( .A1(n1042), .A2(n1186), .ZN(n1195) );
NAND4_X1 U856 ( .A1(n1051), .A2(n1184), .A3(n1196), .A4(n1067), .ZN(n1186) );
INV_X1 U857 ( .A(n1180), .ZN(n1042) );
XOR2_X1 U858 ( .A(G134), .B(n1178), .Z(G36) );
AND4_X1 U859 ( .A1(n1043), .A2(n1184), .A3(n1060), .A4(n1180), .ZN(n1178) );
XOR2_X1 U860 ( .A(n1176), .B(n1197), .Z(G33) );
NOR2_X1 U861 ( .A1(KEYINPUT3), .A2(n1198), .ZN(n1197) );
XOR2_X1 U862 ( .A(KEYINPUT32), .B(G131), .Z(n1198) );
AND4_X1 U863 ( .A1(n1043), .A2(n1184), .A3(n1056), .A4(n1180), .ZN(n1176) );
NAND2_X1 U864 ( .A1(n1199), .A2(n1200), .ZN(n1180) );
NAND3_X1 U865 ( .A1(n1040), .A2(n1039), .A3(n1201), .ZN(n1200) );
INV_X1 U866 ( .A(KEYINPUT60), .ZN(n1201) );
NAND2_X1 U867 ( .A1(KEYINPUT60), .A2(n1036), .ZN(n1199) );
XNOR2_X1 U868 ( .A(n1202), .B(n1175), .ZN(G30) );
AND3_X1 U869 ( .A1(n1184), .A2(n1060), .A3(n1189), .ZN(n1175) );
AND3_X1 U870 ( .A1(n1049), .A2(n1203), .A3(n1204), .ZN(n1184) );
XNOR2_X1 U871 ( .A(G101), .B(n1205), .ZN(G3) );
NAND3_X1 U872 ( .A1(n1160), .A2(n1206), .A3(KEYINPUT53), .ZN(n1205) );
XOR2_X1 U873 ( .A(KEYINPUT6), .B(n1169), .Z(n1206) );
AND3_X1 U874 ( .A1(n1043), .A2(n1168), .A3(n1051), .ZN(n1169) );
XOR2_X1 U875 ( .A(G125), .B(n1174), .Z(G27) );
AND4_X1 U876 ( .A1(n1036), .A2(n1204), .A3(n1056), .A4(n1207), .ZN(n1174) );
AND2_X1 U877 ( .A1(n1045), .A2(n1044), .ZN(n1207) );
NAND2_X1 U878 ( .A1(n1024), .A2(n1208), .ZN(n1204) );
NAND3_X1 U879 ( .A1(G902), .A2(n1209), .A3(n1093), .ZN(n1208) );
AND2_X1 U880 ( .A1(n1210), .A2(n1087), .ZN(n1093) );
INV_X1 U881 ( .A(G900), .ZN(n1087) );
XOR2_X1 U882 ( .A(G122), .B(n1211), .Z(G24) );
NOR2_X1 U883 ( .A1(KEYINPUT49), .A2(n1166), .ZN(n1211) );
NAND3_X1 U884 ( .A1(n1191), .A2(n1059), .A3(n1212), .ZN(n1166) );
NOR2_X1 U885 ( .A1(n1067), .A2(n1196), .ZN(n1059) );
AND3_X1 U886 ( .A1(n1213), .A2(n1214), .A3(n1036), .ZN(n1191) );
XNOR2_X1 U887 ( .A(G119), .B(n1215), .ZN(G21) );
NAND2_X1 U888 ( .A1(KEYINPUT4), .A2(n1216), .ZN(n1215) );
INV_X1 U889 ( .A(n1165), .ZN(n1216) );
NAND3_X1 U890 ( .A1(n1051), .A2(n1189), .A3(n1212), .ZN(n1165) );
AND3_X1 U891 ( .A1(n1036), .A2(n1067), .A3(n1196), .ZN(n1189) );
INV_X1 U892 ( .A(n1217), .ZN(n1196) );
XOR2_X1 U893 ( .A(G116), .B(n1218), .Z(G18) );
NOR2_X1 U894 ( .A1(KEYINPUT25), .A2(n1162), .ZN(n1218) );
NAND4_X1 U895 ( .A1(n1212), .A2(n1043), .A3(n1060), .A4(n1036), .ZN(n1162) );
INV_X1 U896 ( .A(n1057), .ZN(n1060) );
NAND2_X1 U897 ( .A1(n1061), .A2(n1214), .ZN(n1057) );
XNOR2_X1 U898 ( .A(G113), .B(n1167), .ZN(G15) );
NAND4_X1 U899 ( .A1(n1212), .A2(n1043), .A3(n1160), .A4(n1056), .ZN(n1167) );
NOR2_X1 U900 ( .A1(n1214), .A2(n1061), .ZN(n1056) );
INV_X1 U901 ( .A(n1213), .ZN(n1061) );
AND2_X1 U902 ( .A1(n1217), .A2(n1067), .ZN(n1043) );
AND2_X1 U903 ( .A1(n1045), .A2(n1219), .ZN(n1212) );
NOR2_X1 U904 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
INV_X1 U905 ( .A(n1203), .ZN(n1050) );
NAND2_X1 U906 ( .A1(n1220), .A2(n1221), .ZN(G12) );
NAND2_X1 U907 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U908 ( .A(KEYINPUT36), .B(n1224), .Z(n1220) );
NOR2_X1 U909 ( .A1(n1222), .A2(n1223), .ZN(n1224) );
INV_X1 U910 ( .A(G110), .ZN(n1223) );
AND2_X1 U911 ( .A1(n1161), .A2(n1225), .ZN(n1222) );
XNOR2_X1 U912 ( .A(KEYINPUT14), .B(n1160), .ZN(n1225) );
XNOR2_X1 U913 ( .A(n1036), .B(KEYINPUT2), .ZN(n1160) );
NOR2_X1 U914 ( .A1(n1080), .A2(n1040), .ZN(n1036) );
NOR2_X1 U915 ( .A1(n1081), .A2(n1226), .ZN(n1040) );
AND2_X1 U916 ( .A1(n1078), .A2(n1079), .ZN(n1226) );
NOR2_X1 U917 ( .A1(n1079), .A2(n1078), .ZN(n1081) );
INV_X1 U918 ( .A(n1156), .ZN(n1078) );
NAND2_X1 U919 ( .A1(G210), .A2(n1227), .ZN(n1156) );
OR2_X1 U920 ( .A1(n1155), .A2(n1228), .ZN(n1079) );
XNOR2_X1 U921 ( .A(n1229), .B(n1230), .ZN(n1155) );
XNOR2_X1 U922 ( .A(n1231), .B(n1232), .ZN(n1230) );
XOR2_X1 U923 ( .A(n1233), .B(n1234), .Z(n1229) );
NOR2_X1 U924 ( .A1(G953), .A2(n1116), .ZN(n1234) );
INV_X1 U925 ( .A(G224), .ZN(n1116) );
XOR2_X1 U926 ( .A(n1235), .B(n1236), .Z(n1233) );
NAND3_X1 U927 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1235) );
OR2_X1 U928 ( .A1(n1240), .A2(KEYINPUT13), .ZN(n1239) );
INV_X1 U929 ( .A(n1110), .ZN(n1240) );
NAND3_X1 U930 ( .A1(KEYINPUT13), .A2(n1241), .A3(n1111), .ZN(n1238) );
OR2_X1 U931 ( .A1(n1111), .A2(n1241), .ZN(n1237) );
NOR2_X1 U932 ( .A1(KEYINPUT33), .A2(n1110), .ZN(n1241) );
XOR2_X1 U933 ( .A(G110), .B(G122), .Z(n1110) );
XOR2_X1 U934 ( .A(n1242), .B(n1243), .Z(n1111) );
XNOR2_X1 U935 ( .A(n1244), .B(G104), .ZN(n1243) );
XOR2_X1 U936 ( .A(n1245), .B(G101), .Z(n1242) );
NAND3_X1 U937 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1245) );
NAND2_X1 U938 ( .A1(KEYINPUT31), .A2(n1249), .ZN(n1248) );
OR3_X1 U939 ( .A1(n1249), .A2(KEYINPUT31), .A3(G113), .ZN(n1247) );
NAND2_X1 U940 ( .A1(G113), .A2(n1250), .ZN(n1246) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U942 ( .A(KEYINPUT31), .ZN(n1252) );
XOR2_X1 U943 ( .A(KEYINPUT23), .B(n1249), .Z(n1251) );
XOR2_X1 U944 ( .A(n1253), .B(n1254), .Z(n1249) );
NOR2_X1 U945 ( .A1(KEYINPUT22), .A2(n1255), .ZN(n1254) );
INV_X1 U946 ( .A(n1039), .ZN(n1080) );
NAND2_X1 U947 ( .A1(n1256), .A2(G214), .ZN(n1039) );
XOR2_X1 U948 ( .A(n1227), .B(KEYINPUT16), .Z(n1256) );
NAND2_X1 U949 ( .A1(n1257), .A2(n1188), .ZN(n1227) );
INV_X1 U950 ( .A(G237), .ZN(n1257) );
AND3_X1 U951 ( .A1(n1044), .A2(n1168), .A3(n1051), .ZN(n1161) );
NOR2_X1 U952 ( .A1(n1214), .A2(n1213), .ZN(n1051) );
XOR2_X1 U953 ( .A(n1258), .B(n1130), .Z(n1213) );
INV_X1 U954 ( .A(G475), .ZN(n1130) );
NAND2_X1 U955 ( .A1(n1131), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U956 ( .A(n1260), .B(n1261), .ZN(n1131) );
XOR2_X1 U957 ( .A(G113), .B(n1262), .Z(n1261) );
XNOR2_X1 U958 ( .A(n1194), .B(G122), .ZN(n1262) );
XOR2_X1 U959 ( .A(n1263), .B(n1264), .Z(n1260) );
XOR2_X1 U960 ( .A(n1265), .B(G104), .Z(n1263) );
NAND2_X1 U961 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U962 ( .A1(n1268), .A2(G131), .ZN(n1267) );
XOR2_X1 U963 ( .A(n1269), .B(KEYINPUT5), .Z(n1266) );
OR2_X1 U964 ( .A1(n1268), .A2(G131), .ZN(n1269) );
XOR2_X1 U965 ( .A(n1270), .B(G143), .Z(n1268) );
NAND3_X1 U966 ( .A1(n1271), .A2(n1272), .A3(G214), .ZN(n1270) );
XNOR2_X1 U967 ( .A(KEYINPUT61), .B(n1085), .ZN(n1272) );
NAND2_X1 U968 ( .A1(n1273), .A2(n1274), .ZN(n1214) );
NAND2_X1 U969 ( .A1(n1070), .A2(n1275), .ZN(n1274) );
XOR2_X1 U970 ( .A(KEYINPUT63), .B(n1276), .Z(n1273) );
NOR2_X1 U971 ( .A1(n1070), .A2(n1275), .ZN(n1276) );
XNOR2_X1 U972 ( .A(KEYINPUT29), .B(n1069), .ZN(n1275) );
INV_X1 U973 ( .A(G478), .ZN(n1069) );
NOR2_X1 U974 ( .A1(n1125), .A2(n1228), .ZN(n1070) );
INV_X1 U975 ( .A(n1259), .ZN(n1228) );
XOR2_X1 U976 ( .A(n1277), .B(n1278), .Z(n1125) );
XOR2_X1 U977 ( .A(G116), .B(n1279), .Z(n1278) );
XOR2_X1 U978 ( .A(KEYINPUT54), .B(G122), .Z(n1279) );
XOR2_X1 U979 ( .A(n1280), .B(n1281), .Z(n1277) );
AND2_X1 U980 ( .A1(n1282), .A2(G217), .ZN(n1281) );
XNOR2_X1 U981 ( .A(G107), .B(n1283), .ZN(n1280) );
NOR2_X1 U982 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U983 ( .A(KEYINPUT56), .B(n1286), .Z(n1285) );
NOR2_X1 U984 ( .A1(G134), .A2(n1287), .ZN(n1286) );
AND2_X1 U985 ( .A1(n1287), .A2(G134), .ZN(n1284) );
NAND2_X1 U986 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U987 ( .A1(n1290), .A2(n1192), .ZN(n1289) );
NAND2_X1 U988 ( .A1(G143), .A2(n1291), .ZN(n1288) );
NAND2_X1 U989 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U990 ( .A1(KEYINPUT43), .A2(G128), .ZN(n1293) );
OR2_X1 U991 ( .A1(n1290), .A2(KEYINPUT43), .ZN(n1292) );
AND2_X1 U992 ( .A1(KEYINPUT24), .A2(G128), .ZN(n1290) );
AND3_X1 U993 ( .A1(n1049), .A2(n1203), .A3(n1219), .ZN(n1168) );
NAND2_X1 U994 ( .A1(n1024), .A2(n1294), .ZN(n1219) );
NAND3_X1 U995 ( .A1(G902), .A2(n1209), .A3(n1108), .ZN(n1294) );
AND2_X1 U996 ( .A1(n1210), .A2(n1117), .ZN(n1108) );
INV_X1 U997 ( .A(G898), .ZN(n1117) );
XNOR2_X1 U998 ( .A(KEYINPUT35), .B(n1085), .ZN(n1210) );
NAND3_X1 U999 ( .A1(n1209), .A2(n1085), .A3(G952), .ZN(n1024) );
NAND2_X1 U1000 ( .A1(G237), .A2(G234), .ZN(n1209) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1295), .ZN(n1203) );
NAND2_X1 U1002 ( .A1(n1077), .A2(n1062), .ZN(n1049) );
NAND2_X1 U1003 ( .A1(G469), .A2(n1296), .ZN(n1062) );
OR2_X1 U1004 ( .A1(n1296), .A2(G469), .ZN(n1077) );
NAND2_X1 U1005 ( .A1(n1297), .A2(n1259), .ZN(n1296) );
XOR2_X1 U1006 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U1007 ( .A(KEYINPUT17), .B(n1300), .Z(n1299) );
NOR3_X1 U1008 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
AND2_X1 U1009 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NOR3_X1 U1010 ( .A1(n1305), .A2(KEYINPUT19), .A3(n1304), .ZN(n1302) );
NAND2_X1 U1011 ( .A1(KEYINPUT21), .A2(n1151), .ZN(n1304) );
NOR2_X1 U1012 ( .A1(n1151), .A2(n1306), .ZN(n1301) );
INV_X1 U1013 ( .A(KEYINPUT19), .ZN(n1306) );
NOR2_X1 U1014 ( .A1(n1086), .A2(G953), .ZN(n1151) );
INV_X1 U1015 ( .A(G227), .ZN(n1086) );
NAND2_X1 U1016 ( .A1(n1307), .A2(n1308), .ZN(n1298) );
NAND2_X1 U1017 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XNOR2_X1 U1018 ( .A(n1231), .B(n1311), .ZN(n1310) );
INV_X1 U1019 ( .A(n1145), .ZN(n1311) );
XNOR2_X1 U1020 ( .A(n1312), .B(n1313), .ZN(n1309) );
INV_X1 U1021 ( .A(n1314), .ZN(n1312) );
XOR2_X1 U1022 ( .A(n1315), .B(KEYINPUT46), .Z(n1307) );
NAND2_X1 U1023 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XNOR2_X1 U1024 ( .A(n1314), .B(n1313), .ZN(n1317) );
XNOR2_X1 U1025 ( .A(n1231), .B(n1145), .ZN(n1316) );
XNOR2_X1 U1026 ( .A(n1318), .B(n1319), .ZN(n1145) );
XNOR2_X1 U1027 ( .A(n1244), .B(G101), .ZN(n1319) );
INV_X1 U1028 ( .A(G107), .ZN(n1244) );
XOR2_X1 U1029 ( .A(n1320), .B(n1100), .Z(n1318) );
NOR2_X1 U1030 ( .A1(KEYINPUT48), .A2(G128), .ZN(n1100) );
NAND2_X1 U1031 ( .A1(KEYINPUT11), .A2(G104), .ZN(n1320) );
NOR2_X1 U1032 ( .A1(n1217), .A2(n1067), .ZN(n1044) );
XOR2_X1 U1033 ( .A(n1321), .B(n1141), .Z(n1067) );
INV_X1 U1034 ( .A(G472), .ZN(n1141) );
NAND2_X1 U1035 ( .A1(n1322), .A2(n1259), .ZN(n1321) );
XNOR2_X1 U1036 ( .A(n1323), .B(n1324), .ZN(n1322) );
XNOR2_X1 U1037 ( .A(G101), .B(n1137), .ZN(n1324) );
NAND3_X1 U1038 ( .A1(n1271), .A2(n1085), .A3(G210), .ZN(n1137) );
XNOR2_X1 U1039 ( .A(G237), .B(KEYINPUT30), .ZN(n1271) );
INV_X1 U1040 ( .A(n1139), .ZN(n1323) );
XNOR2_X1 U1041 ( .A(n1325), .B(n1326), .ZN(n1139) );
XOR2_X1 U1042 ( .A(n1255), .B(n1148), .Z(n1326) );
XOR2_X1 U1043 ( .A(n1313), .B(n1102), .Z(n1148) );
XNOR2_X1 U1044 ( .A(n1314), .B(n1231), .ZN(n1102) );
XNOR2_X1 U1045 ( .A(G146), .B(n1192), .ZN(n1231) );
INV_X1 U1046 ( .A(G143), .ZN(n1192) );
XNOR2_X1 U1047 ( .A(G137), .B(G134), .ZN(n1314) );
XOR2_X1 U1048 ( .A(G131), .B(KEYINPUT40), .Z(n1313) );
XOR2_X1 U1049 ( .A(G116), .B(KEYINPUT34), .Z(n1255) );
XOR2_X1 U1050 ( .A(n1327), .B(n1328), .Z(n1325) );
NOR2_X1 U1051 ( .A1(KEYINPUT7), .A2(n1253), .ZN(n1328) );
XNOR2_X1 U1052 ( .A(G113), .B(n1236), .ZN(n1327) );
NOR2_X1 U1053 ( .A1(KEYINPUT62), .A2(n1202), .ZN(n1236) );
XNOR2_X1 U1054 ( .A(n1073), .B(n1329), .ZN(n1217) );
NOR2_X1 U1055 ( .A1(n1071), .A2(KEYINPUT42), .ZN(n1329) );
INV_X1 U1056 ( .A(n1122), .ZN(n1071) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1295), .ZN(n1122) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1188), .ZN(n1295) );
INV_X1 U1059 ( .A(G902), .ZN(n1188) );
NAND2_X1 U1060 ( .A1(n1330), .A2(n1120), .ZN(n1073) );
XNOR2_X1 U1061 ( .A(n1331), .B(n1332), .ZN(n1120) );
XNOR2_X1 U1062 ( .A(n1305), .B(n1333), .ZN(n1332) );
XNOR2_X1 U1063 ( .A(n1334), .B(n1264), .ZN(n1333) );
XNOR2_X1 U1064 ( .A(G146), .B(n1232), .ZN(n1264) );
INV_X1 U1065 ( .A(n1101), .ZN(n1232) );
XOR2_X1 U1066 ( .A(G125), .B(KEYINPUT41), .Z(n1101) );
NAND2_X1 U1067 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1068 ( .A1(n1253), .A2(n1202), .ZN(n1336) );
XOR2_X1 U1069 ( .A(n1337), .B(KEYINPUT1), .Z(n1335) );
OR2_X1 U1070 ( .A1(n1253), .A2(n1202), .ZN(n1337) );
INV_X1 U1071 ( .A(G128), .ZN(n1202) );
XOR2_X1 U1072 ( .A(G119), .B(KEYINPUT18), .Z(n1253) );
INV_X1 U1073 ( .A(n1147), .ZN(n1305) );
XNOR2_X1 U1074 ( .A(G110), .B(n1194), .ZN(n1147) );
INV_X1 U1075 ( .A(G140), .ZN(n1194) );
XOR2_X1 U1076 ( .A(n1338), .B(n1339), .Z(n1331) );
XOR2_X1 U1077 ( .A(KEYINPUT28), .B(G137), .Z(n1339) );
NAND2_X1 U1078 ( .A1(n1282), .A2(G221), .ZN(n1338) );
AND2_X1 U1079 ( .A1(G234), .A2(n1085), .ZN(n1282) );
INV_X1 U1080 ( .A(G953), .ZN(n1085) );
XNOR2_X1 U1081 ( .A(n1259), .B(KEYINPUT51), .ZN(n1330) );
XOR2_X1 U1082 ( .A(G902), .B(KEYINPUT59), .Z(n1259) );
endmodule


