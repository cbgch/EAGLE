//Key = 1011100110001011000001101100001000010111011110010100111011010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387;

XOR2_X1 U759 ( .A(G107), .B(n1043), .Z(G9) );
NOR2_X1 U760 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR3_X1 U761 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND3_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1046) );
NAND2_X1 U763 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U764 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U765 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1059) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND3_X1 U772 ( .A1(n1065), .A2(n1071), .A3(n1061), .ZN(n1054) );
NAND3_X1 U773 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NAND2_X1 U774 ( .A1(n1056), .A2(n1075), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1058), .A2(n1076), .ZN(n1072) );
NAND2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U778 ( .A(n1081), .ZN(n1052) );
AND3_X1 U779 ( .A1(n1049), .A2(n1050), .A3(n1082), .ZN(n1044) );
NAND4_X1 U780 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1049) );
NOR4_X1 U781 ( .A1(n1070), .A2(n1079), .A3(n1087), .A4(n1088), .ZN(n1086) );
XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(n1088) );
XNOR2_X1 U783 ( .A(KEYINPUT2), .B(n1091), .ZN(n1090) );
XOR2_X1 U784 ( .A(n1092), .B(n1093), .Z(n1087) );
NOR2_X1 U785 ( .A1(G469), .A2(KEYINPUT9), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1085) );
XNOR2_X1 U787 ( .A(n1096), .B(KEYINPUT63), .ZN(n1094) );
XNOR2_X1 U788 ( .A(n1097), .B(n1098), .ZN(n1083) );
NAND2_X1 U789 ( .A1(KEYINPUT15), .A2(n1099), .ZN(n1097) );
XOR2_X1 U790 ( .A(n1100), .B(n1101), .Z(G72) );
XOR2_X1 U791 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U793 ( .A(KEYINPUT16), .B(n1106), .Z(n1105) );
NOR2_X1 U794 ( .A1(G900), .A2(n1050), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1104) );
XOR2_X1 U796 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U797 ( .A1(KEYINPUT5), .A2(n1111), .ZN(n1110) );
XNOR2_X1 U798 ( .A(G140), .B(n1112), .ZN(n1111) );
NOR2_X1 U799 ( .A1(G125), .A2(KEYINPUT55), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1113), .A2(n1050), .ZN(n1102) );
XOR2_X1 U801 ( .A(n1047), .B(KEYINPUT40), .Z(n1113) );
NAND2_X1 U802 ( .A1(G953), .A2(n1114), .ZN(n1100) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND2_X1 U804 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U806 ( .A1(G953), .A2(n1119), .ZN(n1118) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1119) );
NAND2_X1 U808 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U810 ( .A1(G953), .A2(n1124), .ZN(n1123) );
INV_X1 U811 ( .A(n1117), .ZN(n1120) );
XNOR2_X1 U812 ( .A(n1125), .B(n1126), .ZN(n1117) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U814 ( .A(G953), .B(KEYINPUT43), .ZN(n1128) );
INV_X1 U815 ( .A(n1048), .ZN(n1127) );
NAND2_X1 U816 ( .A1(n1129), .A2(n1122), .ZN(n1125) );
NAND2_X1 U817 ( .A1(G953), .A2(n1130), .ZN(n1122) );
XOR2_X1 U818 ( .A(n1131), .B(n1132), .Z(n1129) );
NAND2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
NAND2_X1 U820 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U821 ( .A(KEYINPUT4), .B(n1137), .Z(n1133) );
NOR2_X1 U822 ( .A1(n1136), .A2(n1135), .ZN(n1137) );
NOR2_X1 U823 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U824 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U825 ( .A1(n1098), .A2(n1142), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1138), .A2(n1143), .ZN(G63) );
NOR2_X1 U827 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U828 ( .A(KEYINPUT33), .B(n1146), .Z(n1145) );
AND2_X1 U829 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U830 ( .A1(n1148), .A2(n1147), .ZN(n1144) );
NAND2_X1 U831 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
XOR2_X1 U832 ( .A(KEYINPUT18), .B(G478), .Z(n1150) );
NOR2_X1 U833 ( .A1(n1138), .A2(n1151), .ZN(G60) );
XOR2_X1 U834 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U835 ( .A1(n1154), .A2(KEYINPUT32), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1091), .A2(n1142), .ZN(n1154) );
XNOR2_X1 U837 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U838 ( .A1(n1138), .A2(n1156), .ZN(G57) );
XOR2_X1 U839 ( .A(n1157), .B(KEYINPUT39), .Z(n1156) );
NAND2_X1 U840 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U841 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U842 ( .A(n1162), .B(KEYINPUT13), .Z(n1158) );
OR2_X1 U843 ( .A1(n1161), .A2(n1160), .ZN(n1162) );
NAND2_X1 U844 ( .A1(n1163), .A2(n1164), .ZN(n1160) );
OR3_X1 U845 ( .A1(n1142), .A2(n1165), .A3(n1166), .ZN(n1164) );
NAND2_X1 U846 ( .A1(n1167), .A2(n1166), .ZN(n1163) );
XNOR2_X1 U847 ( .A(n1168), .B(n1169), .ZN(n1166) );
NAND2_X1 U848 ( .A1(KEYINPUT42), .A2(n1170), .ZN(n1168) );
XNOR2_X1 U849 ( .A(n1171), .B(n1172), .ZN(n1170) );
XOR2_X1 U850 ( .A(KEYINPUT3), .B(n1173), .Z(n1167) );
NOR2_X1 U851 ( .A1(n1165), .A2(n1142), .ZN(n1173) );
XNOR2_X1 U852 ( .A(n1174), .B(G101), .ZN(n1161) );
NAND2_X1 U853 ( .A1(KEYINPUT49), .A2(n1175), .ZN(n1174) );
NOR2_X1 U854 ( .A1(n1138), .A2(n1176), .ZN(G54) );
XOR2_X1 U855 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U856 ( .A(n1172), .B(n1179), .Z(n1178) );
XNOR2_X1 U857 ( .A(n1180), .B(n1181), .ZN(n1177) );
NAND2_X1 U858 ( .A1(KEYINPUT41), .A2(n1182), .ZN(n1181) );
NAND2_X1 U859 ( .A1(KEYINPUT21), .A2(n1183), .ZN(n1180) );
NAND2_X1 U860 ( .A1(n1149), .A2(G469), .ZN(n1183) );
INV_X1 U861 ( .A(n1142), .ZN(n1149) );
NOR2_X1 U862 ( .A1(n1138), .A2(n1184), .ZN(G51) );
XOR2_X1 U863 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U864 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U865 ( .A1(KEYINPUT11), .A2(n1171), .ZN(n1188) );
NOR2_X1 U866 ( .A1(n1189), .A2(n1142), .ZN(n1187) );
NAND2_X1 U867 ( .A1(G902), .A2(n1190), .ZN(n1142) );
OR2_X1 U868 ( .A1(n1048), .A2(n1047), .ZN(n1190) );
NAND4_X1 U869 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1047) );
NOR4_X1 U870 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR2_X1 U871 ( .A1(n1199), .A2(n1200), .ZN(n1193) );
NOR2_X1 U872 ( .A1(n1067), .A2(n1201), .ZN(n1200) );
NOR4_X1 U873 ( .A1(n1202), .A2(n1203), .A3(n1063), .A4(n1204), .ZN(n1199) );
XNOR2_X1 U874 ( .A(n1061), .B(KEYINPUT27), .ZN(n1202) );
NAND4_X1 U875 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1048) );
NOR4_X1 U876 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NOR3_X1 U877 ( .A1(n1073), .A2(n1213), .A3(n1064), .ZN(n1212) );
NOR3_X1 U878 ( .A1(n1063), .A2(n1214), .A3(n1215), .ZN(n1211) );
XNOR2_X1 U879 ( .A(n1216), .B(KEYINPUT58), .ZN(n1214) );
INV_X1 U880 ( .A(n1217), .ZN(n1063) );
INV_X1 U881 ( .A(n1155), .ZN(n1210) );
NAND4_X1 U882 ( .A1(n1218), .A2(n1216), .A3(n1219), .A4(n1065), .ZN(n1155) );
INV_X1 U883 ( .A(n1220), .ZN(n1209) );
NOR2_X1 U884 ( .A1(n1221), .A2(n1043), .ZN(n1207) );
AND4_X1 U885 ( .A1(n1216), .A2(n1219), .A3(n1075), .A4(n1065), .ZN(n1043) );
XOR2_X1 U886 ( .A(n1222), .B(n1223), .Z(n1185) );
XNOR2_X1 U887 ( .A(G125), .B(n1224), .ZN(n1223) );
AND2_X1 U888 ( .A1(n1225), .A2(n1082), .ZN(n1138) );
INV_X1 U889 ( .A(G952), .ZN(n1082) );
XNOR2_X1 U890 ( .A(G953), .B(KEYINPUT62), .ZN(n1225) );
XNOR2_X1 U891 ( .A(G146), .B(n1192), .ZN(G48) );
NAND3_X1 U892 ( .A1(n1218), .A2(n1226), .A3(n1227), .ZN(n1192) );
NAND3_X1 U893 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(G45) );
NAND2_X1 U894 ( .A1(KEYINPUT6), .A2(n1231), .ZN(n1230) );
NAND2_X1 U895 ( .A1(G143), .A2(n1232), .ZN(n1231) );
NAND3_X1 U896 ( .A1(n1233), .A2(n1234), .A3(G143), .ZN(n1229) );
INV_X1 U897 ( .A(KEYINPUT6), .ZN(n1234) );
NAND2_X1 U898 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
NAND3_X1 U899 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1228) );
INV_X1 U900 ( .A(KEYINPUT17), .ZN(n1236) );
INV_X1 U901 ( .A(n1232), .ZN(n1235) );
NAND2_X1 U902 ( .A1(n1238), .A2(n1226), .ZN(n1232) );
XOR2_X1 U903 ( .A(n1201), .B(KEYINPUT37), .Z(n1238) );
NAND4_X1 U904 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1201) );
XNOR2_X1 U905 ( .A(G140), .B(n1243), .ZN(G42) );
NAND4_X1 U906 ( .A1(n1061), .A2(n1240), .A3(n1217), .A4(n1218), .ZN(n1243) );
XNOR2_X1 U907 ( .A(G137), .B(n1244), .ZN(G39) );
NAND2_X1 U908 ( .A1(KEYINPUT14), .A2(n1198), .ZN(n1244) );
AND3_X1 U909 ( .A1(n1227), .A2(n1058), .A3(n1061), .ZN(n1198) );
INV_X1 U910 ( .A(n1245), .ZN(n1061) );
XOR2_X1 U911 ( .A(G134), .B(n1197), .Z(G36) );
AND2_X1 U912 ( .A1(n1246), .A2(n1075), .ZN(n1197) );
XOR2_X1 U913 ( .A(G131), .B(n1196), .Z(G33) );
AND2_X1 U914 ( .A1(n1246), .A2(n1218), .ZN(n1196) );
NOR3_X1 U915 ( .A1(n1204), .A2(n1064), .A3(n1245), .ZN(n1246) );
NAND2_X1 U916 ( .A1(n1069), .A2(n1247), .ZN(n1245) );
INV_X1 U917 ( .A(n1096), .ZN(n1069) );
XOR2_X1 U918 ( .A(n1248), .B(n1195), .Z(G30) );
AND3_X1 U919 ( .A1(n1075), .A2(n1226), .A3(n1227), .ZN(n1195) );
AND3_X1 U920 ( .A1(n1249), .A2(n1095), .A3(n1240), .ZN(n1227) );
INV_X1 U921 ( .A(n1204), .ZN(n1240) );
NAND2_X1 U922 ( .A1(n1216), .A2(n1250), .ZN(n1204) );
NAND2_X1 U923 ( .A1(KEYINPUT35), .A2(n1251), .ZN(n1248) );
XOR2_X1 U924 ( .A(G101), .B(n1221), .Z(G3) );
NOR3_X1 U925 ( .A1(n1064), .A2(n1077), .A3(n1215), .ZN(n1221) );
INV_X1 U926 ( .A(n1216), .ZN(n1077) );
XNOR2_X1 U927 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U928 ( .A1(n1252), .A2(n1217), .A3(n1226), .A4(n1250), .ZN(n1191) );
NAND2_X1 U929 ( .A1(n1081), .A2(n1253), .ZN(n1250) );
NAND4_X1 U930 ( .A1(G902), .A2(G953), .A3(n1254), .A4(n1255), .ZN(n1253) );
INV_X1 U931 ( .A(G900), .ZN(n1255) );
XNOR2_X1 U932 ( .A(G122), .B(n1220), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1239), .A2(n1056), .A3(n1256), .A4(n1219), .ZN(n1220) );
AND2_X1 U934 ( .A1(n1242), .A2(n1065), .ZN(n1256) );
NOR2_X1 U935 ( .A1(n1095), .A2(n1249), .ZN(n1065) );
XOR2_X1 U936 ( .A(n1205), .B(n1257), .Z(G21) );
NAND2_X1 U937 ( .A1(KEYINPUT38), .A2(G119), .ZN(n1257) );
NAND4_X1 U938 ( .A1(n1258), .A2(n1056), .A3(n1249), .A4(n1095), .ZN(n1205) );
XNOR2_X1 U939 ( .A(G116), .B(n1206), .ZN(G18) );
NAND4_X1 U940 ( .A1(n1056), .A2(n1241), .A3(n1219), .A4(n1075), .ZN(n1206) );
NOR2_X1 U941 ( .A1(n1239), .A2(n1084), .ZN(n1075) );
XNOR2_X1 U942 ( .A(G113), .B(n1259), .ZN(G15) );
NAND4_X1 U943 ( .A1(n1252), .A2(n1241), .A3(n1260), .A4(n1261), .ZN(n1259) );
XNOR2_X1 U944 ( .A(KEYINPUT46), .B(n1067), .ZN(n1260) );
INV_X1 U945 ( .A(n1064), .ZN(n1241) );
NAND2_X1 U946 ( .A1(n1262), .A2(n1095), .ZN(n1064) );
INV_X1 U947 ( .A(n1073), .ZN(n1252) );
NAND2_X1 U948 ( .A1(n1218), .A2(n1056), .ZN(n1073) );
NOR2_X1 U949 ( .A1(n1263), .A2(n1079), .ZN(n1056) );
INV_X1 U950 ( .A(n1203), .ZN(n1218) );
NAND2_X1 U951 ( .A1(n1239), .A2(n1084), .ZN(n1203) );
INV_X1 U952 ( .A(n1242), .ZN(n1084) );
XNOR2_X1 U953 ( .A(G110), .B(n1264), .ZN(G12) );
NAND3_X1 U954 ( .A1(n1258), .A2(n1216), .A3(n1217), .ZN(n1264) );
NOR2_X1 U955 ( .A1(n1095), .A2(n1262), .ZN(n1217) );
INV_X1 U956 ( .A(n1249), .ZN(n1262) );
XNOR2_X1 U957 ( .A(n1099), .B(n1098), .ZN(n1249) );
NAND2_X1 U958 ( .A1(G217), .A2(n1265), .ZN(n1098) );
NOR2_X1 U959 ( .A1(n1141), .A2(G902), .ZN(n1099) );
XNOR2_X1 U960 ( .A(n1266), .B(n1267), .ZN(n1141) );
AND3_X1 U961 ( .A1(G221), .A2(n1050), .A3(G234), .ZN(n1267) );
XOR2_X1 U962 ( .A(n1268), .B(G137), .Z(n1266) );
NAND2_X1 U963 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U964 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U965 ( .A(n1273), .B(KEYINPUT26), .Z(n1269) );
OR2_X1 U966 ( .A1(n1272), .A2(n1271), .ZN(n1273) );
XNOR2_X1 U967 ( .A(n1274), .B(n1275), .ZN(n1271) );
NOR2_X1 U968 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
AND3_X1 U969 ( .A1(KEYINPUT51), .A2(n1278), .A3(G140), .ZN(n1277) );
NOR2_X1 U970 ( .A1(KEYINPUT51), .A2(n1279), .ZN(n1276) );
NAND2_X1 U971 ( .A1(KEYINPUT61), .A2(n1280), .ZN(n1274) );
XOR2_X1 U972 ( .A(G110), .B(n1281), .Z(n1272) );
XNOR2_X1 U973 ( .A(n1251), .B(G119), .ZN(n1281) );
INV_X1 U974 ( .A(G128), .ZN(n1251) );
XOR2_X1 U975 ( .A(n1282), .B(n1165), .Z(n1095) );
INV_X1 U976 ( .A(G472), .ZN(n1165) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U978 ( .A(n1285), .B(n1286), .Z(n1283) );
XOR2_X1 U979 ( .A(n1172), .B(n1169), .Z(n1286) );
XOR2_X1 U980 ( .A(n1287), .B(n1288), .Z(n1169) );
XNOR2_X1 U981 ( .A(G113), .B(KEYINPUT48), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1289), .B(n1290), .Z(n1285) );
XOR2_X1 U983 ( .A(G101), .B(n1175), .Z(n1290) );
AND3_X1 U984 ( .A1(n1291), .A2(n1050), .A3(n1292), .ZN(n1175) );
XOR2_X1 U985 ( .A(KEYINPUT10), .B(G210), .Z(n1292) );
NAND2_X1 U986 ( .A1(KEYINPUT59), .A2(n1293), .ZN(n1289) );
NOR2_X1 U987 ( .A1(n1080), .A2(n1079), .ZN(n1216) );
AND2_X1 U988 ( .A1(G221), .A2(n1265), .ZN(n1079) );
NAND2_X1 U989 ( .A1(G234), .A2(n1284), .ZN(n1265) );
INV_X1 U990 ( .A(n1263), .ZN(n1080) );
XNOR2_X1 U991 ( .A(n1092), .B(G469), .ZN(n1263) );
NAND2_X1 U992 ( .A1(n1294), .A2(n1284), .ZN(n1092) );
XOR2_X1 U993 ( .A(n1179), .B(n1295), .Z(n1294) );
XOR2_X1 U994 ( .A(n1296), .B(n1182), .Z(n1295) );
XOR2_X1 U995 ( .A(n1297), .B(n1109), .Z(n1182) );
AND2_X1 U996 ( .A1(n1298), .A2(n1299), .ZN(n1109) );
NAND2_X1 U997 ( .A1(G128), .A2(n1300), .ZN(n1299) );
XOR2_X1 U998 ( .A(n1301), .B(KEYINPUT20), .Z(n1298) );
OR2_X1 U999 ( .A1(n1300), .A2(G128), .ZN(n1301) );
NAND3_X1 U1000 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1300) );
OR2_X1 U1001 ( .A1(n1305), .A2(G143), .ZN(n1304) );
NAND2_X1 U1002 ( .A1(n1306), .A2(n1307), .ZN(n1303) );
INV_X1 U1003 ( .A(KEYINPUT47), .ZN(n1307) );
NAND2_X1 U1004 ( .A1(n1308), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U1005 ( .A(KEYINPUT24), .B(G143), .ZN(n1308) );
NAND2_X1 U1006 ( .A1(KEYINPUT47), .A2(n1309), .ZN(n1302) );
NAND2_X1 U1007 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
OR2_X1 U1008 ( .A1(G143), .A2(KEYINPUT24), .ZN(n1311) );
NAND3_X1 U1009 ( .A1(G143), .A2(n1305), .A3(KEYINPUT24), .ZN(n1310) );
XOR2_X1 U1010 ( .A(n1280), .B(KEYINPUT23), .Z(n1305) );
NOR2_X1 U1011 ( .A1(KEYINPUT50), .A2(n1172), .ZN(n1296) );
XOR2_X1 U1012 ( .A(n1107), .B(KEYINPUT56), .Z(n1172) );
XNOR2_X1 U1013 ( .A(G131), .B(n1312), .ZN(n1107) );
XOR2_X1 U1014 ( .A(G137), .B(G134), .Z(n1312) );
XOR2_X1 U1015 ( .A(n1313), .B(n1314), .Z(n1179) );
XOR2_X1 U1016 ( .A(G140), .B(G110), .Z(n1314) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1050), .ZN(n1313) );
INV_X1 U1018 ( .A(n1215), .ZN(n1258) );
NAND2_X1 U1019 ( .A1(n1058), .A2(n1219), .ZN(n1215) );
INV_X1 U1020 ( .A(n1213), .ZN(n1219) );
NAND2_X1 U1021 ( .A1(n1226), .A2(n1261), .ZN(n1213) );
NAND2_X1 U1022 ( .A1(n1315), .A2(n1081), .ZN(n1261) );
NAND3_X1 U1023 ( .A1(n1254), .A2(n1050), .A3(G952), .ZN(n1081) );
NAND4_X1 U1024 ( .A1(n1316), .A2(G902), .A3(n1254), .A4(n1130), .ZN(n1315) );
INV_X1 U1025 ( .A(G898), .ZN(n1130) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1254) );
XNOR2_X1 U1027 ( .A(G953), .B(KEYINPUT52), .ZN(n1316) );
INV_X1 U1028 ( .A(n1067), .ZN(n1226) );
NAND2_X1 U1029 ( .A1(n1247), .A2(n1096), .ZN(n1067) );
XNOR2_X1 U1030 ( .A(n1189), .B(n1317), .ZN(n1096) );
NOR2_X1 U1031 ( .A1(G902), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1032 ( .A(n1222), .B(n1319), .Z(n1318) );
NOR2_X1 U1033 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NOR2_X1 U1034 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1035 ( .A(KEYINPUT0), .B(n1224), .Z(n1323) );
INV_X1 U1036 ( .A(n1324), .ZN(n1322) );
NOR2_X1 U1037 ( .A1(n1224), .A2(n1324), .ZN(n1320) );
NAND2_X1 U1038 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1039 ( .A1(G125), .A2(n1293), .ZN(n1326) );
XOR2_X1 U1040 ( .A(KEYINPUT12), .B(n1327), .Z(n1325) );
NOR2_X1 U1041 ( .A1(G125), .A2(n1293), .ZN(n1327) );
INV_X1 U1042 ( .A(n1171), .ZN(n1293) );
XNOR2_X1 U1043 ( .A(n1328), .B(n1280), .ZN(n1171) );
NOR2_X1 U1044 ( .A1(n1124), .A2(G953), .ZN(n1224) );
INV_X1 U1045 ( .A(G224), .ZN(n1124) );
NAND3_X1 U1046 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1222) );
NAND2_X1 U1047 ( .A1(n1132), .A2(n1332), .ZN(n1331) );
INV_X1 U1048 ( .A(KEYINPUT7), .ZN(n1332) );
NAND3_X1 U1049 ( .A1(KEYINPUT7), .A2(n1333), .A3(n1334), .ZN(n1330) );
OR2_X1 U1050 ( .A1(n1334), .A2(n1333), .ZN(n1329) );
NOR2_X1 U1051 ( .A1(n1335), .A2(n1132), .ZN(n1333) );
XOR2_X1 U1052 ( .A(G110), .B(n1336), .Z(n1132) );
XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n1337), .ZN(n1336) );
INV_X1 U1054 ( .A(KEYINPUT53), .ZN(n1335) );
NAND3_X1 U1055 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1334) );
OR2_X1 U1056 ( .A1(n1341), .A2(n1136), .ZN(n1340) );
NAND3_X1 U1057 ( .A1(n1136), .A2(n1341), .A3(n1135), .ZN(n1339) );
NAND2_X1 U1058 ( .A1(n1342), .A2(n1343), .ZN(n1338) );
NAND2_X1 U1059 ( .A1(n1344), .A2(n1341), .ZN(n1343) );
INV_X1 U1060 ( .A(KEYINPUT34), .ZN(n1341) );
XOR2_X1 U1061 ( .A(n1136), .B(KEYINPUT31), .Z(n1344) );
XOR2_X1 U1062 ( .A(n1345), .B(KEYINPUT45), .Z(n1136) );
NAND2_X1 U1063 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND3_X1 U1064 ( .A1(G101), .A2(n1348), .A3(n1349), .ZN(n1347) );
INV_X1 U1065 ( .A(KEYINPUT22), .ZN(n1349) );
NAND2_X1 U1066 ( .A1(n1297), .A2(KEYINPUT22), .ZN(n1346) );
XOR2_X1 U1067 ( .A(G101), .B(n1348), .Z(n1297) );
XNOR2_X1 U1068 ( .A(G107), .B(n1350), .ZN(n1348) );
INV_X1 U1069 ( .A(n1135), .ZN(n1342) );
XOR2_X1 U1070 ( .A(G113), .B(n1351), .Z(n1135) );
NOR2_X1 U1071 ( .A1(KEYINPUT1), .A2(n1288), .ZN(n1351) );
XNOR2_X1 U1072 ( .A(G116), .B(G119), .ZN(n1288) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1352), .ZN(n1189) );
XOR2_X1 U1074 ( .A(n1070), .B(KEYINPUT57), .Z(n1247) );
AND2_X1 U1075 ( .A1(G214), .A2(n1352), .ZN(n1070) );
NAND2_X1 U1076 ( .A1(n1291), .A2(n1284), .ZN(n1352) );
NOR2_X1 U1077 ( .A1(n1242), .A2(n1239), .ZN(n1058) );
XNOR2_X1 U1078 ( .A(n1353), .B(n1089), .ZN(n1239) );
NAND2_X1 U1079 ( .A1(n1152), .A2(n1284), .ZN(n1089) );
XOR2_X1 U1080 ( .A(n1354), .B(n1355), .Z(n1152) );
NOR2_X1 U1081 ( .A1(KEYINPUT19), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1082 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1083 ( .A(n1359), .B(n1279), .Z(n1358) );
XNOR2_X1 U1084 ( .A(G140), .B(n1278), .ZN(n1279) );
INV_X1 U1085 ( .A(G125), .ZN(n1278) );
AND3_X1 U1086 ( .A1(G214), .A2(n1050), .A3(n1291), .ZN(n1359) );
INV_X1 U1087 ( .A(G237), .ZN(n1291) );
XOR2_X1 U1088 ( .A(n1360), .B(n1361), .Z(n1357) );
XNOR2_X1 U1089 ( .A(n1237), .B(G131), .ZN(n1361) );
NAND2_X1 U1090 ( .A1(KEYINPUT8), .A2(n1280), .ZN(n1360) );
XNOR2_X1 U1091 ( .A(G146), .B(KEYINPUT29), .ZN(n1280) );
NAND3_X1 U1092 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1354) );
NAND2_X1 U1093 ( .A1(n1365), .A2(G104), .ZN(n1364) );
NAND2_X1 U1094 ( .A1(n1366), .A2(n1367), .ZN(n1363) );
INV_X1 U1095 ( .A(KEYINPUT25), .ZN(n1367) );
NAND2_X1 U1096 ( .A1(n1368), .A2(n1350), .ZN(n1366) );
INV_X1 U1097 ( .A(G104), .ZN(n1350) );
XNOR2_X1 U1098 ( .A(KEYINPUT36), .B(n1365), .ZN(n1368) );
NAND2_X1 U1099 ( .A1(KEYINPUT25), .A2(n1369), .ZN(n1362) );
NAND2_X1 U1100 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1101 ( .A1(KEYINPUT36), .A2(n1365), .ZN(n1371) );
OR3_X1 U1102 ( .A1(G104), .A2(KEYINPUT36), .A3(n1365), .ZN(n1370) );
XNOR2_X1 U1103 ( .A(n1372), .B(n1373), .ZN(n1365) );
INV_X1 U1104 ( .A(G113), .ZN(n1373) );
NAND2_X1 U1105 ( .A1(KEYINPUT54), .A2(n1337), .ZN(n1372) );
NAND2_X1 U1106 ( .A1(KEYINPUT44), .A2(n1091), .ZN(n1353) );
INV_X1 U1107 ( .A(G475), .ZN(n1091) );
XNOR2_X1 U1108 ( .A(n1374), .B(G478), .ZN(n1242) );
NAND2_X1 U1109 ( .A1(n1284), .A2(n1148), .ZN(n1374) );
NAND2_X1 U1110 ( .A1(n1375), .A2(n1376), .ZN(n1148) );
NAND4_X1 U1111 ( .A1(G217), .A2(G234), .A3(n1377), .A4(n1378), .ZN(n1376) );
NOR2_X1 U1112 ( .A1(G953), .A2(n1379), .ZN(n1377) );
NAND2_X1 U1113 ( .A1(n1380), .A2(n1381), .ZN(n1375) );
NAND3_X1 U1114 ( .A1(G234), .A2(n1050), .A3(G217), .ZN(n1381) );
INV_X1 U1115 ( .A(G953), .ZN(n1050) );
NAND2_X1 U1116 ( .A1(n1378), .A2(n1382), .ZN(n1380) );
INV_X1 U1117 ( .A(n1379), .ZN(n1382) );
NOR2_X1 U1118 ( .A1(n1383), .A2(n1384), .ZN(n1379) );
XNOR2_X1 U1119 ( .A(n1385), .B(KEYINPUT30), .ZN(n1378) );
NAND2_X1 U1120 ( .A1(n1384), .A2(n1383), .ZN(n1385) );
XNOR2_X1 U1121 ( .A(n1386), .B(n1387), .ZN(n1383) );
XNOR2_X1 U1122 ( .A(KEYINPUT28), .B(n1337), .ZN(n1387) );
INV_X1 U1123 ( .A(G122), .ZN(n1337) );
XNOR2_X1 U1124 ( .A(G107), .B(G116), .ZN(n1386) );
XNOR2_X1 U1125 ( .A(G134), .B(n1328), .ZN(n1384) );
XNOR2_X1 U1126 ( .A(G128), .B(n1237), .ZN(n1328) );
INV_X1 U1127 ( .A(G143), .ZN(n1237) );
INV_X1 U1128 ( .A(G902), .ZN(n1284) );
endmodule


