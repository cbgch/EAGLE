//Key = 0101001000110010010101100011101110000100101010110101001001010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343;

XOR2_X1 U739 ( .A(n1025), .B(n1026), .Z(G9) );
NOR2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U742 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1029) );
NAND2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND4_X1 U745 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
NAND3_X1 U746 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
NAND2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NAND2_X1 U749 ( .A1(n1050), .A2(n1051), .ZN(n1043) );
NAND3_X1 U750 ( .A1(n1050), .A2(n1052), .A3(n1048), .ZN(n1037) );
NAND2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1039), .ZN(n1054) );
NAND2_X1 U753 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XOR2_X1 U754 ( .A(n1059), .B(KEYINPUT18), .Z(n1058) );
NAND3_X1 U755 ( .A1(n1060), .A2(n1061), .A3(n1042), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
INV_X1 U757 ( .A(n1064), .ZN(n1062) );
NAND2_X1 U758 ( .A1(n1040), .A2(n1065), .ZN(n1053) );
INV_X1 U759 ( .A(n1066), .ZN(n1035) );
AND3_X1 U760 ( .A1(n1034), .A2(n1067), .A3(n1033), .ZN(n1027) );
NAND4_X1 U761 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1033) );
NOR3_X1 U762 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
NAND3_X1 U765 ( .A1(n1064), .A2(n1079), .A3(n1042), .ZN(n1072) );
NOR3_X1 U766 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1083), .B(n1084), .Z(n1081) );
NOR2_X1 U768 ( .A1(KEYINPUT25), .A2(n1085), .ZN(n1084) );
XOR2_X1 U769 ( .A(n1086), .B(n1087), .Z(n1080) );
NOR2_X1 U770 ( .A1(KEYINPUT33), .A2(n1088), .ZN(n1087) );
XOR2_X1 U771 ( .A(n1089), .B(G472), .Z(n1069) );
NAND2_X1 U772 ( .A1(KEYINPUT21), .A2(n1090), .ZN(n1089) );
XOR2_X1 U773 ( .A(n1091), .B(KEYINPUT7), .Z(n1068) );
NAND2_X1 U774 ( .A1(n1075), .A2(n1076), .ZN(n1091) );
INV_X1 U775 ( .A(G952), .ZN(n1067) );
XOR2_X1 U776 ( .A(n1092), .B(n1093), .Z(G72) );
XOR2_X1 U777 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U778 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U779 ( .A(KEYINPUT58), .B(G953), .Z(n1097) );
INV_X1 U780 ( .A(n1031), .ZN(n1096) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
INV_X1 U782 ( .A(n1100), .ZN(n1099) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1098) );
XNOR2_X1 U784 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U785 ( .A1(KEYINPUT39), .A2(n1105), .ZN(n1104) );
XOR2_X1 U786 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U787 ( .A1(KEYINPUT5), .A2(n1108), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1109), .B(G140), .Z(n1101) );
NAND2_X1 U789 ( .A1(G953), .A2(n1110), .ZN(n1092) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1110) );
NAND2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(G69) );
NAND2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U793 ( .A(n1115), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
NAND2_X1 U795 ( .A1(n1117), .A2(n1114), .ZN(n1116) );
NAND2_X1 U796 ( .A1(G953), .A2(n1118), .ZN(n1114) );
INV_X1 U797 ( .A(n1119), .ZN(n1117) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(n1115) );
NOR4_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1119), .A4(n1124), .ZN(n1121) );
INV_X1 U800 ( .A(n1125), .ZN(n1124) );
NOR2_X1 U801 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
XOR2_X1 U802 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U803 ( .A(n1130), .B(KEYINPUT59), .Z(n1128) );
NOR3_X1 U804 ( .A1(n1131), .A2(n1129), .A3(n1130), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1030), .ZN(n1120) );
NOR3_X1 U806 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(G66) );
AND2_X1 U807 ( .A1(KEYINPUT30), .A2(n1136), .ZN(n1135) );
NOR3_X1 U808 ( .A1(KEYINPUT30), .A2(G953), .A3(G952), .ZN(n1134) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1133) );
NOR2_X1 U810 ( .A1(n1078), .A2(n1139), .ZN(n1138) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1140), .ZN(G63) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U813 ( .A1(n1088), .A2(n1139), .ZN(n1141) );
INV_X1 U814 ( .A(G478), .ZN(n1088) );
NOR2_X1 U815 ( .A1(n1136), .A2(n1143), .ZN(G60) );
XOR2_X1 U816 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U817 ( .A1(n1146), .A2(KEYINPUT56), .ZN(n1145) );
AND2_X1 U818 ( .A1(G475), .A2(n1147), .ZN(n1146) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(G6) );
NAND2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U821 ( .A(KEYINPUT14), .B(n1152), .Z(n1148) );
NOR2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1136), .A2(n1153), .ZN(G57) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U826 ( .A1(KEYINPUT47), .A2(n1158), .ZN(n1156) );
XOR2_X1 U827 ( .A(n1159), .B(n1160), .Z(n1154) );
NOR2_X1 U828 ( .A1(KEYINPUT53), .A2(n1161), .ZN(n1160) );
XOR2_X1 U829 ( .A(n1162), .B(KEYINPUT4), .Z(n1159) );
NAND2_X1 U830 ( .A1(n1147), .A2(G472), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1136), .A2(n1163), .ZN(G54) );
NOR2_X1 U832 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
XOR2_X1 U835 ( .A(KEYINPUT17), .B(n1167), .Z(n1169) );
XNOR2_X1 U836 ( .A(n1170), .B(n1171), .ZN(n1167) );
XNOR2_X1 U837 ( .A(n1172), .B(n1173), .ZN(n1170) );
NOR2_X1 U838 ( .A1(KEYINPUT24), .A2(n1174), .ZN(n1173) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U840 ( .A(G140), .B(n1177), .Z(n1176) );
NAND2_X1 U841 ( .A1(KEYINPUT57), .A2(n1178), .ZN(n1175) );
XNOR2_X1 U842 ( .A(n1166), .B(KEYINPUT35), .ZN(n1168) );
NOR2_X1 U843 ( .A1(n1139), .A2(n1076), .ZN(n1166) );
INV_X1 U844 ( .A(G469), .ZN(n1076) );
NOR2_X1 U845 ( .A1(n1136), .A2(n1179), .ZN(G51) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U847 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND3_X1 U848 ( .A1(n1147), .A2(G210), .A3(KEYINPUT46), .ZN(n1182) );
INV_X1 U849 ( .A(n1139), .ZN(n1147) );
NAND2_X1 U850 ( .A1(G902), .A2(n1184), .ZN(n1139) );
OR2_X1 U851 ( .A1(n1031), .A2(n1030), .ZN(n1184) );
NAND4_X1 U852 ( .A1(n1185), .A2(n1026), .A3(n1186), .A4(n1187), .ZN(n1030) );
NOR3_X1 U853 ( .A1(n1150), .A2(n1188), .A3(n1189), .ZN(n1187) );
AND3_X1 U854 ( .A1(n1190), .A2(n1050), .A3(n1191), .ZN(n1150) );
NAND3_X1 U855 ( .A1(n1065), .A2(n1192), .A3(n1193), .ZN(n1186) );
NAND2_X1 U856 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NAND2_X1 U857 ( .A1(n1049), .A2(n1051), .ZN(n1195) );
NAND2_X1 U858 ( .A1(n1196), .A2(n1197), .ZN(n1051) );
NAND2_X1 U859 ( .A1(n1046), .A2(n1198), .ZN(n1194) );
NAND3_X1 U860 ( .A1(n1050), .A2(n1199), .A3(n1190), .ZN(n1026) );
NAND4_X1 U861 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1031) );
NOR4_X1 U862 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
INV_X1 U863 ( .A(n1208), .ZN(n1204) );
NOR2_X1 U864 ( .A1(n1209), .A2(n1210), .ZN(n1202) );
NOR3_X1 U865 ( .A1(n1211), .A2(n1061), .A3(n1197), .ZN(n1210) );
NOR4_X1 U866 ( .A1(n1212), .A2(n1198), .A3(n1213), .A4(n1214), .ZN(n1209) );
XOR2_X1 U867 ( .A(KEYINPUT62), .B(n1191), .Z(n1214) );
NOR2_X1 U868 ( .A1(n1132), .A2(G952), .ZN(n1136) );
XNOR2_X1 U869 ( .A(G146), .B(n1201), .ZN(G48) );
OR3_X1 U870 ( .A1(n1196), .A2(n1061), .A3(n1211), .ZN(n1201) );
XOR2_X1 U871 ( .A(n1215), .B(n1200), .Z(G45) );
NAND4_X1 U872 ( .A1(n1216), .A2(n1049), .A3(n1217), .A4(n1218), .ZN(n1200) );
XOR2_X1 U873 ( .A(G140), .B(n1219), .Z(G42) );
NOR4_X1 U874 ( .A1(n1212), .A2(n1198), .A3(n1196), .A4(n1213), .ZN(n1219) );
XOR2_X1 U875 ( .A(G137), .B(n1207), .Z(G39) );
NOR3_X1 U876 ( .A1(n1047), .A2(n1213), .A3(n1220), .ZN(n1207) );
XOR2_X1 U877 ( .A(G134), .B(n1206), .Z(G36) );
NOR3_X1 U878 ( .A1(n1221), .A2(n1197), .A3(n1213), .ZN(n1206) );
XOR2_X1 U879 ( .A(n1222), .B(n1205), .Z(G33) );
NOR3_X1 U880 ( .A1(n1221), .A2(n1196), .A3(n1213), .ZN(n1205) );
NAND4_X1 U881 ( .A1(n1039), .A2(n1217), .A3(n1218), .A4(n1042), .ZN(n1213) );
NAND2_X1 U882 ( .A1(KEYINPUT40), .A2(n1223), .ZN(n1222) );
XOR2_X1 U883 ( .A(G128), .B(n1224), .Z(G30) );
NOR3_X1 U884 ( .A1(n1225), .A2(n1197), .A3(n1211), .ZN(n1224) );
NAND4_X1 U885 ( .A1(n1198), .A2(n1065), .A3(n1218), .A4(n1226), .ZN(n1211) );
INV_X1 U886 ( .A(n1199), .ZN(n1197) );
XOR2_X1 U887 ( .A(KEYINPUT28), .B(n1217), .Z(n1225) );
INV_X1 U888 ( .A(n1061), .ZN(n1217) );
XOR2_X1 U889 ( .A(n1189), .B(n1227), .Z(G3) );
NOR2_X1 U890 ( .A1(KEYINPUT34), .A2(n1158), .ZN(n1227) );
INV_X1 U891 ( .A(G101), .ZN(n1158) );
AND3_X1 U892 ( .A1(n1049), .A2(n1190), .A3(n1048), .ZN(n1189) );
XOR2_X1 U893 ( .A(n1109), .B(n1208), .Z(G27) );
NAND4_X1 U894 ( .A1(n1191), .A2(n1065), .A3(n1040), .A4(n1228), .ZN(n1208) );
AND3_X1 U895 ( .A1(n1047), .A2(n1226), .A3(n1218), .ZN(n1228) );
NAND2_X1 U896 ( .A1(n1066), .A2(n1229), .ZN(n1218) );
NAND3_X1 U897 ( .A1(G902), .A2(n1230), .A3(n1100), .ZN(n1229) );
NOR2_X1 U898 ( .A1(n1132), .A2(G900), .ZN(n1100) );
INV_X1 U899 ( .A(n1059), .ZN(n1040) );
XOR2_X1 U900 ( .A(n1231), .B(n1185), .Z(G24) );
NAND3_X1 U901 ( .A1(n1216), .A2(n1050), .A3(n1193), .ZN(n1185) );
NOR2_X1 U902 ( .A1(n1226), .A2(n1198), .ZN(n1050) );
NOR3_X1 U903 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1216) );
XNOR2_X1 U904 ( .A(G119), .B(n1235), .ZN(G21) );
NAND4_X1 U905 ( .A1(n1193), .A2(n1046), .A3(n1198), .A4(n1236), .ZN(n1235) );
XOR2_X1 U906 ( .A(KEYINPUT8), .B(n1065), .Z(n1236) );
XNOR2_X1 U907 ( .A(G116), .B(n1237), .ZN(G18) );
NAND4_X1 U908 ( .A1(n1238), .A2(n1049), .A3(n1239), .A4(n1199), .ZN(n1237) );
NOR2_X1 U909 ( .A1(n1233), .A2(n1240), .ZN(n1199) );
NOR2_X1 U910 ( .A1(n1241), .A2(n1232), .ZN(n1239) );
INV_X1 U911 ( .A(n1221), .ZN(n1049) );
XOR2_X1 U912 ( .A(n1059), .B(KEYINPUT49), .Z(n1238) );
XOR2_X1 U913 ( .A(n1242), .B(n1243), .Z(G15) );
NAND4_X1 U914 ( .A1(n1244), .A2(n1193), .A3(n1191), .A4(n1065), .ZN(n1243) );
INV_X1 U915 ( .A(n1196), .ZN(n1191) );
NAND2_X1 U916 ( .A1(n1245), .A2(n1240), .ZN(n1196) );
XOR2_X1 U917 ( .A(n1233), .B(KEYINPUT13), .Z(n1245) );
NOR2_X1 U918 ( .A1(n1059), .A2(n1241), .ZN(n1193) );
NAND2_X1 U919 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
XNOR2_X1 U920 ( .A(n1246), .B(KEYINPUT50), .ZN(n1063) );
XOR2_X1 U921 ( .A(n1221), .B(KEYINPUT37), .Z(n1244) );
NAND2_X1 U922 ( .A1(n1198), .A2(n1212), .ZN(n1221) );
INV_X1 U923 ( .A(n1226), .ZN(n1212) );
XOR2_X1 U924 ( .A(n1188), .B(n1247), .Z(G12) );
NOR2_X1 U925 ( .A1(KEYINPUT36), .A2(n1248), .ZN(n1247) );
XOR2_X1 U926 ( .A(KEYINPUT32), .B(G110), .Z(n1248) );
AND3_X1 U927 ( .A1(n1190), .A2(n1047), .A3(n1046), .ZN(n1188) );
INV_X1 U928 ( .A(n1220), .ZN(n1046) );
NAND2_X1 U929 ( .A1(n1048), .A2(n1226), .ZN(n1220) );
NAND3_X1 U930 ( .A1(n1249), .A2(n1250), .A3(n1079), .ZN(n1226) );
NAND2_X1 U931 ( .A1(n1077), .A2(n1078), .ZN(n1079) );
OR3_X1 U932 ( .A1(n1078), .A2(n1077), .A3(KEYINPUT38), .ZN(n1250) );
NAND2_X1 U933 ( .A1(G217), .A2(n1251), .ZN(n1078) );
NAND2_X1 U934 ( .A1(KEYINPUT38), .A2(n1077), .ZN(n1249) );
NOR2_X1 U935 ( .A1(n1137), .A2(G902), .ZN(n1077) );
XOR2_X1 U936 ( .A(n1252), .B(n1253), .Z(n1137) );
XOR2_X1 U937 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND3_X1 U938 ( .A1(G234), .A2(n1132), .A3(G221), .ZN(n1255) );
NAND2_X1 U939 ( .A1(n1256), .A2(KEYINPUT44), .ZN(n1254) );
XOR2_X1 U940 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U941 ( .A(G128), .B(G119), .Z(n1258) );
XOR2_X1 U942 ( .A(n1178), .B(n1259), .Z(n1257) );
NOR2_X1 U943 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U944 ( .A(KEYINPUT27), .B(KEYINPUT22), .Z(n1261) );
XOR2_X1 U945 ( .A(n1262), .B(n1263), .Z(n1260) );
NOR2_X1 U946 ( .A1(KEYINPUT2), .A2(n1264), .ZN(n1263) );
XOR2_X1 U947 ( .A(G146), .B(n1109), .Z(n1262) );
INV_X1 U948 ( .A(G125), .ZN(n1109) );
XNOR2_X1 U949 ( .A(G137), .B(KEYINPUT3), .ZN(n1252) );
AND2_X1 U950 ( .A1(n1233), .A2(n1234), .ZN(n1048) );
INV_X1 U951 ( .A(n1240), .ZN(n1234) );
XNOR2_X1 U952 ( .A(n1082), .B(KEYINPUT51), .ZN(n1240) );
XNOR2_X1 U953 ( .A(n1265), .B(G475), .ZN(n1082) );
NAND2_X1 U954 ( .A1(n1144), .A2(n1266), .ZN(n1265) );
XOR2_X1 U955 ( .A(n1267), .B(n1268), .Z(n1144) );
XOR2_X1 U956 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U957 ( .A(G113), .B(G104), .Z(n1270) );
XOR2_X1 U958 ( .A(G131), .B(G125), .Z(n1269) );
XOR2_X1 U959 ( .A(n1271), .B(n1272), .Z(n1267) );
XOR2_X1 U960 ( .A(n1273), .B(n1264), .Z(n1272) );
XOR2_X1 U961 ( .A(G140), .B(KEYINPUT26), .Z(n1264) );
XOR2_X1 U962 ( .A(n1274), .B(n1275), .Z(n1271) );
NOR2_X1 U963 ( .A1(KEYINPUT20), .A2(n1231), .ZN(n1275) );
INV_X1 U964 ( .A(G122), .ZN(n1231) );
NAND2_X1 U965 ( .A1(n1276), .A2(G214), .ZN(n1274) );
XNOR2_X1 U966 ( .A(n1086), .B(G478), .ZN(n1233) );
NOR2_X1 U967 ( .A1(n1142), .A2(G902), .ZN(n1086) );
XNOR2_X1 U968 ( .A(n1277), .B(n1278), .ZN(n1142) );
XOR2_X1 U969 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U970 ( .A(G134), .B(G128), .Z(n1280) );
XOR2_X1 U971 ( .A(KEYINPUT52), .B(G143), .Z(n1279) );
XOR2_X1 U972 ( .A(n1281), .B(n1282), .Z(n1277) );
XOR2_X1 U973 ( .A(G122), .B(G107), .Z(n1282) );
XOR2_X1 U974 ( .A(n1283), .B(n1284), .Z(n1281) );
NOR2_X1 U975 ( .A1(G116), .A2(KEYINPUT48), .ZN(n1284) );
NAND3_X1 U976 ( .A1(G234), .A2(n1132), .A3(G217), .ZN(n1283) );
INV_X1 U977 ( .A(n1198), .ZN(n1047) );
XOR2_X1 U978 ( .A(n1285), .B(n1286), .Z(n1198) );
NOR2_X1 U979 ( .A1(KEYINPUT45), .A2(G472), .ZN(n1286) );
XNOR2_X1 U980 ( .A(n1090), .B(KEYINPUT23), .ZN(n1285) );
AND2_X1 U981 ( .A1(n1287), .A2(n1266), .ZN(n1090) );
XOR2_X1 U982 ( .A(n1288), .B(n1289), .Z(n1287) );
INV_X1 U983 ( .A(n1161), .ZN(n1289) );
XOR2_X1 U984 ( .A(n1157), .B(G101), .Z(n1288) );
XNOR2_X1 U985 ( .A(n1172), .B(n1290), .ZN(n1157) );
XOR2_X1 U986 ( .A(n1291), .B(n1292), .Z(n1290) );
INV_X1 U987 ( .A(n1130), .ZN(n1292) );
AND2_X1 U988 ( .A1(G210), .A2(n1276), .ZN(n1291) );
NOR2_X1 U989 ( .A1(G953), .A2(G237), .ZN(n1276) );
NOR3_X1 U990 ( .A1(n1061), .A2(n1241), .A3(n1232), .ZN(n1190) );
INV_X1 U991 ( .A(n1065), .ZN(n1232) );
NOR2_X1 U992 ( .A1(n1039), .A2(n1057), .ZN(n1065) );
INV_X1 U993 ( .A(n1042), .ZN(n1057) );
NAND2_X1 U994 ( .A1(G214), .A2(n1293), .ZN(n1042) );
XNOR2_X1 U995 ( .A(n1294), .B(n1083), .ZN(n1039) );
NAND2_X1 U996 ( .A1(G210), .A2(n1293), .ZN(n1083) );
NAND2_X1 U997 ( .A1(n1295), .A2(n1266), .ZN(n1293) );
XOR2_X1 U998 ( .A(KEYINPUT6), .B(G237), .Z(n1295) );
NAND2_X1 U999 ( .A1(KEYINPUT1), .A2(n1085), .ZN(n1294) );
AND2_X1 U1000 ( .A1(n1296), .A2(n1266), .ZN(n1085) );
XOR2_X1 U1001 ( .A(n1183), .B(n1297), .Z(n1296) );
NOR2_X1 U1002 ( .A1(KEYINPUT61), .A2(n1298), .ZN(n1297) );
XOR2_X1 U1003 ( .A(n1180), .B(KEYINPUT29), .Z(n1298) );
XOR2_X1 U1004 ( .A(n1299), .B(n1300), .Z(n1180) );
XOR2_X1 U1005 ( .A(KEYINPUT0), .B(G125), .Z(n1300) );
XOR2_X1 U1006 ( .A(n1161), .B(n1301), .Z(n1299) );
NOR2_X1 U1007 ( .A1(G953), .A2(n1118), .ZN(n1301) );
INV_X1 U1008 ( .A(G224), .ZN(n1118) );
XOR2_X1 U1009 ( .A(n1302), .B(n1303), .Z(n1161) );
NOR2_X1 U1010 ( .A1(KEYINPUT15), .A2(n1304), .ZN(n1303) );
NAND3_X1 U1011 ( .A1(n1305), .A2(n1306), .A3(n1125), .ZN(n1183) );
NAND3_X1 U1012 ( .A1(n1129), .A2(n1126), .A3(n1130), .ZN(n1125) );
NAND3_X1 U1013 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
NAND2_X1 U1014 ( .A1(n1130), .A2(n1126), .ZN(n1308) );
OR2_X1 U1015 ( .A1(n1309), .A2(n1307), .ZN(n1305) );
INV_X1 U1016 ( .A(n1129), .ZN(n1307) );
XNOR2_X1 U1017 ( .A(n1178), .B(G122), .ZN(n1129) );
XNOR2_X1 U1018 ( .A(n1310), .B(KEYINPUT42), .ZN(n1309) );
NAND2_X1 U1019 ( .A1(n1311), .A2(n1131), .ZN(n1310) );
INV_X1 U1020 ( .A(n1126), .ZN(n1131) );
NAND2_X1 U1021 ( .A1(n1312), .A2(n1313), .ZN(n1126) );
INV_X1 U1022 ( .A(n1314), .ZN(n1312) );
XOR2_X1 U1023 ( .A(n1130), .B(KEYINPUT10), .Z(n1311) );
XOR2_X1 U1024 ( .A(n1242), .B(n1315), .Z(n1130) );
XOR2_X1 U1025 ( .A(G119), .B(G116), .Z(n1315) );
INV_X1 U1026 ( .A(G113), .ZN(n1242) );
AND2_X1 U1027 ( .A1(n1066), .A2(n1316), .ZN(n1241) );
NAND3_X1 U1028 ( .A1(n1119), .A2(n1230), .A3(G902), .ZN(n1316) );
NOR2_X1 U1029 ( .A1(G898), .A2(n1132), .ZN(n1119) );
NAND3_X1 U1030 ( .A1(n1034), .A2(n1230), .A3(G952), .ZN(n1066) );
NAND2_X1 U1031 ( .A1(G234), .A2(G237), .ZN(n1230) );
XNOR2_X1 U1032 ( .A(G953), .B(KEYINPUT16), .ZN(n1034) );
NAND2_X1 U1033 ( .A1(n1246), .A2(n1064), .ZN(n1061) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1251), .ZN(n1064) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1266), .ZN(n1251) );
XOR2_X1 U1036 ( .A(n1075), .B(G469), .Z(n1246) );
AND2_X1 U1037 ( .A1(n1317), .A2(n1266), .ZN(n1075) );
INV_X1 U1038 ( .A(G902), .ZN(n1266) );
XOR2_X1 U1039 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1040 ( .A(n1320), .B(n1171), .Z(n1319) );
XNOR2_X1 U1041 ( .A(n1321), .B(n1103), .ZN(n1171) );
XNOR2_X1 U1042 ( .A(n1322), .B(KEYINPUT60), .ZN(n1103) );
NAND2_X1 U1043 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1044 ( .A1(n1304), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1045 ( .A1(KEYINPUT19), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1046 ( .A1(G128), .A2(n1327), .ZN(n1326) );
NAND2_X1 U1047 ( .A1(n1328), .A2(n1302), .ZN(n1323) );
INV_X1 U1048 ( .A(G128), .ZN(n1302) );
NAND2_X1 U1049 ( .A1(n1327), .A2(n1329), .ZN(n1328) );
NAND2_X1 U1050 ( .A1(KEYINPUT19), .A2(n1273), .ZN(n1329) );
INV_X1 U1051 ( .A(n1304), .ZN(n1273) );
XOR2_X1 U1052 ( .A(n1215), .B(G146), .Z(n1304) );
INV_X1 U1053 ( .A(G143), .ZN(n1215) );
INV_X1 U1054 ( .A(KEYINPUT43), .ZN(n1327) );
NAND3_X1 U1055 ( .A1(n1330), .A2(n1331), .A3(n1313), .ZN(n1321) );
NAND3_X1 U1056 ( .A1(n1332), .A2(n1025), .A3(G101), .ZN(n1313) );
NAND2_X1 U1057 ( .A1(n1333), .A2(n1334), .ZN(n1331) );
INV_X1 U1058 ( .A(KEYINPUT31), .ZN(n1334) );
XOR2_X1 U1059 ( .A(G101), .B(n1335), .Z(n1333) );
NOR2_X1 U1060 ( .A1(n1332), .A2(n1025), .ZN(n1335) );
INV_X1 U1061 ( .A(G107), .ZN(n1025) );
NAND2_X1 U1062 ( .A1(KEYINPUT31), .A2(n1314), .ZN(n1330) );
NAND2_X1 U1063 ( .A1(n1336), .A2(n1337), .ZN(n1314) );
OR3_X1 U1064 ( .A1(n1332), .A2(G101), .A3(G107), .ZN(n1337) );
NAND2_X1 U1065 ( .A1(n1338), .A2(G107), .ZN(n1336) );
XOR2_X1 U1066 ( .A(G101), .B(n1332), .Z(n1338) );
XNOR2_X1 U1067 ( .A(n1151), .B(KEYINPUT55), .ZN(n1332) );
INV_X1 U1068 ( .A(G104), .ZN(n1151) );
NOR2_X1 U1069 ( .A1(KEYINPUT63), .A2(n1172), .ZN(n1320) );
XNOR2_X1 U1070 ( .A(n1339), .B(n1108), .ZN(n1172) );
XOR2_X1 U1071 ( .A(G134), .B(KEYINPUT9), .Z(n1108) );
XOR2_X1 U1072 ( .A(n1106), .B(KEYINPUT41), .Z(n1339) );
XOR2_X1 U1073 ( .A(n1223), .B(n1340), .Z(n1106) );
XOR2_X1 U1074 ( .A(KEYINPUT11), .B(G137), .Z(n1340) );
INV_X1 U1075 ( .A(G131), .ZN(n1223) );
XOR2_X1 U1076 ( .A(n1341), .B(n1342), .Z(n1318) );
XOR2_X1 U1077 ( .A(KEYINPUT54), .B(n1177), .Z(n1342) );
AND2_X1 U1078 ( .A1(G227), .A2(n1132), .ZN(n1177) );
INV_X1 U1079 ( .A(G953), .ZN(n1132) );
NOR2_X1 U1080 ( .A1(KEYINPUT12), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1081 ( .A(n1178), .B(G140), .Z(n1343) );
INV_X1 U1082 ( .A(G110), .ZN(n1178) );
endmodule


