//Key = 1000100010010001010100001001101010101110001100010110000011001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;

XNOR2_X1 U768 ( .A(n1061), .B(n1062), .ZN(G9) );
NOR3_X1 U769 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
INV_X1 U770 ( .A(n1066), .ZN(n1065) );
XOR2_X1 U771 ( .A(KEYINPUT11), .B(n1067), .Z(n1063) );
NOR2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(G75) );
NOR3_X1 U773 ( .A1(n1070), .A2(G953), .A3(n1071), .ZN(n1069) );
XOR2_X1 U774 ( .A(KEYINPUT43), .B(n1072), .Z(n1070) );
NOR3_X1 U775 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR3_X1 U779 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
AND2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR3_X1 U781 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
NOR3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(n1089), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1093), .A2(n1066), .ZN(n1092) );
INV_X1 U784 ( .A(n1094), .ZN(n1076) );
NOR4_X1 U785 ( .A1(n1095), .A2(n1089), .A3(n1091), .A4(n1082), .ZN(n1074) );
INV_X1 U786 ( .A(n1096), .ZN(n1082) );
INV_X1 U787 ( .A(n1086), .ZN(n1091) );
INV_X1 U788 ( .A(n1097), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XNOR2_X1 U791 ( .A(KEYINPUT54), .B(n1102), .ZN(n1101) );
NOR3_X1 U792 ( .A1(n1103), .A2(n1077), .A3(n1104), .ZN(n1098) );
NOR3_X1 U793 ( .A1(n1071), .A2(G953), .A3(G952), .ZN(n1068) );
AND4_X1 U794 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1071) );
NOR4_X1 U795 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
XNOR2_X1 U796 ( .A(KEYINPUT10), .B(n1113), .ZN(n1112) );
XNOR2_X1 U797 ( .A(G469), .B(n1114), .ZN(n1111) );
NAND2_X1 U798 ( .A1(KEYINPUT47), .A2(n1115), .ZN(n1114) );
NOR3_X1 U799 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1107) );
XOR2_X1 U800 ( .A(KEYINPUT39), .B(n1119), .Z(n1105) );
NOR3_X1 U801 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NOR3_X1 U802 ( .A1(n1123), .A2(KEYINPUT22), .A3(n1124), .ZN(n1122) );
AND2_X1 U803 ( .A1(n1123), .A2(KEYINPUT22), .ZN(n1121) );
INV_X1 U804 ( .A(n1125), .ZN(n1120) );
NAND3_X1 U805 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(G72) );
XOR2_X1 U806 ( .A(n1129), .B(KEYINPUT5), .Z(n1128) );
NAND2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND3_X1 U808 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1127) );
INV_X1 U809 ( .A(n1135), .ZN(n1134) );
OR2_X1 U810 ( .A1(n1131), .A2(n1130), .ZN(n1126) );
AND2_X1 U811 ( .A1(G953), .A2(n1136), .ZN(n1130) );
NAND2_X1 U812 ( .A1(G900), .A2(G227), .ZN(n1136) );
NAND3_X1 U813 ( .A1(n1135), .A2(n1137), .A3(n1138), .ZN(n1131) );
XOR2_X1 U814 ( .A(n1139), .B(KEYINPUT26), .Z(n1138) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1132), .ZN(n1139) );
NAND3_X1 U816 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1143), .B(KEYINPUT59), .Z(n1142) );
OR2_X1 U818 ( .A1(n1133), .A2(G900), .ZN(n1137) );
XNOR2_X1 U819 ( .A(n1144), .B(n1145), .ZN(n1135) );
XNOR2_X1 U820 ( .A(n1146), .B(n1147), .ZN(n1145) );
INV_X1 U821 ( .A(n1148), .ZN(n1146) );
XNOR2_X1 U822 ( .A(G131), .B(n1149), .ZN(n1144) );
NOR2_X1 U823 ( .A1(KEYINPUT29), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U824 ( .A(G137), .B(n1151), .ZN(n1150) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(G69) );
XOR2_X1 U826 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U827 ( .A1(G953), .A2(n1156), .ZN(n1155) );
XOR2_X1 U828 ( .A(KEYINPUT48), .B(n1157), .Z(n1156) );
NAND2_X1 U829 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
INV_X1 U830 ( .A(n1160), .ZN(n1159) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1158) );
XNOR2_X1 U832 ( .A(n1163), .B(n1164), .ZN(n1162) );
NAND2_X1 U833 ( .A1(KEYINPUT19), .A2(n1165), .ZN(n1164) );
NOR2_X1 U834 ( .A1(KEYINPUT23), .A2(n1166), .ZN(n1161) );
NAND2_X1 U835 ( .A1(G953), .A2(n1167), .ZN(n1152) );
NAND2_X1 U836 ( .A1(G898), .A2(G224), .ZN(n1167) );
NOR2_X1 U837 ( .A1(n1168), .A2(n1169), .ZN(G66) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1168), .A2(n1174), .ZN(G63) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND3_X1 U842 ( .A1(n1177), .A2(G478), .A3(KEYINPUT4), .ZN(n1175) );
NOR2_X1 U843 ( .A1(n1168), .A2(n1178), .ZN(G60) );
XOR2_X1 U844 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U845 ( .A1(n1123), .A2(n1173), .ZN(n1179) );
XNOR2_X1 U846 ( .A(G104), .B(n1181), .ZN(G6) );
NOR2_X1 U847 ( .A1(n1168), .A2(n1182), .ZN(G57) );
XOR2_X1 U848 ( .A(n1183), .B(n1184), .Z(n1182) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(n1184) );
AND2_X1 U850 ( .A1(G472), .A2(n1177), .ZN(n1185) );
INV_X1 U851 ( .A(n1173), .ZN(n1177) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1183) );
XNOR2_X1 U853 ( .A(G101), .B(n1189), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1168), .A2(n1190), .ZN(G54) );
XOR2_X1 U855 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U856 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U857 ( .A1(n1195), .A2(n1173), .ZN(n1194) );
NOR3_X1 U858 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U860 ( .A(n1201), .ZN(n1200) );
NOR2_X1 U861 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
XOR2_X1 U862 ( .A(n1204), .B(KEYINPUT16), .Z(n1202) );
NOR3_X1 U863 ( .A1(n1201), .A2(n1204), .A3(n1203), .ZN(n1197) );
AND2_X1 U864 ( .A1(n1203), .A2(n1204), .ZN(n1196) );
NAND3_X1 U865 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1204) );
OR2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U867 ( .A1(KEYINPUT2), .A2(n1210), .ZN(n1206) );
NAND2_X1 U868 ( .A1(n1211), .A2(n1209), .ZN(n1210) );
XNOR2_X1 U869 ( .A(KEYINPUT50), .B(n1208), .ZN(n1211) );
NAND2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1205) );
INV_X1 U871 ( .A(KEYINPUT2), .ZN(n1213) );
NAND2_X1 U872 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
OR2_X1 U873 ( .A1(n1208), .A2(KEYINPUT50), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1208), .A2(n1209), .A3(KEYINPUT50), .ZN(n1214) );
XOR2_X1 U875 ( .A(n1148), .B(KEYINPUT33), .Z(n1208) );
INV_X1 U876 ( .A(KEYINPUT56), .ZN(n1203) );
NOR2_X1 U877 ( .A1(KEYINPUT13), .A2(n1216), .ZN(n1191) );
NOR2_X1 U878 ( .A1(n1168), .A2(n1217), .ZN(G51) );
XOR2_X1 U879 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U880 ( .A(n1220), .B(n1221), .Z(n1218) );
NOR2_X1 U881 ( .A1(n1222), .A2(n1173), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1223), .A2(n1073), .ZN(n1173) );
NAND4_X1 U883 ( .A1(n1157), .A2(n1140), .A3(n1224), .A4(n1143), .ZN(n1073) );
XNOR2_X1 U884 ( .A(KEYINPUT28), .B(n1141), .ZN(n1224) );
AND3_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1140) );
NOR3_X1 U886 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
INV_X1 U887 ( .A(n1231), .ZN(n1228) );
NAND2_X1 U888 ( .A1(n1094), .A2(n1232), .ZN(n1225) );
NAND2_X1 U889 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U890 ( .A(n1235), .B(KEYINPUT40), .Z(n1234) );
NAND3_X1 U891 ( .A1(n1096), .A2(n1236), .A3(n1237), .ZN(n1235) );
XOR2_X1 U892 ( .A(KEYINPUT51), .B(n1238), .Z(n1236) );
XNOR2_X1 U893 ( .A(n1239), .B(KEYINPUT3), .ZN(n1233) );
AND4_X1 U894 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1157) );
AND4_X1 U895 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1181), .ZN(n1243) );
NAND3_X1 U896 ( .A1(n1247), .A2(n1067), .A3(n1093), .ZN(n1181) );
NAND3_X1 U897 ( .A1(n1248), .A2(n1083), .A3(n1066), .ZN(n1242) );
NAND2_X1 U898 ( .A1(n1249), .A2(n1250), .ZN(n1083) );
NAND2_X1 U899 ( .A1(n1067), .A2(n1097), .ZN(n1250) );
NAND2_X1 U900 ( .A1(n1251), .A2(n1086), .ZN(n1249) );
NAND2_X1 U901 ( .A1(n1252), .A2(n1253), .ZN(n1241) );
NAND2_X1 U902 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U903 ( .A1(n1067), .A2(n1256), .A3(n1251), .ZN(n1255) );
INV_X1 U904 ( .A(KEYINPUT44), .ZN(n1256) );
NAND2_X1 U905 ( .A1(KEYINPUT17), .A2(n1257), .ZN(n1254) );
INV_X1 U906 ( .A(n1258), .ZN(n1257) );
NAND4_X1 U907 ( .A1(n1096), .A2(n1259), .A3(n1260), .A4(n1100), .ZN(n1240) );
NAND2_X1 U908 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
NAND3_X1 U909 ( .A1(n1251), .A2(n1067), .A3(KEYINPUT44), .ZN(n1262) );
OR2_X1 U910 ( .A1(n1258), .A2(KEYINPUT17), .ZN(n1261) );
XNOR2_X1 U911 ( .A(KEYINPUT25), .B(n1263), .ZN(n1223) );
NAND3_X1 U912 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1220) );
NAND2_X1 U913 ( .A1(KEYINPUT41), .A2(n1267), .ZN(n1265) );
NAND3_X1 U914 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
INV_X1 U915 ( .A(n1271), .ZN(n1270) );
NAND2_X1 U916 ( .A1(G125), .A2(n1272), .ZN(n1269) );
NAND3_X1 U917 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1268) );
OR2_X1 U918 ( .A1(n1276), .A2(KEYINPUT41), .ZN(n1264) );
NOR2_X1 U919 ( .A1(n1133), .A2(G952), .ZN(n1168) );
XOR2_X1 U920 ( .A(n1226), .B(n1277), .Z(G48) );
XOR2_X1 U921 ( .A(KEYINPUT24), .B(G146), .Z(n1277) );
NAND3_X1 U922 ( .A1(n1093), .A2(n1278), .A3(n1279), .ZN(n1226) );
XNOR2_X1 U923 ( .A(G143), .B(n1141), .ZN(G45) );
NAND4_X1 U924 ( .A1(n1237), .A2(n1251), .A3(n1280), .A4(n1278), .ZN(n1141) );
NOR2_X1 U925 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XNOR2_X1 U926 ( .A(G140), .B(n1283), .ZN(G42) );
NAND3_X1 U927 ( .A1(n1239), .A2(n1094), .A3(KEYINPUT15), .ZN(n1283) );
AND3_X1 U928 ( .A1(n1093), .A2(n1087), .A3(n1237), .ZN(n1239) );
XOR2_X1 U929 ( .A(n1284), .B(n1285), .Z(G39) );
NAND3_X1 U930 ( .A1(n1279), .A2(n1096), .A3(n1094), .ZN(n1285) );
NAND2_X1 U931 ( .A1(KEYINPUT8), .A2(G137), .ZN(n1284) );
XNOR2_X1 U932 ( .A(n1151), .B(n1230), .ZN(G36) );
AND2_X1 U933 ( .A1(n1286), .A2(n1066), .ZN(n1230) );
XNOR2_X1 U934 ( .A(n1287), .B(n1229), .ZN(G33) );
AND2_X1 U935 ( .A1(n1286), .A2(n1093), .ZN(n1229) );
AND3_X1 U936 ( .A1(n1237), .A2(n1251), .A3(n1094), .ZN(n1286) );
NOR2_X1 U937 ( .A1(n1104), .A2(n1116), .ZN(n1094) );
XNOR2_X1 U938 ( .A(G128), .B(n1143), .ZN(G30) );
NAND3_X1 U939 ( .A1(n1066), .A2(n1278), .A3(n1279), .ZN(n1143) );
AND2_X1 U940 ( .A1(n1237), .A2(n1238), .ZN(n1279) );
AND2_X1 U941 ( .A1(n1067), .A2(n1288), .ZN(n1237) );
OR2_X1 U942 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U943 ( .A(G101), .B(n1291), .ZN(G3) );
NAND2_X1 U944 ( .A1(n1251), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U945 ( .A(G125), .B(n1231), .ZN(G27) );
NAND4_X1 U946 ( .A1(n1093), .A2(n1087), .A3(n1293), .A4(n1086), .ZN(n1231) );
NOR2_X1 U947 ( .A1(n1294), .A2(n1100), .ZN(n1293) );
NOR2_X1 U948 ( .A1(n1289), .A2(n1290), .ZN(n1294) );
NOR4_X1 U949 ( .A1(n1263), .A2(n1133), .A3(n1077), .A4(G900), .ZN(n1290) );
INV_X1 U950 ( .A(n1102), .ZN(n1077) );
INV_X1 U951 ( .A(n1295), .ZN(n1289) );
XOR2_X1 U952 ( .A(n1246), .B(n1296), .Z(G24) );
XNOR2_X1 U953 ( .A(KEYINPUT63), .B(n1297), .ZN(n1296) );
NAND4_X1 U954 ( .A1(n1086), .A2(n1247), .A3(n1110), .A4(n1298), .ZN(n1246) );
INV_X1 U955 ( .A(n1064), .ZN(n1247) );
NAND2_X1 U956 ( .A1(n1248), .A2(n1097), .ZN(n1064) );
NOR2_X1 U957 ( .A1(n1299), .A2(n1109), .ZN(n1097) );
XNOR2_X1 U958 ( .A(G119), .B(n1300), .ZN(G21) );
NOR2_X1 U959 ( .A1(KEYINPUT58), .A2(n1301), .ZN(n1300) );
NOR2_X1 U960 ( .A1(n1302), .A2(n1258), .ZN(n1301) );
NAND2_X1 U961 ( .A1(n1238), .A2(n1086), .ZN(n1258) );
NOR2_X1 U962 ( .A1(n1303), .A2(n1304), .ZN(n1238) );
XNOR2_X1 U963 ( .A(G116), .B(n1305), .ZN(G18) );
NAND4_X1 U964 ( .A1(n1306), .A2(n1260), .A3(n1066), .A4(n1307), .ZN(n1305) );
AND2_X1 U965 ( .A1(n1086), .A2(n1251), .ZN(n1307) );
NOR2_X1 U966 ( .A1(n1298), .A2(n1282), .ZN(n1066) );
INV_X1 U967 ( .A(n1110), .ZN(n1282) );
XNOR2_X1 U968 ( .A(KEYINPUT20), .B(n1100), .ZN(n1306) );
INV_X1 U969 ( .A(n1278), .ZN(n1100) );
XNOR2_X1 U970 ( .A(G113), .B(n1245), .ZN(G15) );
NAND4_X1 U971 ( .A1(n1093), .A2(n1251), .A3(n1086), .A4(n1248), .ZN(n1245) );
NOR2_X1 U972 ( .A1(n1090), .A2(n1118), .ZN(n1086) );
INV_X1 U973 ( .A(n1088), .ZN(n1118) );
NOR2_X1 U974 ( .A1(n1299), .A2(n1303), .ZN(n1251) );
INV_X1 U975 ( .A(n1109), .ZN(n1303) );
NOR2_X1 U976 ( .A1(n1110), .A2(n1281), .ZN(n1093) );
INV_X1 U977 ( .A(n1298), .ZN(n1281) );
XNOR2_X1 U978 ( .A(G110), .B(n1244), .ZN(G12) );
NAND2_X1 U979 ( .A1(n1292), .A2(n1087), .ZN(n1244) );
NOR2_X1 U980 ( .A1(n1109), .A2(n1304), .ZN(n1087) );
INV_X1 U981 ( .A(n1299), .ZN(n1304) );
NAND3_X1 U982 ( .A1(n1308), .A2(n1309), .A3(n1106), .ZN(n1299) );
NAND2_X1 U983 ( .A1(n1310), .A2(n1311), .ZN(n1106) );
NAND2_X1 U984 ( .A1(n1117), .A2(KEYINPUT61), .ZN(n1309) );
NOR2_X1 U985 ( .A1(n1311), .A2(n1310), .ZN(n1117) );
INV_X1 U986 ( .A(n1172), .ZN(n1310) );
NAND2_X1 U987 ( .A1(G217), .A2(n1312), .ZN(n1172) );
INV_X1 U988 ( .A(n1313), .ZN(n1311) );
OR2_X1 U989 ( .A1(n1313), .A2(KEYINPUT61), .ZN(n1308) );
NOR2_X1 U990 ( .A1(n1171), .A2(G902), .ZN(n1313) );
XNOR2_X1 U991 ( .A(n1314), .B(n1315), .ZN(n1171) );
XOR2_X1 U992 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U993 ( .A(n1147), .B(n1318), .ZN(n1317) );
NOR2_X1 U994 ( .A1(G146), .A2(KEYINPUT46), .ZN(n1318) );
XNOR2_X1 U995 ( .A(G140), .B(n1274), .ZN(n1147) );
NAND2_X1 U996 ( .A1(n1319), .A2(n1320), .ZN(n1316) );
NAND2_X1 U997 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U998 ( .A(KEYINPUT14), .B(n1323), .Z(n1321) );
NAND2_X1 U999 ( .A1(G110), .A2(n1324), .ZN(n1319) );
XNOR2_X1 U1000 ( .A(n1323), .B(KEYINPUT1), .ZN(n1324) );
XOR2_X1 U1001 ( .A(G119), .B(G128), .Z(n1323) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1314) );
XOR2_X1 U1003 ( .A(KEYINPUT0), .B(G137), .Z(n1326) );
NAND2_X1 U1004 ( .A1(G221), .A2(n1327), .ZN(n1325) );
XNOR2_X1 U1005 ( .A(n1328), .B(G472), .ZN(n1109) );
NAND3_X1 U1006 ( .A1(n1329), .A2(n1263), .A3(n1330), .ZN(n1328) );
NAND3_X1 U1007 ( .A1(n1189), .A2(n1331), .A3(n1332), .ZN(n1330) );
XNOR2_X1 U1008 ( .A(n1333), .B(n1334), .ZN(n1332) );
NAND2_X1 U1009 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
OR2_X1 U1010 ( .A1(n1186), .A2(KEYINPUT49), .ZN(n1336) );
OR2_X1 U1011 ( .A1(n1337), .A2(KEYINPUT18), .ZN(n1335) );
NAND2_X1 U1012 ( .A1(n1338), .A2(n1339), .ZN(n1329) );
NAND2_X1 U1013 ( .A1(n1189), .A2(n1331), .ZN(n1339) );
INV_X1 U1014 ( .A(KEYINPUT21), .ZN(n1331) );
NAND2_X1 U1015 ( .A1(n1340), .A2(n1341), .ZN(n1189) );
NAND2_X1 U1016 ( .A1(G113), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1017 ( .A(n1343), .B(n1344), .ZN(n1338) );
INV_X1 U1018 ( .A(n1334), .ZN(n1344) );
XOR2_X1 U1019 ( .A(n1345), .B(n1187), .Z(n1334) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1346), .ZN(n1187) );
NAND2_X1 U1021 ( .A1(KEYINPUT60), .A2(n1347), .ZN(n1345) );
INV_X1 U1022 ( .A(G101), .ZN(n1347) );
NAND2_X1 U1023 ( .A1(n1348), .A2(n1349), .ZN(n1343) );
NAND2_X1 U1024 ( .A1(n1186), .A2(KEYINPUT49), .ZN(n1349) );
INV_X1 U1025 ( .A(n1337), .ZN(n1186) );
NAND2_X1 U1026 ( .A1(n1337), .A2(KEYINPUT18), .ZN(n1348) );
XNOR2_X1 U1027 ( .A(n1350), .B(n1273), .ZN(n1337) );
XNOR2_X1 U1028 ( .A(n1201), .B(KEYINPUT30), .ZN(n1350) );
AND2_X1 U1029 ( .A1(n1252), .A2(n1067), .ZN(n1292) );
AND2_X1 U1030 ( .A1(n1090), .A2(n1088), .ZN(n1067) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1312), .ZN(n1088) );
NAND2_X1 U1032 ( .A1(G234), .A2(n1263), .ZN(n1312) );
XNOR2_X1 U1033 ( .A(n1115), .B(n1195), .ZN(n1090) );
INV_X1 U1034 ( .A(G469), .ZN(n1195) );
AND2_X1 U1035 ( .A1(n1351), .A2(n1263), .ZN(n1115) );
XOR2_X1 U1036 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1037 ( .A(n1209), .B(n1216), .ZN(n1353) );
XNOR2_X1 U1038 ( .A(n1354), .B(n1355), .ZN(n1216) );
XNOR2_X1 U1039 ( .A(G140), .B(n1322), .ZN(n1355) );
NAND2_X1 U1040 ( .A1(G227), .A2(n1133), .ZN(n1354) );
XNOR2_X1 U1041 ( .A(n1356), .B(n1357), .ZN(n1209) );
NOR2_X1 U1042 ( .A1(KEYINPUT55), .A2(n1061), .ZN(n1357) );
XNOR2_X1 U1043 ( .A(n1201), .B(n1358), .ZN(n1352) );
NOR2_X1 U1044 ( .A1(KEYINPUT53), .A2(n1148), .ZN(n1358) );
XNOR2_X1 U1045 ( .A(n1359), .B(G128), .ZN(n1148) );
NAND2_X1 U1046 ( .A1(KEYINPUT57), .A2(n1360), .ZN(n1359) );
NAND2_X1 U1047 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1048 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XNOR2_X1 U1049 ( .A(G143), .B(KEYINPUT12), .ZN(n1364) );
XNOR2_X1 U1050 ( .A(G146), .B(KEYINPUT27), .ZN(n1363) );
XOR2_X1 U1051 ( .A(KEYINPUT42), .B(n1365), .Z(n1361) );
NOR2_X1 U1052 ( .A1(G146), .A2(n1366), .ZN(n1365) );
XNOR2_X1 U1053 ( .A(n1367), .B(n1368), .ZN(n1201) );
XNOR2_X1 U1054 ( .A(G137), .B(n1287), .ZN(n1368) );
NAND2_X1 U1055 ( .A1(KEYINPUT36), .A2(n1151), .ZN(n1367) );
INV_X1 U1056 ( .A(n1302), .ZN(n1252) );
NAND2_X1 U1057 ( .A1(n1096), .A2(n1248), .ZN(n1302) );
AND2_X1 U1058 ( .A1(n1278), .A2(n1260), .ZN(n1248) );
NAND2_X1 U1059 ( .A1(n1295), .A2(n1369), .ZN(n1260) );
NAND3_X1 U1060 ( .A1(n1160), .A2(n1102), .A3(G902), .ZN(n1369) );
NOR2_X1 U1061 ( .A1(n1133), .A2(G898), .ZN(n1160) );
NAND3_X1 U1062 ( .A1(G952), .A2(n1102), .A3(n1370), .ZN(n1295) );
XNOR2_X1 U1063 ( .A(G953), .B(KEYINPUT9), .ZN(n1370) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1102) );
NOR2_X1 U1065 ( .A1(n1113), .A2(n1116), .ZN(n1278) );
INV_X1 U1066 ( .A(n1103), .ZN(n1116) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1371), .ZN(n1103) );
INV_X1 U1068 ( .A(n1104), .ZN(n1113) );
XOR2_X1 U1069 ( .A(n1372), .B(n1222), .Z(n1104) );
NAND2_X1 U1070 ( .A1(G210), .A2(n1371), .ZN(n1222) );
NAND2_X1 U1071 ( .A1(n1373), .A2(n1263), .ZN(n1371) );
INV_X1 U1072 ( .A(G237), .ZN(n1373) );
NAND2_X1 U1073 ( .A1(n1374), .A2(n1263), .ZN(n1372) );
XOR2_X1 U1074 ( .A(n1375), .B(n1376), .Z(n1374) );
NOR2_X1 U1075 ( .A1(KEYINPUT31), .A2(n1219), .ZN(n1376) );
XOR2_X1 U1076 ( .A(n1377), .B(n1166), .Z(n1219) );
XNOR2_X1 U1077 ( .A(n1378), .B(n1322), .ZN(n1166) );
INV_X1 U1078 ( .A(G110), .ZN(n1322) );
NAND2_X1 U1079 ( .A1(KEYINPUT32), .A2(n1297), .ZN(n1378) );
XOR2_X1 U1080 ( .A(n1165), .B(n1379), .Z(n1377) );
NOR2_X1 U1081 ( .A1(n1163), .A2(KEYINPUT35), .ZN(n1379) );
AND2_X1 U1082 ( .A1(n1380), .A2(n1341), .ZN(n1163) );
OR2_X1 U1083 ( .A1(n1342), .A2(G113), .ZN(n1341) );
NAND2_X1 U1084 ( .A1(n1381), .A2(n1342), .ZN(n1380) );
XOR2_X1 U1085 ( .A(G116), .B(G119), .Z(n1342) );
XNOR2_X1 U1086 ( .A(G113), .B(KEYINPUT37), .ZN(n1381) );
XOR2_X1 U1087 ( .A(n1356), .B(n1382), .Z(n1165) );
XNOR2_X1 U1088 ( .A(KEYINPUT34), .B(n1061), .ZN(n1382) );
XNOR2_X1 U1089 ( .A(G101), .B(n1383), .ZN(n1356) );
XOR2_X1 U1090 ( .A(KEYINPUT52), .B(G104), .Z(n1383) );
NAND2_X1 U1091 ( .A1(n1276), .A2(n1266), .ZN(n1375) );
NAND2_X1 U1092 ( .A1(n1271), .A2(G125), .ZN(n1266) );
NOR2_X1 U1093 ( .A1(n1273), .A2(n1275), .ZN(n1271) );
AND2_X1 U1094 ( .A1(n1384), .A2(n1385), .ZN(n1276) );
NAND2_X1 U1095 ( .A1(n1386), .A2(n1274), .ZN(n1385) );
XNOR2_X1 U1096 ( .A(n1272), .B(n1273), .ZN(n1386) );
NAND3_X1 U1097 ( .A1(n1275), .A2(n1273), .A3(G125), .ZN(n1384) );
XNOR2_X1 U1098 ( .A(n1387), .B(n1388), .ZN(n1273) );
XNOR2_X1 U1099 ( .A(G146), .B(KEYINPUT7), .ZN(n1387) );
INV_X1 U1100 ( .A(n1272), .ZN(n1275) );
NAND2_X1 U1101 ( .A1(G224), .A2(n1133), .ZN(n1272) );
NOR2_X1 U1102 ( .A1(n1110), .A2(n1298), .ZN(n1096) );
NAND2_X1 U1103 ( .A1(n1389), .A2(n1125), .ZN(n1298) );
NAND2_X1 U1104 ( .A1(n1124), .A2(n1123), .ZN(n1125) );
OR2_X1 U1105 ( .A1(n1123), .A2(n1124), .ZN(n1389) );
NOR2_X1 U1106 ( .A1(n1180), .A2(G902), .ZN(n1124) );
XNOR2_X1 U1107 ( .A(n1390), .B(n1391), .ZN(n1180) );
XOR2_X1 U1108 ( .A(n1392), .B(n1393), .Z(n1391) );
XNOR2_X1 U1109 ( .A(n1394), .B(n1395), .ZN(n1393) );
NOR2_X1 U1110 ( .A1(KEYINPUT6), .A2(n1396), .ZN(n1395) );
NOR2_X1 U1111 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1399), .Z(n1398) );
NOR2_X1 U1113 ( .A1(n1400), .A2(n1287), .ZN(n1399) );
AND2_X1 U1114 ( .A1(n1287), .A2(n1400), .ZN(n1397) );
XOR2_X1 U1115 ( .A(n1401), .B(n1366), .Z(n1400) );
NAND2_X1 U1116 ( .A1(G214), .A2(n1346), .ZN(n1401) );
NOR2_X1 U1117 ( .A1(G953), .A2(G237), .ZN(n1346) );
INV_X1 U1118 ( .A(G131), .ZN(n1287) );
NAND2_X1 U1119 ( .A1(KEYINPUT38), .A2(n1402), .ZN(n1394) );
XNOR2_X1 U1120 ( .A(n1297), .B(G113), .ZN(n1402) );
INV_X1 U1121 ( .A(G122), .ZN(n1297) );
NOR2_X1 U1122 ( .A1(G140), .A2(KEYINPUT45), .ZN(n1392) );
XNOR2_X1 U1123 ( .A(G104), .B(n1403), .ZN(n1390) );
XNOR2_X1 U1124 ( .A(G146), .B(n1274), .ZN(n1403) );
INV_X1 U1125 ( .A(G125), .ZN(n1274) );
INV_X1 U1126 ( .A(G475), .ZN(n1123) );
XNOR2_X1 U1127 ( .A(n1404), .B(G478), .ZN(n1110) );
NAND2_X1 U1128 ( .A1(n1176), .A2(n1263), .ZN(n1404) );
INV_X1 U1129 ( .A(G902), .ZN(n1263) );
XNOR2_X1 U1130 ( .A(n1405), .B(n1406), .ZN(n1176) );
XOR2_X1 U1131 ( .A(G116), .B(n1407), .Z(n1406) );
XNOR2_X1 U1132 ( .A(n1151), .B(G122), .ZN(n1407) );
INV_X1 U1133 ( .A(G134), .ZN(n1151) );
XOR2_X1 U1134 ( .A(n1408), .B(n1388), .Z(n1405) );
XNOR2_X1 U1135 ( .A(G128), .B(n1366), .ZN(n1388) );
INV_X1 U1136 ( .A(G143), .ZN(n1366) );
XNOR2_X1 U1137 ( .A(n1409), .B(n1061), .ZN(n1408) );
INV_X1 U1138 ( .A(G107), .ZN(n1061) );
NAND2_X1 U1139 ( .A1(G217), .A2(n1327), .ZN(n1409) );
AND2_X1 U1140 ( .A1(G234), .A2(n1133), .ZN(n1327) );
INV_X1 U1141 ( .A(G953), .ZN(n1133) );
endmodule


