//Key = 0001111111000001011001000000000110110011010101101000101101110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;

XNOR2_X1 U726 ( .A(n1001), .B(n1002), .ZN(G9) );
NOR2_X1 U727 ( .A1(KEYINPUT1), .A2(n1003), .ZN(n1002) );
INV_X1 U728 ( .A(G107), .ZN(n1003) );
NOR2_X1 U729 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR3_X1 U730 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
NOR2_X1 U731 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U732 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U733 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
INV_X1 U734 ( .A(n1015), .ZN(n1014) );
NOR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1013) );
NOR2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U738 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U740 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
XNOR2_X1 U741 ( .A(n1028), .B(KEYINPUT60), .ZN(n1026) );
NOR2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(n1020) );
NOR2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U745 ( .A1(n1030), .A2(n1035), .A3(n1023), .ZN(n1016) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR4_X1 U748 ( .A1(n1040), .A2(n1023), .A3(n1019), .A4(n1030), .ZN(n1011) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U750 ( .A1(G952), .A2(n1008), .ZN(n1004) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1008) );
NAND4_X1 U752 ( .A1(n1045), .A2(n1033), .A3(n1046), .A4(n1047), .ZN(n1044) );
NOR4_X1 U753 ( .A1(n1028), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1047) );
XOR2_X1 U754 ( .A(n1051), .B(n1052), .Z(n1049) );
NOR2_X1 U755 ( .A1(n1053), .A2(KEYINPUT2), .ZN(n1052) );
NOR3_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1048) );
NOR2_X1 U757 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR3_X1 U758 ( .A1(G478), .A2(KEYINPUT44), .A3(n1059), .ZN(n1055) );
INV_X1 U759 ( .A(n1057), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1060), .A2(KEYINPUT22), .ZN(n1057) );
AND2_X1 U761 ( .A1(n1060), .A2(KEYINPUT44), .ZN(n1054) );
XOR2_X1 U762 ( .A(n1061), .B(n1062), .Z(G72) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XOR2_X1 U765 ( .A(KEYINPUT20), .B(n1067), .Z(n1066) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XOR2_X1 U767 ( .A(KEYINPUT13), .B(n1043), .Z(n1065) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1063) );
XOR2_X1 U769 ( .A(KEYINPUT21), .B(G953), .Z(n1070) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1061) );
NAND2_X1 U771 ( .A1(G953), .A2(n1069), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1074), .B(n1075), .Z(n1072) );
NAND2_X1 U773 ( .A1(n1076), .A2(KEYINPUT46), .ZN(n1074) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(G69) );
XOR2_X1 U776 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U778 ( .A1(G898), .A2(G224), .ZN(n1084) );
XOR2_X1 U779 ( .A(KEYINPUT13), .B(G953), .Z(n1083) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1087), .B(KEYINPUT24), .Z(n1085) );
NAND2_X1 U782 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NOR3_X1 U783 ( .A1(n1089), .A2(KEYINPUT23), .A3(G953), .ZN(n1079) );
INV_X1 U784 ( .A(n1090), .ZN(n1089) );
NOR3_X1 U785 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(G66) );
NOR3_X1 U786 ( .A1(n1094), .A2(G953), .A3(G952), .ZN(n1093) );
AND2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
INV_X1 U788 ( .A(KEYINPUT30), .ZN(n1094) );
XOR2_X1 U789 ( .A(n1096), .B(n1097), .Z(n1091) );
NAND3_X1 U790 ( .A1(n1098), .A2(G217), .A3(KEYINPUT8), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1099), .ZN(G63) );
NOR3_X1 U792 ( .A1(n1060), .A2(n1100), .A3(n1101), .ZN(n1099) );
AND3_X1 U793 ( .A1(n1102), .A2(G478), .A3(n1098), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1103), .A2(n1102), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1104), .A2(n1058), .ZN(n1103) );
INV_X1 U796 ( .A(G478), .ZN(n1058) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1106), .ZN(G60) );
XOR2_X1 U798 ( .A(n1107), .B(KEYINPUT54), .Z(n1106) );
NAND2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U800 ( .A(n1043), .B(KEYINPUT31), .Z(n1108) );
NOR2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
XOR2_X1 U802 ( .A(n1112), .B(KEYINPUT17), .Z(n1111) );
NAND2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XNOR2_X1 U805 ( .A(n1115), .B(KEYINPUT42), .ZN(n1114) );
AND2_X1 U806 ( .A1(n1098), .A2(G475), .ZN(n1113) );
XNOR2_X1 U807 ( .A(G104), .B(n1116), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1095), .A2(n1117), .ZN(G57) );
XOR2_X1 U809 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U810 ( .A(n1078), .B(n1120), .ZN(n1118) );
AND2_X1 U811 ( .A1(G472), .A2(n1098), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1095), .A2(n1121), .ZN(G54) );
XOR2_X1 U813 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U814 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U815 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U816 ( .A1(n1128), .A2(KEYINPUT32), .ZN(n1127) );
XOR2_X1 U817 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U818 ( .A1(KEYINPUT41), .A2(G110), .ZN(n1129) );
NAND3_X1 U819 ( .A1(n1131), .A2(n1006), .A3(G469), .ZN(n1126) );
INV_X1 U820 ( .A(n1104), .ZN(n1006) );
XOR2_X1 U821 ( .A(KEYINPUT56), .B(G902), .Z(n1131) );
NOR2_X1 U822 ( .A1(KEYINPUT14), .A2(n1077), .ZN(n1124) );
XNOR2_X1 U823 ( .A(n1078), .B(n1132), .ZN(n1122) );
NOR2_X1 U824 ( .A1(n1095), .A2(n1133), .ZN(G51) );
NOR3_X1 U825 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR2_X1 U826 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
INV_X1 U827 ( .A(n1139), .ZN(n1138) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
XOR2_X1 U829 ( .A(n1142), .B(KEYINPUT27), .Z(n1140) );
NOR3_X1 U830 ( .A1(n1139), .A2(n1142), .A3(n1141), .ZN(n1135) );
XNOR2_X1 U831 ( .A(n1143), .B(n1086), .ZN(n1139) );
NAND2_X1 U832 ( .A1(n1144), .A2(KEYINPUT35), .ZN(n1143) );
XOR2_X1 U833 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U834 ( .A1(KEYINPUT12), .A2(n1147), .ZN(n1146) );
AND2_X1 U835 ( .A1(n1141), .A2(n1142), .ZN(n1134) );
NAND2_X1 U836 ( .A1(n1098), .A2(n1053), .ZN(n1142) );
NOR2_X1 U837 ( .A1(n1148), .A2(n1104), .ZN(n1098) );
NOR2_X1 U838 ( .A1(n1090), .A2(n1071), .ZN(n1104) );
NAND2_X1 U839 ( .A1(n1149), .A2(n1150), .ZN(n1071) );
NOR4_X1 U840 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NOR4_X1 U841 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1149) );
NOR3_X1 U842 ( .A1(n1159), .A2(n1019), .A3(n1160), .ZN(n1158) );
XOR2_X1 U843 ( .A(KEYINPUT4), .B(n1025), .Z(n1159) );
INV_X1 U844 ( .A(n1161), .ZN(n1155) );
NAND2_X1 U845 ( .A1(n1162), .A2(n1163), .ZN(n1090) );
AND4_X1 U846 ( .A1(n1164), .A2(n1165), .A3(n1001), .A4(n1166), .ZN(n1163) );
NAND3_X1 U847 ( .A1(n1167), .A2(n1168), .A3(n1042), .ZN(n1001) );
AND4_X1 U848 ( .A1(n1169), .A2(n1170), .A3(n1116), .A4(n1171), .ZN(n1162) );
NAND3_X1 U849 ( .A1(n1041), .A2(n1172), .A3(n1032), .ZN(n1171) );
NAND3_X1 U850 ( .A1(n1167), .A2(n1168), .A3(n1041), .ZN(n1116) );
INV_X1 U851 ( .A(KEYINPUT45), .ZN(n1141) );
NOR2_X1 U852 ( .A1(n1043), .A2(G952), .ZN(n1095) );
XOR2_X1 U853 ( .A(n1173), .B(n1161), .Z(G48) );
NAND4_X1 U854 ( .A1(n1174), .A2(n1041), .A3(n1025), .A4(n1037), .ZN(n1161) );
XNOR2_X1 U855 ( .A(n1157), .B(n1175), .ZN(G45) );
NAND2_X1 U856 ( .A1(KEYINPUT3), .A2(G143), .ZN(n1175) );
AND4_X1 U857 ( .A1(n1025), .A2(n1037), .A3(n1032), .A4(n1176), .ZN(n1157) );
AND3_X1 U858 ( .A1(n1177), .A2(n1178), .A3(n1050), .ZN(n1176) );
XOR2_X1 U859 ( .A(G140), .B(n1156), .Z(G42) );
NOR3_X1 U860 ( .A1(n1030), .A2(n1179), .A3(n1160), .ZN(n1156) );
INV_X1 U861 ( .A(n1037), .ZN(n1179) );
NAND2_X1 U862 ( .A1(n1180), .A2(n1181), .ZN(G39) );
NAND2_X1 U863 ( .A1(n1154), .A2(n1182), .ZN(n1181) );
XOR2_X1 U864 ( .A(KEYINPUT18), .B(n1183), .Z(n1180) );
NOR2_X1 U865 ( .A1(n1154), .A2(n1182), .ZN(n1183) );
INV_X1 U866 ( .A(G137), .ZN(n1182) );
AND4_X1 U867 ( .A1(n1184), .A2(n1174), .A3(n1037), .A4(n1015), .ZN(n1154) );
XOR2_X1 U868 ( .A(G134), .B(n1153), .Z(G36) );
AND2_X1 U869 ( .A1(n1185), .A2(n1042), .ZN(n1153) );
NAND2_X1 U870 ( .A1(n1186), .A2(n1187), .ZN(G33) );
NAND2_X1 U871 ( .A1(n1152), .A2(n1188), .ZN(n1187) );
XOR2_X1 U872 ( .A(KEYINPUT6), .B(n1189), .Z(n1186) );
NOR2_X1 U873 ( .A1(n1152), .A2(n1188), .ZN(n1189) );
AND2_X1 U874 ( .A1(n1185), .A2(n1041), .ZN(n1152) );
AND4_X1 U875 ( .A1(n1184), .A2(n1032), .A3(n1037), .A4(n1178), .ZN(n1185) );
XNOR2_X1 U876 ( .A(n1190), .B(KEYINPUT53), .ZN(n1037) );
INV_X1 U877 ( .A(n1030), .ZN(n1184) );
NAND2_X1 U878 ( .A1(n1191), .A2(n1192), .ZN(n1030) );
XOR2_X1 U879 ( .A(n1193), .B(n1194), .Z(G30) );
NAND2_X1 U880 ( .A1(KEYINPUT38), .A2(n1151), .ZN(n1194) );
AND3_X1 U881 ( .A1(n1042), .A2(n1195), .A3(n1174), .ZN(n1151) );
AND3_X1 U882 ( .A1(n1178), .A2(n1196), .A3(n1197), .ZN(n1174) );
XNOR2_X1 U883 ( .A(G101), .B(n1170), .ZN(G3) );
NAND3_X1 U884 ( .A1(n1168), .A2(n1015), .A3(n1032), .ZN(n1170) );
XOR2_X1 U885 ( .A(G125), .B(n1198), .Z(G27) );
NOR3_X1 U886 ( .A1(n1160), .A2(n1199), .A3(n1019), .ZN(n1198) );
INV_X1 U887 ( .A(n1046), .ZN(n1019) );
NAND4_X1 U888 ( .A1(n1045), .A2(n1041), .A3(n1178), .A4(n1196), .ZN(n1160) );
NAND2_X1 U889 ( .A1(n1010), .A2(n1200), .ZN(n1178) );
NAND4_X1 U890 ( .A1(G902), .A2(G953), .A3(n1201), .A4(n1069), .ZN(n1200) );
INV_X1 U891 ( .A(G900), .ZN(n1069) );
XOR2_X1 U892 ( .A(n1202), .B(n1169), .Z(G24) );
NAND4_X1 U893 ( .A1(n1172), .A2(n1167), .A3(n1177), .A4(n1050), .ZN(n1169) );
INV_X1 U894 ( .A(n1023), .ZN(n1167) );
NAND2_X1 U895 ( .A1(n1045), .A2(n1203), .ZN(n1023) );
XOR2_X1 U896 ( .A(n1204), .B(n1166), .Z(G21) );
NAND4_X1 U897 ( .A1(n1197), .A2(n1172), .A3(n1015), .A4(n1196), .ZN(n1166) );
XOR2_X1 U898 ( .A(n1045), .B(KEYINPUT39), .Z(n1197) );
XOR2_X1 U899 ( .A(n1205), .B(n1165), .Z(G18) );
NAND3_X1 U900 ( .A1(n1172), .A2(n1042), .A3(n1032), .ZN(n1165) );
NAND2_X1 U901 ( .A1(n1206), .A2(n1207), .ZN(G15) );
NAND4_X1 U902 ( .A1(n1208), .A2(n1041), .A3(n1209), .A4(n1210), .ZN(n1207) );
XOR2_X1 U903 ( .A(n1211), .B(KEYINPUT19), .Z(n1206) );
NAND2_X1 U904 ( .A1(G113), .A2(n1212), .ZN(n1211) );
NAND3_X1 U905 ( .A1(n1041), .A2(n1209), .A3(n1208), .ZN(n1212) );
XNOR2_X1 U906 ( .A(n1032), .B(KEYINPUT48), .ZN(n1208) );
AND2_X1 U907 ( .A1(n1203), .A2(n1034), .ZN(n1032) );
INV_X1 U908 ( .A(n1045), .ZN(n1034) );
XOR2_X1 U909 ( .A(KEYINPUT0), .B(n1033), .Z(n1203) );
INV_X1 U910 ( .A(n1196), .ZN(n1033) );
NAND2_X1 U911 ( .A1(n1213), .A2(n1214), .ZN(n1209) );
NAND4_X1 U912 ( .A1(n1199), .A2(n1215), .A3(n1046), .A4(n1216), .ZN(n1214) );
INV_X1 U913 ( .A(KEYINPUT15), .ZN(n1216) );
NAND2_X1 U914 ( .A1(KEYINPUT15), .A2(n1172), .ZN(n1213) );
AND3_X1 U915 ( .A1(n1025), .A2(n1215), .A3(n1046), .ZN(n1172) );
NOR2_X1 U916 ( .A1(n1039), .A2(n1217), .ZN(n1046) );
INV_X1 U917 ( .A(n1199), .ZN(n1025) );
AND2_X1 U918 ( .A1(n1218), .A2(n1050), .ZN(n1041) );
XOR2_X1 U919 ( .A(KEYINPUT16), .B(n1219), .Z(n1218) );
XOR2_X1 U920 ( .A(n1164), .B(n1220), .Z(G12) );
NAND2_X1 U921 ( .A1(KEYINPUT9), .A2(n1221), .ZN(n1220) );
XOR2_X1 U922 ( .A(KEYINPUT62), .B(G110), .Z(n1221) );
NAND4_X1 U923 ( .A1(n1045), .A2(n1168), .A3(n1015), .A4(n1196), .ZN(n1164) );
NAND3_X1 U924 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1196) );
NAND2_X1 U925 ( .A1(G902), .A2(G217), .ZN(n1224) );
NAND3_X1 U926 ( .A1(n1097), .A2(n1148), .A3(n1225), .ZN(n1223) );
OR2_X1 U927 ( .A1(n1225), .A2(n1097), .ZN(n1222) );
AND3_X1 U928 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1097) );
NAND2_X1 U929 ( .A1(KEYINPUT10), .A2(n1229), .ZN(n1228) );
NAND3_X1 U930 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1227) );
INV_X1 U931 ( .A(KEYINPUT10), .ZN(n1231) );
OR2_X1 U932 ( .A1(n1232), .A2(n1230), .ZN(n1226) );
NOR2_X1 U933 ( .A1(KEYINPUT28), .A2(n1229), .ZN(n1230) );
XOR2_X1 U934 ( .A(n1233), .B(G137), .Z(n1229) );
NAND3_X1 U935 ( .A1(n1234), .A2(n1043), .A3(G221), .ZN(n1233) );
XNOR2_X1 U936 ( .A(KEYINPUT7), .B(n1235), .ZN(n1234) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1232) );
XNOR2_X1 U938 ( .A(n1238), .B(n1239), .ZN(n1237) );
NOR2_X1 U939 ( .A1(KEYINPUT51), .A2(n1240), .ZN(n1239) );
XOR2_X1 U940 ( .A(n1075), .B(KEYINPUT47), .Z(n1240) );
INV_X1 U941 ( .A(n1241), .ZN(n1075) );
NAND2_X1 U942 ( .A1(n1242), .A2(KEYINPUT43), .ZN(n1238) );
XOR2_X1 U943 ( .A(n1193), .B(G119), .Z(n1242) );
XNOR2_X1 U944 ( .A(G110), .B(n1243), .ZN(n1236) );
XOR2_X1 U945 ( .A(KEYINPUT49), .B(G146), .Z(n1243) );
NAND2_X1 U946 ( .A1(G217), .A2(n1244), .ZN(n1225) );
INV_X1 U947 ( .A(G234), .ZN(n1244) );
NAND2_X1 U948 ( .A1(n1245), .A2(n1246), .ZN(n1015) );
OR3_X1 U949 ( .A1(n1050), .A2(n1177), .A3(KEYINPUT16), .ZN(n1246) );
NAND2_X1 U950 ( .A1(KEYINPUT16), .A2(n1042), .ZN(n1245) );
NOR2_X1 U951 ( .A1(n1050), .A2(n1219), .ZN(n1042) );
INV_X1 U952 ( .A(n1177), .ZN(n1219) );
XOR2_X1 U953 ( .A(n1060), .B(G478), .Z(n1177) );
NOR2_X1 U954 ( .A1(n1102), .A2(G902), .ZN(n1060) );
XNOR2_X1 U955 ( .A(n1247), .B(n1248), .ZN(n1102) );
XOR2_X1 U956 ( .A(G128), .B(n1249), .Z(n1248) );
XOR2_X1 U957 ( .A(G143), .B(G134), .Z(n1249) );
XOR2_X1 U958 ( .A(n1250), .B(n1251), .Z(n1247) );
XOR2_X1 U959 ( .A(n1252), .B(G116), .Z(n1250) );
NAND3_X1 U960 ( .A1(n1235), .A2(n1253), .A3(G217), .ZN(n1252) );
XOR2_X1 U961 ( .A(KEYINPUT59), .B(G953), .Z(n1253) );
XNOR2_X1 U962 ( .A(G234), .B(KEYINPUT58), .ZN(n1235) );
XNOR2_X1 U963 ( .A(n1254), .B(G475), .ZN(n1050) );
NAND2_X1 U964 ( .A1(n1115), .A2(n1148), .ZN(n1254) );
XOR2_X1 U965 ( .A(n1255), .B(n1256), .Z(n1115) );
XOR2_X1 U966 ( .A(KEYINPUT49), .B(G131), .Z(n1256) );
XOR2_X1 U967 ( .A(n1257), .B(G122), .Z(n1255) );
XOR2_X1 U968 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U969 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U970 ( .A(KEYINPUT36), .B(G113), .Z(n1261) );
XOR2_X1 U971 ( .A(KEYINPUT61), .B(KEYINPUT55), .Z(n1260) );
XOR2_X1 U972 ( .A(n1262), .B(n1263), .Z(n1258) );
XOR2_X1 U973 ( .A(n1264), .B(n1241), .Z(n1263) );
XOR2_X1 U974 ( .A(G125), .B(G140), .Z(n1241) );
XOR2_X1 U975 ( .A(n1265), .B(G104), .Z(n1262) );
NAND2_X1 U976 ( .A1(G214), .A2(n1266), .ZN(n1265) );
AND2_X1 U977 ( .A1(n1195), .A2(n1215), .ZN(n1168) );
NAND2_X1 U978 ( .A1(n1267), .A2(n1010), .ZN(n1215) );
NAND3_X1 U979 ( .A1(n1201), .A2(n1043), .A3(n1268), .ZN(n1010) );
XOR2_X1 U980 ( .A(n1109), .B(KEYINPUT52), .Z(n1268) );
INV_X1 U981 ( .A(G952), .ZN(n1109) );
NAND4_X1 U982 ( .A1(G902), .A2(n1269), .A3(n1201), .A4(n1088), .ZN(n1267) );
INV_X1 U983 ( .A(G898), .ZN(n1088) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1201) );
XOR2_X1 U985 ( .A(KEYINPUT26), .B(G953), .Z(n1269) );
NOR2_X1 U986 ( .A1(n1199), .A2(n1190), .ZN(n1195) );
NAND2_X1 U987 ( .A1(n1270), .A2(n1039), .ZN(n1190) );
XNOR2_X1 U988 ( .A(n1271), .B(G469), .ZN(n1039) );
NAND2_X1 U989 ( .A1(n1272), .A2(n1148), .ZN(n1271) );
XOR2_X1 U990 ( .A(n1130), .B(n1273), .Z(n1272) );
XOR2_X1 U991 ( .A(G110), .B(n1274), .Z(n1273) );
NOR2_X1 U992 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U993 ( .A(KEYINPUT37), .B(n1277), .Z(n1276) );
NOR2_X1 U994 ( .A1(n1078), .A2(n1278), .ZN(n1277) );
AND2_X1 U995 ( .A1(n1278), .A2(n1078), .ZN(n1275) );
NAND2_X1 U996 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U997 ( .A1(n1077), .A2(n1281), .ZN(n1280) );
NAND2_X1 U998 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
OR2_X1 U999 ( .A1(n1132), .A2(KEYINPUT25), .ZN(n1283) );
NAND2_X1 U1000 ( .A1(n1132), .A2(n1284), .ZN(n1279) );
NAND2_X1 U1001 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U1002 ( .A1(n1287), .A2(n1282), .ZN(n1286) );
INV_X1 U1003 ( .A(KEYINPUT50), .ZN(n1282) );
INV_X1 U1004 ( .A(n1077), .ZN(n1287) );
XOR2_X1 U1005 ( .A(n1288), .B(KEYINPUT29), .Z(n1077) );
INV_X1 U1006 ( .A(KEYINPUT25), .ZN(n1285) );
XOR2_X1 U1007 ( .A(n1289), .B(n1290), .Z(n1132) );
XOR2_X1 U1008 ( .A(G140), .B(n1291), .Z(n1130) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1068), .ZN(n1291) );
INV_X1 U1010 ( .A(G227), .ZN(n1068) );
XOR2_X1 U1011 ( .A(KEYINPUT57), .B(n1217), .Z(n1270) );
INV_X1 U1012 ( .A(n1038), .ZN(n1217) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1292), .ZN(n1038) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1148), .ZN(n1292) );
NAND2_X1 U1015 ( .A1(n1192), .A2(n1027), .ZN(n1199) );
INV_X1 U1016 ( .A(n1191), .ZN(n1027) );
XOR2_X1 U1017 ( .A(n1051), .B(n1053), .Z(n1191) );
AND2_X1 U1018 ( .A1(G210), .A2(n1293), .ZN(n1053) );
NAND2_X1 U1019 ( .A1(n1294), .A2(n1148), .ZN(n1051) );
XOR2_X1 U1020 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1021 ( .A(n1086), .B(n1145), .Z(n1296) );
XOR2_X1 U1022 ( .A(n1288), .B(G125), .Z(n1145) );
XOR2_X1 U1023 ( .A(n1297), .B(n1298), .Z(n1086) );
XOR2_X1 U1024 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1025 ( .A(KEYINPUT34), .B(G110), .Z(n1300) );
NOR2_X1 U1026 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
INV_X1 U1027 ( .A(n1303), .ZN(n1301) );
XNOR2_X1 U1028 ( .A(n1251), .B(n1289), .ZN(n1297) );
XOR2_X1 U1029 ( .A(G101), .B(G104), .Z(n1289) );
XNOR2_X1 U1030 ( .A(n1202), .B(n1290), .ZN(n1251) );
XOR2_X1 U1031 ( .A(G107), .B(KEYINPUT5), .Z(n1290) );
INV_X1 U1032 ( .A(G122), .ZN(n1202) );
XNOR2_X1 U1033 ( .A(KEYINPUT11), .B(n1147), .ZN(n1295) );
NAND2_X1 U1034 ( .A1(G224), .A2(n1043), .ZN(n1147) );
INV_X1 U1035 ( .A(G953), .ZN(n1043) );
XNOR2_X1 U1036 ( .A(n1028), .B(KEYINPUT63), .ZN(n1192) );
AND2_X1 U1037 ( .A1(G214), .A2(n1293), .ZN(n1028) );
OR2_X1 U1038 ( .A1(G902), .A2(G237), .ZN(n1293) );
XOR2_X1 U1039 ( .A(n1304), .B(G472), .Z(n1045) );
NAND2_X1 U1040 ( .A1(n1305), .A2(n1148), .ZN(n1304) );
INV_X1 U1041 ( .A(G902), .ZN(n1148) );
XNOR2_X1 U1042 ( .A(n1119), .B(n1306), .ZN(n1305) );
NOR2_X1 U1043 ( .A1(KEYINPUT40), .A2(n1078), .ZN(n1306) );
XNOR2_X1 U1044 ( .A(n1188), .B(n1307), .ZN(n1078) );
XOR2_X1 U1045 ( .A(G137), .B(G134), .Z(n1307) );
INV_X1 U1046 ( .A(G131), .ZN(n1188) );
XNOR2_X1 U1047 ( .A(n1308), .B(n1309), .ZN(n1119) );
XOR2_X1 U1048 ( .A(n1310), .B(n1311), .Z(n1309) );
INV_X1 U1049 ( .A(n1288), .ZN(n1311) );
XOR2_X1 U1050 ( .A(n1193), .B(n1264), .Z(n1288) );
XNOR2_X1 U1051 ( .A(G143), .B(n1173), .ZN(n1264) );
INV_X1 U1052 ( .A(G146), .ZN(n1173) );
INV_X1 U1053 ( .A(G128), .ZN(n1193) );
AND2_X1 U1054 ( .A1(n1266), .A2(G210), .ZN(n1310) );
NOR2_X1 U1055 ( .A1(G953), .A2(G237), .ZN(n1266) );
XOR2_X1 U1056 ( .A(n1312), .B(G101), .Z(n1308) );
NAND3_X1 U1057 ( .A1(n1313), .A2(n1314), .A3(n1303), .ZN(n1312) );
NAND3_X1 U1058 ( .A1(G113), .A2(n1204), .A3(G116), .ZN(n1303) );
NAND2_X1 U1059 ( .A1(n1302), .A2(n1315), .ZN(n1314) );
INV_X1 U1060 ( .A(KEYINPUT33), .ZN(n1315) );
NAND2_X1 U1061 ( .A1(n1316), .A2(n1317), .ZN(n1302) );
NAND3_X1 U1062 ( .A1(n1210), .A2(n1205), .A3(n1204), .ZN(n1317) );
INV_X1 U1063 ( .A(G116), .ZN(n1205) );
INV_X1 U1064 ( .A(G113), .ZN(n1210) );
NAND2_X1 U1065 ( .A1(n1318), .A2(G119), .ZN(n1316) );
XOR2_X1 U1066 ( .A(G116), .B(G113), .Z(n1318) );
NAND2_X1 U1067 ( .A1(n1319), .A2(KEYINPUT33), .ZN(n1313) );
XOR2_X1 U1068 ( .A(G113), .B(n1320), .Z(n1319) );
NOR2_X1 U1069 ( .A1(G116), .A2(n1204), .ZN(n1320) );
INV_X1 U1070 ( .A(G119), .ZN(n1204) );
endmodule


