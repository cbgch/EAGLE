//Key = 0011101101010100110100001011101101111000101000010011010101111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271;

XOR2_X1 U695 ( .A(G107), .B(n959), .Z(G9) );
NOR2_X1 U696 ( .A1(n960), .A2(n961), .ZN(G75) );
NOR4_X1 U697 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n961) );
NOR2_X1 U698 ( .A1(n966), .A2(n967), .ZN(n964) );
NOR2_X1 U699 ( .A1(n968), .A2(n969), .ZN(n966) );
NAND3_X1 U700 ( .A1(n970), .A2(n971), .A3(n972), .ZN(n962) );
NAND3_X1 U701 ( .A1(n973), .A2(n974), .A3(n975), .ZN(n972) );
NAND2_X1 U702 ( .A1(n976), .A2(n977), .ZN(n973) );
NAND3_X1 U703 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NAND2_X1 U704 ( .A1(n981), .A2(n982), .ZN(n979) );
NAND2_X1 U705 ( .A1(n983), .A2(n984), .ZN(n982) );
OR2_X1 U706 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND2_X1 U707 ( .A1(n987), .A2(n988), .ZN(n981) );
NAND2_X1 U708 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND2_X1 U709 ( .A1(n991), .A2(n992), .ZN(n990) );
XNOR2_X1 U710 ( .A(n993), .B(KEYINPUT15), .ZN(n989) );
NAND2_X1 U711 ( .A1(n994), .A2(n995), .ZN(n976) );
NAND2_X1 U712 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND2_X1 U713 ( .A1(n998), .A2(n967), .ZN(n997) );
INV_X1 U714 ( .A(KEYINPUT18), .ZN(n967) );
NAND3_X1 U715 ( .A1(n978), .A2(n999), .A3(n994), .ZN(n970) );
INV_X1 U716 ( .A(n969), .ZN(n994) );
NAND3_X1 U717 ( .A1(n983), .A2(n987), .A3(n980), .ZN(n969) );
INV_X1 U718 ( .A(n1000), .ZN(n980) );
NAND2_X1 U719 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND2_X1 U720 ( .A1(n1003), .A2(n975), .ZN(n1002) );
NOR3_X1 U721 ( .A1(n965), .A2(G952), .A3(n1004), .ZN(n960) );
INV_X1 U722 ( .A(n971), .ZN(n1004) );
NAND4_X1 U723 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n971) );
NOR3_X1 U724 ( .A1(n1009), .A2(n991), .A3(n1003), .ZN(n1008) );
NOR2_X1 U725 ( .A1(G469), .A2(n1010), .ZN(n1009) );
NOR3_X1 U726 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1007) );
NOR2_X1 U727 ( .A1(KEYINPUT59), .A2(n1014), .ZN(n1013) );
XNOR2_X1 U728 ( .A(n1015), .B(n1016), .ZN(n1014) );
NOR2_X1 U729 ( .A1(n1017), .A2(n1018), .ZN(n1012) );
INV_X1 U730 ( .A(KEYINPUT59), .ZN(n1018) );
NOR2_X1 U731 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
INV_X1 U732 ( .A(n1021), .ZN(n1020) );
XOR2_X1 U733 ( .A(KEYINPUT50), .B(n1022), .Z(n1011) );
NOR3_X1 U734 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
XOR2_X1 U735 ( .A(n1026), .B(n1027), .Z(n1024) );
NOR2_X1 U736 ( .A1(n1028), .A2(KEYINPUT0), .ZN(n1027) );
INV_X1 U737 ( .A(n1029), .ZN(n1028) );
XOR2_X1 U738 ( .A(G472), .B(n1030), .Z(n1023) );
NOR2_X1 U739 ( .A1(KEYINPUT1), .A2(n1031), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1006) );
INV_X1 U741 ( .A(KEYINPUT4), .ZN(n1033) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1010), .ZN(n1032) );
XNOR2_X1 U743 ( .A(KEYINPUT2), .B(G469), .ZN(n1034) );
NAND2_X1 U744 ( .A1(KEYINPUT4), .A2(n1035), .ZN(n1005) );
NAND2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
OR2_X1 U746 ( .A1(G469), .A2(KEYINPUT2), .ZN(n1037) );
NAND3_X1 U747 ( .A1(G469), .A2(n1010), .A3(KEYINPUT2), .ZN(n1036) );
XOR2_X1 U748 ( .A(n1038), .B(n1039), .Z(G72) );
XOR2_X1 U749 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U750 ( .A1(G953), .A2(n1042), .ZN(n1041) );
XOR2_X1 U751 ( .A(n1043), .B(KEYINPUT60), .Z(n1042) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1040) );
NAND2_X1 U754 ( .A1(G953), .A2(n1048), .ZN(n1047) );
XOR2_X1 U755 ( .A(n1049), .B(n1050), .Z(n1046) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U757 ( .A(KEYINPUT46), .B(KEYINPUT34), .ZN(n1051) );
XOR2_X1 U758 ( .A(n1053), .B(KEYINPUT56), .Z(n1049) );
NAND3_X1 U759 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U761 ( .A1(KEYINPUT16), .A2(n1059), .ZN(n1058) );
XNOR2_X1 U762 ( .A(KEYINPUT12), .B(n1060), .ZN(n1057) );
OR2_X1 U763 ( .A1(n1059), .A2(KEYINPUT55), .ZN(n1055) );
NAND4_X1 U764 ( .A1(n1059), .A2(n1061), .A3(KEYINPUT16), .A4(KEYINPUT55), .ZN(n1054) );
XOR2_X1 U765 ( .A(KEYINPUT12), .B(n1060), .Z(n1061) );
XOR2_X1 U766 ( .A(G131), .B(n1062), .Z(n1059) );
NAND2_X1 U767 ( .A1(G953), .A2(n1063), .ZN(n1038) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(G69) );
NAND2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1064) );
NAND2_X1 U772 ( .A1(n1070), .A2(n1067), .ZN(n1069) );
NAND2_X1 U773 ( .A1(G953), .A2(n1071), .ZN(n1067) );
INV_X1 U774 ( .A(n1072), .ZN(n1070) );
INV_X1 U775 ( .A(n1066), .ZN(n1068) );
XNOR2_X1 U776 ( .A(n1073), .B(n1074), .ZN(n1066) );
NOR3_X1 U777 ( .A1(n1072), .A2(n1075), .A3(n1076), .ZN(n1074) );
NOR2_X1 U778 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U779 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
AND2_X1 U780 ( .A1(n1078), .A2(n1081), .ZN(n1075) );
INV_X1 U781 ( .A(KEYINPUT44), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1082), .A2(n1083), .ZN(n1073) );
NAND2_X1 U783 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U784 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U785 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U786 ( .A1(n1029), .A2(n1090), .ZN(n1089) );
NAND2_X1 U787 ( .A1(KEYINPUT17), .A2(n1091), .ZN(n1088) );
NOR2_X1 U788 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND3_X1 U790 ( .A1(n1095), .A2(G478), .A3(KEYINPUT57), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1086), .A2(n1096), .ZN(G60) );
NOR2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U793 ( .A(KEYINPUT32), .B(n1099), .Z(n1098) );
NOR2_X1 U794 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
AND2_X1 U795 ( .A1(n1101), .A2(n1100), .ZN(n1097) );
NAND2_X1 U796 ( .A1(n1095), .A2(G475), .ZN(n1101) );
XOR2_X1 U797 ( .A(n1102), .B(n1103), .Z(G6) );
NOR2_X1 U798 ( .A1(KEYINPUT48), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U799 ( .A(KEYINPUT29), .B(n1105), .ZN(n1104) );
NAND2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1102) );
XNOR2_X1 U801 ( .A(n1108), .B(KEYINPUT61), .ZN(n1106) );
NOR2_X1 U802 ( .A1(n1086), .A2(n1109), .ZN(G57) );
XNOR2_X1 U803 ( .A(n1110), .B(n1111), .ZN(n1109) );
XOR2_X1 U804 ( .A(n1112), .B(n1113), .Z(n1111) );
AND2_X1 U805 ( .A1(G472), .A2(n1095), .ZN(n1113) );
NAND2_X1 U806 ( .A1(KEYINPUT28), .A2(n1114), .ZN(n1112) );
NOR2_X1 U807 ( .A1(n1086), .A2(n1115), .ZN(G54) );
XOR2_X1 U808 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U809 ( .A(n1118), .B(n1060), .Z(n1117) );
XOR2_X1 U810 ( .A(n1119), .B(n1120), .Z(n1116) );
XOR2_X1 U811 ( .A(n1121), .B(n1122), .Z(n1120) );
AND2_X1 U812 ( .A1(G469), .A2(n1095), .ZN(n1122) );
INV_X1 U813 ( .A(n1090), .ZN(n1095) );
NAND2_X1 U814 ( .A1(KEYINPUT24), .A2(n1123), .ZN(n1119) );
NOR2_X1 U815 ( .A1(n1082), .A2(G952), .ZN(n1086) );
NOR2_X1 U816 ( .A1(n1124), .A2(n1125), .ZN(G51) );
XOR2_X1 U817 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U818 ( .A(n1081), .B(n1128), .Z(n1127) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U820 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U821 ( .A(KEYINPUT8), .B(n1133), .ZN(n1131) );
NOR2_X1 U822 ( .A1(n1134), .A2(n1135), .ZN(n1129) );
XNOR2_X1 U823 ( .A(n1136), .B(KEYINPUT14), .ZN(n1135) );
XOR2_X1 U824 ( .A(KEYINPUT52), .B(n1137), .Z(n1126) );
NOR2_X1 U825 ( .A1(n1138), .A2(n1090), .ZN(n1137) );
NAND2_X1 U826 ( .A1(G902), .A2(n963), .ZN(n1090) );
NAND4_X1 U827 ( .A1(n1139), .A2(n1084), .A3(n1044), .A4(n1140), .ZN(n963) );
XOR2_X1 U828 ( .A(KEYINPUT62), .B(n1045), .Z(n1140) );
AND4_X1 U829 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1045) );
AND4_X1 U830 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1044) );
NAND2_X1 U831 ( .A1(n1149), .A2(n1150), .ZN(n1145) );
XNOR2_X1 U832 ( .A(KEYINPUT5), .B(n996), .ZN(n1150) );
AND4_X1 U833 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1084) );
NOR4_X1 U834 ( .A1(n959), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1154) );
INV_X1 U835 ( .A(n1158), .ZN(n1155) );
AND3_X1 U836 ( .A1(n1159), .A2(n987), .A3(n1160), .ZN(n959) );
NAND2_X1 U837 ( .A1(n1108), .A2(n1107), .ZN(n1153) );
AND4_X1 U838 ( .A1(n998), .A2(n1161), .A3(n987), .A4(n1162), .ZN(n1108) );
XOR2_X1 U839 ( .A(n1085), .B(KEYINPUT41), .Z(n1139) );
NOR2_X1 U840 ( .A1(n1082), .A2(n1163), .ZN(n1124) );
XOR2_X1 U841 ( .A(KEYINPUT25), .B(G952), .Z(n1163) );
XNOR2_X1 U842 ( .A(G146), .B(n1141), .ZN(G48) );
NAND2_X1 U843 ( .A1(n1164), .A2(n998), .ZN(n1141) );
XNOR2_X1 U844 ( .A(G143), .B(n1142), .ZN(G45) );
NAND3_X1 U845 ( .A1(n1165), .A2(n986), .A3(n1166), .ZN(n1142) );
NOR3_X1 U846 ( .A1(n1001), .A2(n1167), .A3(n1168), .ZN(n1166) );
INV_X1 U847 ( .A(n1161), .ZN(n1001) );
XNOR2_X1 U848 ( .A(G140), .B(n1143), .ZN(G42) );
NAND3_X1 U849 ( .A1(n985), .A2(n998), .A3(n1169), .ZN(n1143) );
XNOR2_X1 U850 ( .A(G137), .B(n1144), .ZN(G39) );
NAND2_X1 U851 ( .A1(n1169), .A2(n1170), .ZN(n1144) );
XNOR2_X1 U852 ( .A(G134), .B(n1171), .ZN(G36) );
NAND2_X1 U853 ( .A1(n1149), .A2(n1160), .ZN(n1171) );
XNOR2_X1 U854 ( .A(G131), .B(n1146), .ZN(G33) );
NAND2_X1 U855 ( .A1(n1149), .A2(n998), .ZN(n1146) );
AND2_X1 U856 ( .A1(n1169), .A2(n986), .ZN(n1149) );
AND3_X1 U857 ( .A1(n1161), .A2(n1172), .A3(n983), .ZN(n1169) );
NOR2_X1 U858 ( .A1(n1173), .A2(n991), .ZN(n983) );
XNOR2_X1 U859 ( .A(G128), .B(n1147), .ZN(G30) );
NAND2_X1 U860 ( .A1(n1164), .A2(n1160), .ZN(n1147) );
AND4_X1 U861 ( .A1(n1165), .A2(n1161), .A3(n1174), .A4(n1175), .ZN(n1164) );
XNOR2_X1 U862 ( .A(G101), .B(n1151), .ZN(G3) );
NAND3_X1 U863 ( .A1(n1159), .A2(n986), .A3(n978), .ZN(n1151) );
XNOR2_X1 U864 ( .A(G125), .B(n1148), .ZN(G27) );
NAND3_X1 U865 ( .A1(n1165), .A2(n1176), .A3(n985), .ZN(n1148) );
AND2_X1 U866 ( .A1(n993), .A2(n1172), .ZN(n1165) );
NAND2_X1 U867 ( .A1(n1000), .A2(n1177), .ZN(n1172) );
NAND4_X1 U868 ( .A1(G902), .A2(G953), .A3(n1178), .A4(n1048), .ZN(n1177) );
INV_X1 U869 ( .A(G900), .ZN(n1048) );
XNOR2_X1 U870 ( .A(G122), .B(n1152), .ZN(G24) );
NAND4_X1 U871 ( .A1(n1179), .A2(n1180), .A3(n987), .A4(n1181), .ZN(n1152) );
NAND2_X1 U872 ( .A1(n1182), .A2(n1183), .ZN(n987) );
OR3_X1 U873 ( .A1(n1174), .A2(n1175), .A3(KEYINPUT43), .ZN(n1183) );
NAND2_X1 U874 ( .A1(KEYINPUT43), .A2(n986), .ZN(n1182) );
XOR2_X1 U875 ( .A(G119), .B(n1157), .Z(G21) );
AND2_X1 U876 ( .A1(n1170), .A2(n1179), .ZN(n1157) );
AND3_X1 U877 ( .A1(n1174), .A2(n1175), .A3(n978), .ZN(n1170) );
XOR2_X1 U878 ( .A(G116), .B(n1156), .Z(G18) );
AND3_X1 U879 ( .A1(n1160), .A2(n986), .A3(n1179), .ZN(n1156) );
AND4_X1 U880 ( .A1(n975), .A2(n993), .A3(n1162), .A4(n974), .ZN(n1179) );
XOR2_X1 U881 ( .A(n1107), .B(KEYINPUT22), .Z(n993) );
INV_X1 U882 ( .A(n996), .ZN(n1160) );
NAND2_X1 U883 ( .A1(n1184), .A2(n1181), .ZN(n996) );
XNOR2_X1 U884 ( .A(G113), .B(n1158), .ZN(G15) );
NAND4_X1 U885 ( .A1(n1176), .A2(n986), .A3(n1107), .A4(n1162), .ZN(n1158) );
NOR2_X1 U886 ( .A1(n1174), .A2(n1185), .ZN(n986) );
INV_X1 U887 ( .A(n1175), .ZN(n1185) );
INV_X1 U888 ( .A(n968), .ZN(n1176) );
NAND3_X1 U889 ( .A1(n975), .A2(n974), .A3(n998), .ZN(n968) );
NOR2_X1 U890 ( .A1(n1181), .A2(n1168), .ZN(n998) );
INV_X1 U891 ( .A(n1180), .ZN(n1168) );
XNOR2_X1 U892 ( .A(n1184), .B(KEYINPUT45), .ZN(n1180) );
XNOR2_X1 U893 ( .A(G110), .B(n1085), .ZN(G12) );
NAND3_X1 U894 ( .A1(n978), .A2(n1159), .A3(n985), .ZN(n1085) );
AND2_X1 U895 ( .A1(n1186), .A2(n1174), .ZN(n985) );
XOR2_X1 U896 ( .A(n1026), .B(n1029), .Z(n1174) );
NAND2_X1 U897 ( .A1(G217), .A2(n1187), .ZN(n1029) );
NAND2_X1 U898 ( .A1(n1091), .A2(n1188), .ZN(n1026) );
XNOR2_X1 U899 ( .A(n1189), .B(n1190), .ZN(n1091) );
XNOR2_X1 U900 ( .A(n1191), .B(n1192), .ZN(n1190) );
NOR2_X1 U901 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U902 ( .A(n1195), .B(KEYINPUT26), .Z(n1194) );
NAND2_X1 U903 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR2_X1 U904 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n1198), .ZN(n1197) );
XNOR2_X1 U906 ( .A(G128), .B(n1199), .ZN(n1196) );
INV_X1 U907 ( .A(G146), .ZN(n1191) );
XNOR2_X1 U908 ( .A(n1200), .B(n1201), .ZN(n1189) );
NAND2_X1 U909 ( .A1(KEYINPUT30), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U910 ( .A(G137), .B(n1203), .ZN(n1202) );
NAND2_X1 U911 ( .A1(G221), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U912 ( .A(KEYINPUT43), .B(n1175), .ZN(n1186) );
XNOR2_X1 U913 ( .A(n1031), .B(G472), .ZN(n1175) );
NAND2_X1 U914 ( .A1(n1205), .A2(n1188), .ZN(n1031) );
XOR2_X1 U915 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U916 ( .A(KEYINPUT23), .B(KEYINPUT19), .Z(n1207) );
XNOR2_X1 U917 ( .A(n1114), .B(n1208), .ZN(n1206) );
INV_X1 U918 ( .A(n1110), .ZN(n1208) );
XNOR2_X1 U919 ( .A(n1209), .B(n1210), .ZN(n1110) );
XNOR2_X1 U920 ( .A(G101), .B(n1211), .ZN(n1210) );
NAND2_X1 U921 ( .A1(G210), .A2(n1212), .ZN(n1211) );
XOR2_X1 U922 ( .A(n1213), .B(n1214), .Z(n1209) );
NAND2_X1 U923 ( .A1(KEYINPUT35), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U924 ( .A(KEYINPUT3), .B(n1216), .ZN(n1215) );
XOR2_X1 U925 ( .A(n1217), .B(n1218), .Z(n1114) );
AND3_X1 U926 ( .A1(n1161), .A2(n1162), .A3(n1107), .ZN(n1159) );
NOR2_X1 U927 ( .A1(n991), .A2(n992), .ZN(n1107) );
INV_X1 U928 ( .A(n1173), .ZN(n992) );
NAND2_X1 U929 ( .A1(n1219), .A2(n1021), .ZN(n1173) );
NAND2_X1 U930 ( .A1(n1016), .A2(n1015), .ZN(n1021) );
XNOR2_X1 U931 ( .A(n1019), .B(KEYINPUT54), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1015), .A2(n1016), .ZN(n1019) );
INV_X1 U933 ( .A(n1138), .ZN(n1016) );
NAND2_X1 U934 ( .A1(G210), .A2(n1220), .ZN(n1138) );
NAND2_X1 U935 ( .A1(n1221), .A2(n1188), .ZN(n1015) );
XNOR2_X1 U936 ( .A(n1081), .B(n1222), .ZN(n1221) );
XNOR2_X1 U937 ( .A(n1223), .B(KEYINPUT38), .ZN(n1222) );
NAND2_X1 U938 ( .A1(KEYINPUT53), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U939 ( .A(n1132), .B(n1225), .ZN(n1224) );
XNOR2_X1 U940 ( .A(KEYINPUT58), .B(n1133), .ZN(n1225) );
INV_X1 U941 ( .A(n1136), .ZN(n1133) );
NOR2_X1 U942 ( .A1(n1071), .A2(G953), .ZN(n1136) );
INV_X1 U943 ( .A(G224), .ZN(n1071) );
INV_X1 U944 ( .A(n1134), .ZN(n1132) );
XOR2_X1 U945 ( .A(G125), .B(n1218), .Z(n1134) );
XNOR2_X1 U946 ( .A(n1226), .B(KEYINPUT39), .ZN(n1218) );
XNOR2_X1 U947 ( .A(n1079), .B(n1080), .ZN(n1081) );
XNOR2_X1 U948 ( .A(n1198), .B(G122), .ZN(n1080) );
INV_X1 U949 ( .A(G110), .ZN(n1198) );
XOR2_X1 U950 ( .A(n1227), .B(n1228), .Z(n1079) );
XNOR2_X1 U951 ( .A(n1229), .B(n1216), .ZN(n1227) );
NAND2_X1 U952 ( .A1(KEYINPUT7), .A2(n1214), .ZN(n1229) );
XOR2_X1 U953 ( .A(G116), .B(n1199), .Z(n1214) );
XOR2_X1 U954 ( .A(G119), .B(KEYINPUT33), .Z(n1199) );
AND2_X1 U955 ( .A1(G214), .A2(n1220), .ZN(n991) );
NAND2_X1 U956 ( .A1(n1230), .A2(n1188), .ZN(n1220) );
INV_X1 U957 ( .A(G237), .ZN(n1230) );
NAND2_X1 U958 ( .A1(n1000), .A2(n1231), .ZN(n1162) );
NAND3_X1 U959 ( .A1(n1072), .A2(n1178), .A3(G902), .ZN(n1231) );
NOR2_X1 U960 ( .A1(G898), .A2(n1082), .ZN(n1072) );
NAND3_X1 U961 ( .A1(n1232), .A2(n1178), .A3(G952), .ZN(n1000) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1178) );
INV_X1 U963 ( .A(n965), .ZN(n1232) );
XOR2_X1 U964 ( .A(G953), .B(KEYINPUT49), .Z(n965) );
NOR2_X1 U965 ( .A1(n975), .A2(n1003), .ZN(n1161) );
INV_X1 U966 ( .A(n974), .ZN(n1003) );
NAND2_X1 U967 ( .A1(G221), .A2(n1187), .ZN(n974) );
NAND2_X1 U968 ( .A1(G234), .A2(n1188), .ZN(n1187) );
XOR2_X1 U969 ( .A(n1010), .B(G469), .Z(n975) );
NAND2_X1 U970 ( .A1(n1233), .A2(n1188), .ZN(n1010) );
XOR2_X1 U971 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U972 ( .A(n1236), .B(n1121), .ZN(n1235) );
NAND2_X1 U973 ( .A1(G227), .A2(n1082), .ZN(n1121) );
NAND2_X1 U974 ( .A1(n1237), .A2(KEYINPUT42), .ZN(n1236) );
XOR2_X1 U975 ( .A(n1238), .B(n1118), .Z(n1237) );
XNOR2_X1 U976 ( .A(n1217), .B(n1228), .ZN(n1118) );
XNOR2_X1 U977 ( .A(n1239), .B(n1240), .ZN(n1228) );
XNOR2_X1 U978 ( .A(KEYINPUT6), .B(n1105), .ZN(n1240) );
XNOR2_X1 U979 ( .A(G101), .B(n1241), .ZN(n1239) );
NAND2_X1 U980 ( .A1(n1242), .A2(n1243), .ZN(n1217) );
NAND2_X1 U981 ( .A1(n1062), .A2(n1244), .ZN(n1243) );
XOR2_X1 U982 ( .A(n1245), .B(KEYINPUT63), .Z(n1242) );
OR2_X1 U983 ( .A1(n1244), .A2(n1062), .ZN(n1245) );
XNOR2_X1 U984 ( .A(G134), .B(G137), .ZN(n1062) );
XOR2_X1 U985 ( .A(G131), .B(KEYINPUT47), .Z(n1244) );
NAND2_X1 U986 ( .A1(KEYINPUT27), .A2(n1060), .ZN(n1238) );
XNOR2_X1 U987 ( .A(n1226), .B(KEYINPUT20), .ZN(n1060) );
XOR2_X1 U988 ( .A(n1246), .B(n1247), .Z(n1226) );
XNOR2_X1 U989 ( .A(G146), .B(KEYINPUT37), .ZN(n1246) );
NAND2_X1 U990 ( .A1(KEYINPUT31), .A2(n1123), .ZN(n1234) );
XOR2_X1 U991 ( .A(G140), .B(G110), .Z(n1123) );
INV_X1 U992 ( .A(n1025), .ZN(n978) );
NAND2_X1 U993 ( .A1(n1167), .A2(n1184), .ZN(n1025) );
XOR2_X1 U994 ( .A(n1248), .B(G475), .Z(n1184) );
NAND2_X1 U995 ( .A1(n1100), .A2(n1188), .ZN(n1248) );
XNOR2_X1 U996 ( .A(n1249), .B(n1250), .ZN(n1100) );
XNOR2_X1 U997 ( .A(G146), .B(n1251), .ZN(n1250) );
NAND2_X1 U998 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND4_X1 U999 ( .A1(KEYINPUT40), .A2(KEYINPUT11), .A3(n1254), .A4(n1105), .ZN(n1253) );
NAND2_X1 U1000 ( .A1(n1255), .A2(n1256), .ZN(n1252) );
NAND2_X1 U1001 ( .A1(n1257), .A2(n1105), .ZN(n1256) );
INV_X1 U1002 ( .A(G104), .ZN(n1105) );
OR2_X1 U1003 ( .A1(n1254), .A2(KEYINPUT11), .ZN(n1257) );
NAND2_X1 U1004 ( .A1(KEYINPUT40), .A2(n1254), .ZN(n1255) );
XOR2_X1 U1005 ( .A(n1258), .B(G122), .Z(n1254) );
NAND2_X1 U1006 ( .A1(KEYINPUT51), .A2(n1216), .ZN(n1258) );
INV_X1 U1007 ( .A(G113), .ZN(n1216) );
XNOR2_X1 U1008 ( .A(n1259), .B(n1260), .ZN(n1249) );
NAND2_X1 U1009 ( .A1(n1261), .A2(KEYINPUT9), .ZN(n1260) );
XOR2_X1 U1010 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U1011 ( .A(G131), .B(n1264), .ZN(n1263) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1212), .ZN(n1264) );
NOR2_X1 U1013 ( .A1(G953), .A2(G237), .ZN(n1212) );
NAND2_X1 U1014 ( .A1(KEYINPUT13), .A2(n1265), .ZN(n1262) );
NAND2_X1 U1015 ( .A1(KEYINPUT36), .A2(n1201), .ZN(n1259) );
INV_X1 U1016 ( .A(n1052), .ZN(n1201) );
XOR2_X1 U1017 ( .A(G125), .B(G140), .Z(n1052) );
INV_X1 U1018 ( .A(n1181), .ZN(n1167) );
XNOR2_X1 U1019 ( .A(n1266), .B(G478), .ZN(n1181) );
NAND2_X1 U1020 ( .A1(n1094), .A2(n1188), .ZN(n1266) );
INV_X1 U1021 ( .A(G902), .ZN(n1188) );
XNOR2_X1 U1022 ( .A(n1267), .B(n1268), .ZN(n1094) );
XOR2_X1 U1023 ( .A(G116), .B(n1269), .Z(n1268) );
XOR2_X1 U1024 ( .A(G134), .B(G122), .Z(n1269) );
XOR2_X1 U1025 ( .A(n1270), .B(n1241), .Z(n1267) );
XOR2_X1 U1026 ( .A(G107), .B(KEYINPUT10), .Z(n1241) );
XOR2_X1 U1027 ( .A(n1271), .B(n1247), .Z(n1270) );
XNOR2_X1 U1028 ( .A(n1265), .B(G128), .ZN(n1247) );
INV_X1 U1029 ( .A(G143), .ZN(n1265) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1204), .ZN(n1271) );
AND2_X1 U1031 ( .A1(G234), .A2(n1082), .ZN(n1204) );
INV_X1 U1032 ( .A(G953), .ZN(n1082) );
endmodule


