//Key = 0100110000101111110000000010100000101000011111001011111110111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;

XOR2_X1 U754 ( .A(n1035), .B(n1036), .Z(G9) );
NOR3_X1 U755 ( .A1(n1037), .A2(KEYINPUT22), .A3(n1038), .ZN(n1036) );
XNOR2_X1 U756 ( .A(G107), .B(KEYINPUT54), .ZN(n1035) );
NOR2_X1 U757 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR3_X1 U758 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1040) );
AND4_X1 U759 ( .A1(n1042), .A2(n1043), .A3(KEYINPUT1), .A4(n1044), .ZN(n1039) );
NOR4_X1 U760 ( .A1(G953), .A2(n1041), .A3(n1045), .A4(n1046), .ZN(n1044) );
NOR4_X1 U761 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR2_X1 U762 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NOR2_X1 U763 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U764 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1051) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1045) );
INV_X1 U769 ( .A(n1065), .ZN(n1064) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1048), .ZN(n1067) );
INV_X1 U772 ( .A(n1069), .ZN(n1048) );
NOR2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U774 ( .A1(KEYINPUT35), .A2(n1072), .ZN(n1071) );
NOR3_X1 U775 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1070) );
NOR2_X1 U776 ( .A1(n1076), .A2(n1049), .ZN(n1066) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
AND4_X1 U778 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1041) );
NOR4_X1 U779 ( .A1(n1083), .A2(n1084), .A3(n1074), .A4(n1085), .ZN(n1082) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U781 ( .A1(KEYINPUT29), .A2(n1088), .ZN(n1087) );
XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(n1081) );
NAND2_X1 U783 ( .A1(KEYINPUT35), .A2(n1091), .ZN(n1043) );
NAND3_X1 U784 ( .A1(n1092), .A2(n1069), .A3(n1065), .ZN(n1091) );
NOR3_X1 U785 ( .A1(n1058), .A2(n1054), .A3(n1050), .ZN(n1065) );
XOR2_X1 U786 ( .A(n1093), .B(n1094), .Z(G72) );
XOR2_X1 U787 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U788 ( .A1(n1097), .A2(G953), .ZN(n1096) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
INV_X1 U790 ( .A(n1100), .ZN(n1099) );
AND2_X1 U791 ( .A1(G227), .A2(G900), .ZN(n1098) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1093) );
XOR2_X1 U793 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U794 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U795 ( .A1(KEYINPUT31), .A2(n1107), .ZN(n1106) );
XNOR2_X1 U796 ( .A(G134), .B(n1108), .ZN(n1107) );
XNOR2_X1 U797 ( .A(n1109), .B(KEYINPUT28), .ZN(n1103) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(G69) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U800 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U802 ( .A(n1117), .B(KEYINPUT19), .Z(n1115) );
NAND4_X1 U803 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1117) );
NAND2_X1 U804 ( .A1(n1100), .A2(n1122), .ZN(n1112) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1122) );
XOR2_X1 U806 ( .A(G953), .B(KEYINPUT21), .Z(n1100) );
NAND3_X1 U807 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1110) );
XOR2_X1 U808 ( .A(n1126), .B(KEYINPUT33), .Z(n1125) );
NAND2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
OR2_X1 U810 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U811 ( .A(n1129), .B(n1130), .ZN(n1127) );
NAND2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1123) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(G66) );
NOR3_X1 U814 ( .A1(n1089), .A2(n1135), .A3(n1136), .ZN(n1134) );
NOR3_X1 U815 ( .A1(n1137), .A2(n1090), .A3(n1138), .ZN(n1136) );
INV_X1 U816 ( .A(n1139), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1139), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1042), .A2(n1090), .ZN(n1140) );
NOR2_X1 U819 ( .A1(n1133), .A2(n1141), .ZN(G63) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U821 ( .A(KEYINPUT44), .B(n1144), .Z(n1143) );
AND2_X1 U822 ( .A1(G478), .A2(n1145), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1133), .A2(n1146), .ZN(G60) );
XOR2_X1 U824 ( .A(n1147), .B(n1148), .Z(n1146) );
AND2_X1 U825 ( .A1(G475), .A2(n1145), .ZN(n1147) );
XNOR2_X1 U826 ( .A(G104), .B(n1149), .ZN(G6) );
NOR2_X1 U827 ( .A1(n1133), .A2(n1150), .ZN(G57) );
XOR2_X1 U828 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U829 ( .A1(KEYINPUT38), .A2(n1153), .ZN(n1152) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(n1153) );
AND2_X1 U831 ( .A1(G472), .A2(n1145), .ZN(n1155) );
NAND3_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
NAND2_X1 U833 ( .A1(KEYINPUT6), .A2(n1159), .ZN(n1158) );
OR3_X1 U834 ( .A1(n1159), .A2(KEYINPUT6), .A3(n1160), .ZN(n1157) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NAND2_X1 U836 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U837 ( .A(KEYINPUT6), .ZN(n1163) );
XNOR2_X1 U838 ( .A(n1159), .B(KEYINPUT24), .ZN(n1162) );
XOR2_X1 U839 ( .A(n1164), .B(n1165), .Z(n1159) );
NOR2_X1 U840 ( .A1(KEYINPUT0), .A2(n1166), .ZN(n1165) );
NOR2_X1 U841 ( .A1(n1133), .A2(n1167), .ZN(G54) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
AND2_X1 U843 ( .A1(G469), .A2(n1145), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
XOR2_X1 U845 ( .A(KEYINPUT9), .B(n1172), .Z(n1171) );
NOR2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(KEYINPUT57), .Z(n1173) );
AND2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
XOR2_X1 U849 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U850 ( .A(n1178), .B(n1166), .ZN(n1174) );
XOR2_X1 U851 ( .A(G131), .B(n1179), .Z(n1166) );
NAND2_X1 U852 ( .A1(KEYINPUT51), .A2(n1180), .ZN(n1178) );
XOR2_X1 U853 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U854 ( .A(KEYINPUT11), .B(n1183), .Z(n1182) );
NOR2_X1 U855 ( .A1(n1133), .A2(n1184), .ZN(G51) );
NOR2_X1 U856 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U857 ( .A(KEYINPUT49), .B(n1187), .Z(n1186) );
AND2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1188), .ZN(n1185) );
XNOR2_X1 U860 ( .A(n1190), .B(n1191), .ZN(n1188) );
XNOR2_X1 U861 ( .A(G125), .B(n1192), .ZN(n1190) );
NOR2_X1 U862 ( .A1(KEYINPUT39), .A2(n1164), .ZN(n1192) );
NOR2_X1 U863 ( .A1(n1138), .A2(n1193), .ZN(n1189) );
INV_X1 U864 ( .A(n1145), .ZN(n1138) );
NOR2_X1 U865 ( .A1(n1194), .A2(n1042), .ZN(n1145) );
AND4_X1 U866 ( .A1(n1195), .A2(n1196), .A3(n1097), .A4(n1197), .ZN(n1042) );
AND3_X1 U867 ( .A1(n1119), .A2(n1121), .A3(n1120), .ZN(n1197) );
AND4_X1 U868 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1097) );
AND4_X1 U869 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NAND2_X1 U870 ( .A1(n1206), .A2(n1207), .ZN(n1200) );
NAND2_X1 U871 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND3_X1 U872 ( .A1(n1210), .A2(n1211), .A3(n1078), .ZN(n1209) );
XNOR2_X1 U873 ( .A(KEYINPUT30), .B(n1212), .ZN(n1211) );
XOR2_X1 U874 ( .A(KEYINPUT58), .B(n1213), .Z(n1208) );
NAND2_X1 U875 ( .A1(n1214), .A2(n1215), .ZN(n1199) );
XNOR2_X1 U876 ( .A(KEYINPUT20), .B(n1049), .ZN(n1215) );
NAND4_X1 U877 ( .A1(n1092), .A2(n1056), .A3(n1216), .A4(n1217), .ZN(n1198) );
NAND2_X1 U878 ( .A1(KEYINPUT13), .A2(n1218), .ZN(n1217) );
NAND2_X1 U879 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
INV_X1 U880 ( .A(KEYINPUT13), .ZN(n1220) );
NAND3_X1 U881 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1219) );
XNOR2_X1 U882 ( .A(KEYINPUT55), .B(n1118), .ZN(n1196) );
INV_X1 U883 ( .A(n1116), .ZN(n1195) );
NAND4_X1 U884 ( .A1(n1224), .A2(n1225), .A3(n1149), .A4(n1226), .ZN(n1116) );
NAND4_X1 U885 ( .A1(n1055), .A2(n1227), .A3(n1069), .A4(n1060), .ZN(n1149) );
NAND2_X1 U886 ( .A1(n1228), .A2(n1092), .ZN(n1225) );
XOR2_X1 U887 ( .A(n1229), .B(KEYINPUT5), .Z(n1228) );
OR2_X1 U888 ( .A1(n1037), .A2(n1038), .ZN(n1224) );
NAND3_X1 U889 ( .A1(n1069), .A2(n1060), .A3(n1056), .ZN(n1037) );
NOR2_X1 U890 ( .A1(n1230), .A2(G952), .ZN(n1133) );
XNOR2_X1 U891 ( .A(G146), .B(n1205), .ZN(G48) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1055), .ZN(n1205) );
NAND2_X1 U893 ( .A1(n1232), .A2(n1233), .ZN(G45) );
OR2_X1 U894 ( .A1(n1204), .A2(G143), .ZN(n1233) );
XOR2_X1 U895 ( .A(n1234), .B(KEYINPUT18), .Z(n1232) );
NAND2_X1 U896 ( .A1(G143), .A2(n1204), .ZN(n1234) );
NAND3_X1 U897 ( .A1(n1078), .A2(n1210), .A3(n1235), .ZN(n1204) );
NOR3_X1 U898 ( .A1(n1072), .A2(n1236), .A3(n1237), .ZN(n1235) );
XNOR2_X1 U899 ( .A(n1203), .B(n1238), .ZN(G42) );
NOR2_X1 U900 ( .A1(KEYINPUT7), .A2(n1239), .ZN(n1238) );
NAND4_X1 U901 ( .A1(n1210), .A2(n1206), .A3(n1055), .A4(n1077), .ZN(n1203) );
XOR2_X1 U902 ( .A(G137), .B(n1240), .Z(G39) );
AND2_X1 U903 ( .A1(n1206), .A2(n1214), .ZN(n1240) );
NOR2_X1 U904 ( .A1(n1058), .A2(n1218), .ZN(n1214) );
INV_X1 U905 ( .A(n1079), .ZN(n1058) );
NAND2_X1 U906 ( .A1(n1241), .A2(n1242), .ZN(G36) );
NAND2_X1 U907 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XNOR2_X1 U908 ( .A(G134), .B(KEYINPUT48), .ZN(n1243) );
XOR2_X1 U909 ( .A(KEYINPUT53), .B(n1245), .Z(n1241) );
NOR2_X1 U910 ( .A1(n1244), .A2(n1246), .ZN(n1245) );
XNOR2_X1 U911 ( .A(KEYINPUT8), .B(n1247), .ZN(n1246) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1206), .ZN(n1244) );
AND3_X1 U913 ( .A1(n1210), .A2(n1056), .A3(n1078), .ZN(n1213) );
XOR2_X1 U914 ( .A(G131), .B(n1248), .Z(G33) );
NOR3_X1 U915 ( .A1(n1249), .A2(n1212), .A3(n1049), .ZN(n1248) );
INV_X1 U916 ( .A(n1206), .ZN(n1049) );
NOR3_X1 U917 ( .A1(n1074), .A2(n1084), .A3(n1075), .ZN(n1206) );
INV_X1 U918 ( .A(n1073), .ZN(n1084) );
INV_X1 U919 ( .A(n1055), .ZN(n1212) );
NAND3_X1 U920 ( .A1(n1250), .A2(n1251), .A3(n1078), .ZN(n1249) );
OR2_X1 U921 ( .A1(n1252), .A2(n1210), .ZN(n1251) );
NAND2_X1 U922 ( .A1(n1253), .A2(n1252), .ZN(n1250) );
INV_X1 U923 ( .A(KEYINPUT15), .ZN(n1252) );
NAND2_X1 U924 ( .A1(n1221), .A2(n1222), .ZN(n1253) );
XNOR2_X1 U925 ( .A(G128), .B(n1254), .ZN(G30) );
NAND2_X1 U926 ( .A1(n1231), .A2(n1056), .ZN(n1254) );
NOR2_X1 U927 ( .A1(n1218), .A2(n1072), .ZN(n1231) );
NAND2_X1 U928 ( .A1(n1223), .A2(n1210), .ZN(n1218) );
NOR2_X1 U929 ( .A1(n1222), .A2(n1255), .ZN(n1210) );
XNOR2_X1 U930 ( .A(G101), .B(n1226), .ZN(G3) );
NAND4_X1 U931 ( .A1(n1079), .A2(n1078), .A3(n1227), .A4(n1060), .ZN(n1226) );
INV_X1 U932 ( .A(n1038), .ZN(n1227) );
XNOR2_X1 U933 ( .A(n1256), .B(n1257), .ZN(G27) );
NOR2_X1 U934 ( .A1(KEYINPUT46), .A2(n1202), .ZN(n1257) );
NAND4_X1 U935 ( .A1(n1055), .A2(n1080), .A3(n1258), .A4(n1077), .ZN(n1202) );
NOR2_X1 U936 ( .A1(n1255), .A2(n1072), .ZN(n1258) );
INV_X1 U937 ( .A(n1221), .ZN(n1255) );
NAND2_X1 U938 ( .A1(n1050), .A2(n1259), .ZN(n1221) );
NAND3_X1 U939 ( .A1(G902), .A2(n1260), .A3(n1101), .ZN(n1259) );
NOR2_X1 U940 ( .A1(n1261), .A2(G900), .ZN(n1101) );
INV_X1 U941 ( .A(n1054), .ZN(n1080) );
XNOR2_X1 U942 ( .A(G122), .B(n1119), .ZN(G24) );
NAND4_X1 U943 ( .A1(n1262), .A2(n1069), .A3(n1263), .A4(n1264), .ZN(n1119) );
NOR2_X1 U944 ( .A1(n1265), .A2(n1266), .ZN(n1069) );
XNOR2_X1 U945 ( .A(G119), .B(n1120), .ZN(G21) );
NAND3_X1 U946 ( .A1(n1079), .A2(n1223), .A3(n1262), .ZN(n1120) );
NOR2_X1 U947 ( .A1(n1267), .A2(n1268), .ZN(n1223) );
XNOR2_X1 U948 ( .A(G116), .B(n1121), .ZN(G18) );
NAND3_X1 U949 ( .A1(n1078), .A2(n1056), .A3(n1262), .ZN(n1121) );
NOR2_X1 U950 ( .A1(n1264), .A2(n1237), .ZN(n1056) );
INV_X1 U951 ( .A(n1263), .ZN(n1237) );
XNOR2_X1 U952 ( .A(G113), .B(n1118), .ZN(G15) );
NAND3_X1 U953 ( .A1(n1078), .A2(n1055), .A3(n1262), .ZN(n1118) );
NOR2_X1 U954 ( .A1(n1054), .A2(n1038), .ZN(n1262) );
NAND2_X1 U955 ( .A1(n1092), .A2(n1269), .ZN(n1038) );
INV_X1 U956 ( .A(n1072), .ZN(n1092) );
NAND2_X1 U957 ( .A1(n1270), .A2(n1062), .ZN(n1054) );
INV_X1 U958 ( .A(n1061), .ZN(n1270) );
NOR2_X1 U959 ( .A1(n1263), .A2(n1236), .ZN(n1055) );
INV_X1 U960 ( .A(n1264), .ZN(n1236) );
NOR2_X1 U961 ( .A1(n1267), .A2(n1265), .ZN(n1078) );
XOR2_X1 U962 ( .A(G110), .B(n1271), .Z(G12) );
NOR2_X1 U963 ( .A1(n1072), .A2(n1229), .ZN(n1271) );
NAND4_X1 U964 ( .A1(n1079), .A2(n1077), .A3(n1060), .A4(n1269), .ZN(n1229) );
NAND2_X1 U965 ( .A1(n1050), .A2(n1272), .ZN(n1269) );
NAND4_X1 U966 ( .A1(G902), .A2(n1131), .A3(n1260), .A4(n1132), .ZN(n1272) );
INV_X1 U967 ( .A(G898), .ZN(n1132) );
INV_X1 U968 ( .A(n1261), .ZN(n1131) );
XOR2_X1 U969 ( .A(n1230), .B(KEYINPUT62), .Z(n1261) );
NAND3_X1 U970 ( .A1(n1260), .A2(n1230), .A3(G952), .ZN(n1050) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1260) );
INV_X1 U972 ( .A(n1222), .ZN(n1060) );
NAND2_X1 U973 ( .A1(n1061), .A2(n1062), .ZN(n1222) );
NAND2_X1 U974 ( .A1(n1273), .A2(n1274), .ZN(n1062) );
XNOR2_X1 U975 ( .A(G221), .B(KEYINPUT60), .ZN(n1273) );
XNOR2_X1 U976 ( .A(n1275), .B(G469), .ZN(n1061) );
NAND2_X1 U977 ( .A1(n1276), .A2(n1194), .ZN(n1275) );
XOR2_X1 U978 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U979 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U980 ( .A(n1176), .B(KEYINPUT17), .Z(n1280) );
NAND2_X1 U981 ( .A1(G227), .A2(n1230), .ZN(n1176) );
NAND2_X1 U982 ( .A1(KEYINPUT56), .A2(n1177), .ZN(n1279) );
XNOR2_X1 U983 ( .A(n1181), .B(n1281), .ZN(n1277) );
XNOR2_X1 U984 ( .A(n1282), .B(n1283), .ZN(n1181) );
XOR2_X1 U985 ( .A(G101), .B(n1109), .Z(n1283) );
NOR2_X1 U986 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1109) );
XNOR2_X1 U987 ( .A(G104), .B(G107), .ZN(n1282) );
NOR2_X1 U988 ( .A1(n1266), .A2(n1268), .ZN(n1077) );
INV_X1 U989 ( .A(n1265), .ZN(n1268) );
NAND2_X1 U990 ( .A1(n1284), .A2(n1285), .ZN(n1265) );
NAND2_X1 U991 ( .A1(n1089), .A2(n1286), .ZN(n1285) );
XOR2_X1 U992 ( .A(KEYINPUT12), .B(n1287), .Z(n1284) );
NOR2_X1 U993 ( .A1(n1089), .A2(n1286), .ZN(n1287) );
XNOR2_X1 U994 ( .A(KEYINPUT36), .B(n1090), .ZN(n1286) );
NAND2_X1 U995 ( .A1(G217), .A2(n1274), .ZN(n1090) );
NAND2_X1 U996 ( .A1(G234), .A2(n1194), .ZN(n1274) );
NOR2_X1 U997 ( .A1(n1139), .A2(G902), .ZN(n1089) );
XNOR2_X1 U998 ( .A(n1288), .B(n1289), .ZN(n1139) );
XOR2_X1 U999 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1000 ( .A(n1292), .B(n1293), .Z(n1291) );
NOR2_X1 U1001 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U1002 ( .A(n1296), .B(KEYINPUT4), .Z(n1295) );
NAND2_X1 U1003 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NOR2_X1 U1004 ( .A1(n1298), .A2(n1297), .ZN(n1294) );
XOR2_X1 U1005 ( .A(KEYINPUT27), .B(G119), .Z(n1297) );
AND3_X1 U1006 ( .A1(G221), .A2(n1230), .A3(G234), .ZN(n1292) );
XOR2_X1 U1007 ( .A(KEYINPUT26), .B(G146), .Z(n1290) );
XNOR2_X1 U1008 ( .A(n1177), .B(n1299), .ZN(n1288) );
XNOR2_X1 U1009 ( .A(n1300), .B(n1301), .ZN(n1299) );
NOR2_X1 U1010 ( .A1(G125), .A2(KEYINPUT32), .ZN(n1301) );
NAND2_X1 U1011 ( .A1(KEYINPUT59), .A2(n1108), .ZN(n1300) );
XNOR2_X1 U1012 ( .A(G110), .B(n1239), .ZN(n1177) );
INV_X1 U1013 ( .A(n1267), .ZN(n1266) );
XOR2_X1 U1014 ( .A(n1086), .B(n1088), .Z(n1267) );
XNOR2_X1 U1015 ( .A(G472), .B(KEYINPUT16), .ZN(n1088) );
NAND2_X1 U1016 ( .A1(n1302), .A2(n1194), .ZN(n1086) );
XOR2_X1 U1017 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1018 ( .A(n1160), .B(n1305), .ZN(n1304) );
XNOR2_X1 U1019 ( .A(G128), .B(KEYINPUT3), .ZN(n1305) );
AND2_X1 U1020 ( .A1(n1306), .A2(n1307), .ZN(n1160) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U1022 ( .A(KEYINPUT52), .B(n1310), .ZN(n1306) );
XOR2_X1 U1023 ( .A(n1151), .B(n1281), .Z(n1303) );
XNOR2_X1 U1024 ( .A(n1311), .B(n1179), .ZN(n1281) );
XNOR2_X1 U1025 ( .A(n1247), .B(n1312), .ZN(n1179) );
NOR2_X1 U1026 ( .A1(KEYINPUT63), .A2(n1108), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(G137), .B(KEYINPUT42), .ZN(n1108) );
XOR2_X1 U1028 ( .A(n1313), .B(G101), .Z(n1151) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1314), .ZN(n1313) );
NOR2_X1 U1030 ( .A1(n1263), .A2(n1264), .ZN(n1079) );
XNOR2_X1 U1031 ( .A(n1315), .B(G475), .ZN(n1264) );
OR2_X1 U1032 ( .A1(n1148), .A2(G902), .ZN(n1315) );
XNOR2_X1 U1033 ( .A(n1316), .B(n1317), .ZN(n1148) );
XOR2_X1 U1034 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1035 ( .A(G104), .B(G122), .ZN(n1319) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1314), .ZN(n1318) );
NOR2_X1 U1037 ( .A1(G953), .A2(G237), .ZN(n1314) );
XNOR2_X1 U1038 ( .A(n1105), .B(n1308), .ZN(n1316) );
XOR2_X1 U1039 ( .A(n1311), .B(n1320), .Z(n1105) );
XNOR2_X1 U1040 ( .A(n1239), .B(G125), .ZN(n1320) );
INV_X1 U1041 ( .A(G140), .ZN(n1239) );
XNOR2_X1 U1042 ( .A(G131), .B(n1183), .ZN(n1311) );
XNOR2_X1 U1043 ( .A(n1321), .B(n1322), .ZN(n1263) );
XOR2_X1 U1044 ( .A(KEYINPUT37), .B(G478), .Z(n1322) );
NAND2_X1 U1045 ( .A1(n1142), .A2(n1194), .ZN(n1321) );
XNOR2_X1 U1046 ( .A(n1323), .B(n1324), .ZN(n1142) );
XOR2_X1 U1047 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1048 ( .A(n1327), .B(n1328), .ZN(n1326) );
NAND2_X1 U1049 ( .A1(KEYINPUT10), .A2(n1247), .ZN(n1328) );
INV_X1 U1050 ( .A(G134), .ZN(n1247) );
NAND2_X1 U1051 ( .A1(KEYINPUT41), .A2(n1329), .ZN(n1327) );
XNOR2_X1 U1052 ( .A(KEYINPUT34), .B(n1330), .ZN(n1329) );
NAND3_X1 U1053 ( .A1(G217), .A2(n1230), .A3(G234), .ZN(n1325) );
XOR2_X1 U1054 ( .A(n1331), .B(n1332), .Z(n1323) );
XNOR2_X1 U1055 ( .A(G143), .B(n1298), .ZN(n1332) );
INV_X1 U1056 ( .A(G128), .ZN(n1298) );
XNOR2_X1 U1057 ( .A(G116), .B(G107), .ZN(n1331) );
NAND2_X1 U1058 ( .A1(n1073), .A2(n1333), .ZN(n1072) );
OR2_X1 U1059 ( .A1(n1075), .A2(n1074), .ZN(n1333) );
NOR2_X1 U1060 ( .A1(n1334), .A2(n1335), .ZN(n1074) );
XOR2_X1 U1061 ( .A(n1083), .B(KEYINPUT47), .Z(n1075) );
AND2_X1 U1062 ( .A1(n1335), .A2(n1334), .ZN(n1083) );
NAND2_X1 U1063 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
XOR2_X1 U1064 ( .A(n1338), .B(n1339), .Z(n1337) );
XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n1256), .ZN(n1339) );
INV_X1 U1066 ( .A(G125), .ZN(n1256) );
XNOR2_X1 U1067 ( .A(n1164), .B(n1191), .ZN(n1338) );
XNOR2_X1 U1068 ( .A(n1340), .B(n1341), .ZN(n1191) );
XOR2_X1 U1069 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1070 ( .A(KEYINPUT2), .B(n1344), .Z(n1343) );
AND2_X1 U1071 ( .A1(n1230), .A2(G224), .ZN(n1344) );
INV_X1 U1072 ( .A(G953), .ZN(n1230) );
NOR2_X1 U1073 ( .A1(n1129), .A2(KEYINPUT25), .ZN(n1342) );
AND2_X1 U1074 ( .A1(n1310), .A2(n1345), .ZN(n1129) );
NAND2_X1 U1075 ( .A1(n1346), .A2(n1309), .ZN(n1345) );
XNOR2_X1 U1076 ( .A(KEYINPUT50), .B(n1308), .ZN(n1346) );
OR2_X1 U1077 ( .A1(n1309), .A2(n1308), .ZN(n1310) );
XNOR2_X1 U1078 ( .A(G113), .B(KEYINPUT14), .ZN(n1308) );
XOR2_X1 U1079 ( .A(G116), .B(G119), .Z(n1309) );
XOR2_X1 U1080 ( .A(n1130), .B(n1128), .Z(n1340) );
XNOR2_X1 U1081 ( .A(G110), .B(n1330), .ZN(n1128) );
INV_X1 U1082 ( .A(G122), .ZN(n1330) );
NAND2_X1 U1083 ( .A1(n1347), .A2(n1348), .ZN(n1130) );
NAND2_X1 U1084 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
INV_X1 U1085 ( .A(G107), .ZN(n1350) );
XOR2_X1 U1086 ( .A(KEYINPUT40), .B(n1351), .Z(n1349) );
NAND2_X1 U1087 ( .A1(n1352), .A2(G107), .ZN(n1347) );
XOR2_X1 U1088 ( .A(KEYINPUT43), .B(n1351), .Z(n1352) );
XOR2_X1 U1089 ( .A(G101), .B(G104), .Z(n1351) );
XOR2_X1 U1090 ( .A(G128), .B(n1183), .Z(n1164) );
XOR2_X1 U1091 ( .A(G146), .B(G143), .Z(n1183) );
XNOR2_X1 U1092 ( .A(KEYINPUT45), .B(n1194), .ZN(n1336) );
INV_X1 U1093 ( .A(n1193), .ZN(n1335) );
NAND2_X1 U1094 ( .A1(G210), .A2(n1353), .ZN(n1193) );
NAND2_X1 U1095 ( .A1(G214), .A2(n1353), .ZN(n1073) );
NAND2_X1 U1096 ( .A1(n1354), .A2(n1194), .ZN(n1353) );
INV_X1 U1097 ( .A(G902), .ZN(n1194) );
INV_X1 U1098 ( .A(G237), .ZN(n1354) );
endmodule


