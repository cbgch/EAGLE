//Key = 1111111001101000111111110011111000010000100110001010101011001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;

XNOR2_X1 U735 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR3_X1 U737 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
AND4_X1 U739 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1034) );
NAND3_X1 U740 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1031) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1043), .ZN(n1042) );
NAND2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U743 ( .A1(n1036), .A2(n1046), .A3(n1037), .ZN(n1045) );
NAND3_X1 U744 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U745 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U746 ( .A1(n1052), .A2(n1053), .ZN(n1048) );
NAND2_X1 U747 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U748 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U749 ( .A1(n1038), .A2(n1035), .ZN(n1047) );
INV_X1 U750 ( .A(KEYINPUT46), .ZN(n1035) );
NAND3_X1 U751 ( .A1(n1052), .A2(n1058), .A3(n1050), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U753 ( .A1(n1036), .A2(n1061), .ZN(n1060) );
OR2_X1 U754 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U755 ( .A1(n1037), .A2(n1064), .ZN(n1059) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U757 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U758 ( .A(n1069), .ZN(n1039) );
NOR3_X1 U759 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1029) );
INV_X1 U760 ( .A(n1040), .ZN(n1070) );
NAND2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1040) );
NOR4_X1 U762 ( .A1(n1057), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XNOR2_X1 U763 ( .A(n1076), .B(n1077), .ZN(n1075) );
NAND2_X1 U764 ( .A1(KEYINPUT12), .A2(n1078), .ZN(n1076) );
AND2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NOR4_X1 U766 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1071) );
XNOR2_X1 U767 ( .A(n1085), .B(n1086), .ZN(n1084) );
XOR2_X1 U768 ( .A(n1087), .B(n1088), .Z(n1081) );
XNOR2_X1 U769 ( .A(KEYINPUT43), .B(n1089), .ZN(n1088) );
XOR2_X1 U770 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U771 ( .A1(n1092), .A2(n1041), .ZN(n1091) );
AND2_X1 U772 ( .A1(G227), .A2(G900), .ZN(n1092) );
NAND2_X1 U773 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U774 ( .A1(n1095), .A2(n1041), .ZN(n1094) );
XOR2_X1 U775 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U776 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NAND3_X1 U777 ( .A1(n1097), .A2(n1100), .A3(G953), .ZN(n1093) );
XNOR2_X1 U778 ( .A(KEYINPUT15), .B(n1101), .ZN(n1100) );
AND2_X1 U779 ( .A1(KEYINPUT4), .A2(n1102), .ZN(n1097) );
XOR2_X1 U780 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U781 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U782 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U783 ( .A(n1109), .ZN(n1108) );
NOR2_X1 U784 ( .A1(KEYINPUT51), .A2(n1110), .ZN(n1107) );
NOR2_X1 U785 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U786 ( .A1(G140), .A2(n1113), .ZN(n1105) );
NOR2_X1 U787 ( .A1(n1114), .A2(n1112), .ZN(n1113) );
INV_X1 U788 ( .A(KEYINPUT0), .ZN(n1112) );
NOR2_X1 U789 ( .A1(KEYINPUT51), .A2(n1109), .ZN(n1114) );
XOR2_X1 U790 ( .A(G125), .B(KEYINPUT24), .Z(n1109) );
XOR2_X1 U791 ( .A(n1115), .B(n1116), .Z(G69) );
NAND2_X1 U792 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1117) );
NAND2_X1 U794 ( .A1(KEYINPUT5), .A2(n1118), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U798 ( .A(n1125), .B(KEYINPUT26), .ZN(n1123) );
XNOR2_X1 U799 ( .A(KEYINPUT1), .B(n1041), .ZN(n1121) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1119) );
NAND2_X1 U801 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1126) );
XOR2_X1 U803 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U804 ( .A1(n1133), .A2(KEYINPUT41), .ZN(n1131) );
INV_X1 U805 ( .A(n1134), .ZN(n1133) );
XOR2_X1 U806 ( .A(KEYINPUT31), .B(n1135), .Z(n1129) );
NOR2_X1 U807 ( .A1(n1136), .A2(n1137), .ZN(G66) );
NOR3_X1 U808 ( .A1(n1085), .A2(n1138), .A3(n1139), .ZN(n1137) );
NOR3_X1 U809 ( .A1(n1140), .A2(n1086), .A3(n1141), .ZN(n1139) );
INV_X1 U810 ( .A(n1142), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1143), .A2(n1142), .ZN(n1138) );
NOR2_X1 U812 ( .A1(n1144), .A2(n1086), .ZN(n1143) );
INV_X1 U813 ( .A(n1033), .ZN(n1144) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1145), .ZN(G63) );
XOR2_X1 U815 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U816 ( .A1(n1079), .A2(n1141), .ZN(n1146) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1148), .ZN(G60) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U819 ( .A1(n1151), .A2(n1141), .ZN(n1149) );
XNOR2_X1 U820 ( .A(G104), .B(n1152), .ZN(G6) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1153), .ZN(G57) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(n1153) );
XNOR2_X1 U823 ( .A(n1156), .B(n1157), .ZN(n1155) );
XOR2_X1 U824 ( .A(n1158), .B(n1159), .Z(n1154) );
XNOR2_X1 U825 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U826 ( .A1(n1141), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U827 ( .A(KEYINPUT50), .B(n1089), .ZN(n1162) );
NAND2_X1 U828 ( .A1(KEYINPUT18), .A2(n1163), .ZN(n1158) );
NOR2_X1 U829 ( .A1(n1136), .A2(n1164), .ZN(G54) );
XOR2_X1 U830 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U831 ( .A1(KEYINPUT58), .A2(n1167), .ZN(n1166) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1141), .ZN(n1165) );
NOR2_X1 U833 ( .A1(n1136), .A2(n1169), .ZN(G51) );
XOR2_X1 U834 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U835 ( .A1(n1077), .A2(n1141), .ZN(n1171) );
NAND2_X1 U836 ( .A1(G902), .A2(n1033), .ZN(n1141) );
NAND4_X1 U837 ( .A1(n1172), .A2(n1125), .A3(n1098), .A4(n1124), .ZN(n1033) );
AND4_X1 U838 ( .A1(n1173), .A2(n1152), .A3(n1174), .A4(n1028), .ZN(n1124) );
NAND3_X1 U839 ( .A1(n1052), .A2(n1062), .A3(n1175), .ZN(n1028) );
NAND3_X1 U840 ( .A1(n1175), .A2(n1052), .A3(n1063), .ZN(n1152) );
NAND3_X1 U841 ( .A1(n1175), .A2(n1176), .A3(n1037), .ZN(n1173) );
AND4_X1 U842 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1098) );
AND3_X1 U843 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1185), .ZN(n1179) );
NAND2_X1 U845 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U846 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
AND3_X1 U847 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1125) );
NOR3_X1 U848 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1192) );
NOR2_X1 U849 ( .A1(n1054), .A2(n1196), .ZN(n1195) );
NOR2_X1 U850 ( .A1(n1184), .A2(n1197), .ZN(n1194) );
NAND4_X1 U851 ( .A1(n1037), .A2(n1189), .A3(n1198), .A4(n1199), .ZN(n1197) );
NOR2_X1 U852 ( .A1(n1200), .A2(n1199), .ZN(n1193) );
INV_X1 U853 ( .A(KEYINPUT56), .ZN(n1199) );
XOR2_X1 U854 ( .A(n1099), .B(KEYINPUT14), .Z(n1172) );
NAND2_X1 U855 ( .A1(n1201), .A2(n1202), .ZN(n1099) );
INV_X1 U856 ( .A(n1203), .ZN(n1202) );
XNOR2_X1 U857 ( .A(n1036), .B(KEYINPUT19), .ZN(n1201) );
INV_X1 U858 ( .A(n1083), .ZN(n1036) );
NAND2_X1 U859 ( .A1(KEYINPUT35), .A2(n1204), .ZN(n1170) );
XOR2_X1 U860 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U861 ( .A(KEYINPUT55), .B(n1207), .Z(n1206) );
NOR2_X1 U862 ( .A1(n1041), .A2(G952), .ZN(n1136) );
XOR2_X1 U863 ( .A(n1208), .B(n1209), .Z(G48) );
NOR3_X1 U864 ( .A1(n1210), .A2(n1211), .A3(n1054), .ZN(n1209) );
XNOR2_X1 U865 ( .A(n1189), .B(KEYINPUT42), .ZN(n1211) );
XNOR2_X1 U866 ( .A(G146), .B(KEYINPUT40), .ZN(n1208) );
XOR2_X1 U867 ( .A(n1212), .B(n1213), .Z(G45) );
NAND2_X1 U868 ( .A1(KEYINPUT57), .A2(G143), .ZN(n1213) );
NAND2_X1 U869 ( .A1(n1214), .A2(n1184), .ZN(n1212) );
XOR2_X1 U870 ( .A(n1186), .B(KEYINPUT29), .Z(n1214) );
NAND4_X1 U871 ( .A1(n1215), .A2(n1176), .A3(n1082), .A4(n1216), .ZN(n1186) );
NAND2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1219), .A2(n1177), .ZN(n1218) );
XNOR2_X1 U874 ( .A(KEYINPUT59), .B(n1111), .ZN(n1219) );
NAND2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
INV_X1 U876 ( .A(n1177), .ZN(n1221) );
NAND3_X1 U877 ( .A1(n1050), .A2(n1051), .A3(n1188), .ZN(n1177) );
XNOR2_X1 U878 ( .A(G140), .B(n1222), .ZN(n1220) );
XNOR2_X1 U879 ( .A(KEYINPUT38), .B(KEYINPUT21), .ZN(n1222) );
XNOR2_X1 U880 ( .A(G137), .B(n1178), .ZN(G39) );
NAND4_X1 U881 ( .A1(n1050), .A2(n1215), .A3(n1037), .A4(n1189), .ZN(n1178) );
XNOR2_X1 U882 ( .A(G134), .B(n1181), .ZN(G36) );
NAND3_X1 U883 ( .A1(n1215), .A2(n1062), .A3(n1038), .ZN(n1181) );
XOR2_X1 U884 ( .A(n1183), .B(n1223), .Z(G33) );
NAND2_X1 U885 ( .A1(KEYINPUT22), .A2(G131), .ZN(n1223) );
NAND2_X1 U886 ( .A1(n1188), .A2(n1038), .ZN(n1183) );
AND2_X1 U887 ( .A1(n1050), .A2(n1176), .ZN(n1038) );
AND2_X1 U888 ( .A1(n1056), .A2(n1224), .ZN(n1050) );
XOR2_X1 U889 ( .A(KEYINPUT54), .B(n1057), .Z(n1224) );
INV_X1 U890 ( .A(n1210), .ZN(n1188) );
NAND2_X1 U891 ( .A1(n1215), .A2(n1063), .ZN(n1210) );
XNOR2_X1 U892 ( .A(G128), .B(n1182), .ZN(G30) );
NAND4_X1 U893 ( .A1(n1215), .A2(n1189), .A3(n1062), .A4(n1184), .ZN(n1182) );
AND2_X1 U894 ( .A1(n1225), .A2(n1226), .ZN(n1215) );
XNOR2_X1 U895 ( .A(G101), .B(n1227), .ZN(G3) );
NAND3_X1 U896 ( .A1(n1228), .A2(n1037), .A3(n1229), .ZN(n1227) );
AND3_X1 U897 ( .A1(n1225), .A2(n1230), .A3(n1176), .ZN(n1229) );
XNOR2_X1 U898 ( .A(n1184), .B(KEYINPUT27), .ZN(n1228) );
XNOR2_X1 U899 ( .A(n1231), .B(n1232), .ZN(G27) );
NOR2_X1 U900 ( .A1(n1083), .A2(n1203), .ZN(n1232) );
NAND4_X1 U901 ( .A1(n1063), .A2(n1184), .A3(n1051), .A4(n1226), .ZN(n1203) );
NAND2_X1 U902 ( .A1(n1069), .A2(n1233), .ZN(n1226) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1101), .ZN(n1233) );
INV_X1 U904 ( .A(G900), .ZN(n1101) );
XNOR2_X1 U905 ( .A(G122), .B(n1190), .ZN(G24) );
NAND3_X1 U906 ( .A1(n1198), .A2(n1052), .A3(n1235), .ZN(n1190) );
NOR3_X1 U907 ( .A1(n1054), .A2(n1236), .A3(n1237), .ZN(n1235) );
XNOR2_X1 U908 ( .A(G119), .B(n1200), .ZN(G21) );
NAND4_X1 U909 ( .A1(n1037), .A2(n1189), .A3(n1198), .A4(n1184), .ZN(n1200) );
AND2_X1 U910 ( .A1(n1238), .A2(n1239), .ZN(n1189) );
XNOR2_X1 U911 ( .A(KEYINPUT28), .B(n1240), .ZN(n1238) );
XNOR2_X1 U912 ( .A(G116), .B(n1191), .ZN(G18) );
NAND3_X1 U913 ( .A1(n1062), .A2(n1184), .A3(n1241), .ZN(n1191) );
NOR2_X1 U914 ( .A1(n1082), .A2(n1236), .ZN(n1062) );
XNOR2_X1 U915 ( .A(n1242), .B(n1243), .ZN(G15) );
NOR2_X1 U916 ( .A1(n1054), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U917 ( .A(KEYINPUT17), .B(n1196), .ZN(n1244) );
NAND2_X1 U918 ( .A1(n1063), .A2(n1241), .ZN(n1196) );
AND2_X1 U919 ( .A1(n1198), .A2(n1176), .ZN(n1241) );
NAND2_X1 U920 ( .A1(n1245), .A2(n1246), .ZN(n1176) );
OR3_X1 U921 ( .A1(n1240), .A2(n1247), .A3(KEYINPUT32), .ZN(n1246) );
NAND2_X1 U922 ( .A1(KEYINPUT32), .A2(n1052), .ZN(n1245) );
NOR2_X1 U923 ( .A1(n1083), .A2(n1248), .ZN(n1198) );
NAND2_X1 U924 ( .A1(n1068), .A2(n1249), .ZN(n1083) );
NOR2_X1 U925 ( .A1(n1216), .A2(n1237), .ZN(n1063) );
INV_X1 U926 ( .A(n1082), .ZN(n1237) );
XNOR2_X1 U927 ( .A(G110), .B(n1174), .ZN(G12) );
NAND3_X1 U928 ( .A1(n1175), .A2(n1051), .A3(n1037), .ZN(n1174) );
NOR2_X1 U929 ( .A1(n1216), .A2(n1082), .ZN(n1037) );
XOR2_X1 U930 ( .A(n1250), .B(n1151), .Z(n1082) );
INV_X1 U931 ( .A(G475), .ZN(n1151) );
OR2_X1 U932 ( .A1(n1150), .A2(G902), .ZN(n1250) );
XNOR2_X1 U933 ( .A(n1251), .B(n1252), .ZN(n1150) );
XNOR2_X1 U934 ( .A(n1253), .B(n1254), .ZN(n1252) );
NOR2_X1 U935 ( .A1(KEYINPUT49), .A2(n1255), .ZN(n1254) );
XOR2_X1 U936 ( .A(n1256), .B(n1257), .Z(n1255) );
XNOR2_X1 U937 ( .A(n1258), .B(n1259), .ZN(n1257) );
NAND3_X1 U938 ( .A1(n1260), .A2(n1041), .A3(n1261), .ZN(n1258) );
XOR2_X1 U939 ( .A(KEYINPUT13), .B(G214), .Z(n1261) );
XNOR2_X1 U940 ( .A(n1231), .B(n1262), .ZN(n1256) );
XNOR2_X1 U941 ( .A(n1111), .B(G131), .ZN(n1262) );
INV_X1 U942 ( .A(G125), .ZN(n1231) );
XNOR2_X1 U943 ( .A(G113), .B(G122), .ZN(n1251) );
INV_X1 U944 ( .A(n1236), .ZN(n1216) );
NOR2_X1 U945 ( .A1(n1263), .A2(n1073), .ZN(n1236) );
NOR2_X1 U946 ( .A1(n1079), .A2(n1080), .ZN(n1073) );
AND2_X1 U947 ( .A1(n1080), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U948 ( .A(KEYINPUT52), .B(n1079), .ZN(n1264) );
INV_X1 U949 ( .A(G478), .ZN(n1079) );
NOR2_X1 U950 ( .A1(n1147), .A2(G902), .ZN(n1080) );
XNOR2_X1 U951 ( .A(n1265), .B(n1266), .ZN(n1147) );
XOR2_X1 U952 ( .A(n1267), .B(n1268), .Z(n1266) );
AND3_X1 U953 ( .A1(G217), .A2(n1041), .A3(G234), .ZN(n1267) );
XOR2_X1 U954 ( .A(n1269), .B(G143), .Z(n1265) );
NAND2_X1 U955 ( .A1(n1270), .A2(KEYINPUT2), .ZN(n1269) );
XNOR2_X1 U956 ( .A(G107), .B(n1271), .ZN(n1270) );
NOR2_X1 U957 ( .A1(KEYINPUT25), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U958 ( .A(G116), .B(G122), .ZN(n1272) );
NAND2_X1 U959 ( .A1(n1273), .A2(n1274), .ZN(n1051) );
NAND2_X1 U960 ( .A1(n1052), .A2(n1275), .ZN(n1274) );
INV_X1 U961 ( .A(KEYINPUT28), .ZN(n1275) );
NOR2_X1 U962 ( .A1(n1239), .A2(n1240), .ZN(n1052) );
NAND3_X1 U963 ( .A1(n1247), .A2(n1240), .A3(KEYINPUT28), .ZN(n1273) );
XNOR2_X1 U964 ( .A(n1276), .B(n1277), .ZN(n1240) );
INV_X1 U965 ( .A(n1085), .ZN(n1277) );
NOR2_X1 U966 ( .A1(n1142), .A2(G902), .ZN(n1085) );
XNOR2_X1 U967 ( .A(n1278), .B(n1279), .ZN(n1142) );
XOR2_X1 U968 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U969 ( .A(G128), .B(G119), .Z(n1281) );
XOR2_X1 U970 ( .A(G146), .B(G137), .Z(n1280) );
XOR2_X1 U971 ( .A(n1282), .B(n1283), .Z(n1278) );
XOR2_X1 U972 ( .A(G110), .B(n1284), .Z(n1283) );
AND3_X1 U973 ( .A1(G221), .A2(n1041), .A3(G234), .ZN(n1284) );
NAND3_X1 U974 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1282) );
OR2_X1 U975 ( .A1(G125), .A2(KEYINPUT10), .ZN(n1287) );
NAND3_X1 U976 ( .A1(KEYINPUT10), .A2(G125), .A3(n1111), .ZN(n1286) );
NAND2_X1 U977 ( .A1(G140), .A2(n1288), .ZN(n1285) );
NAND2_X1 U978 ( .A1(n1289), .A2(KEYINPUT10), .ZN(n1288) );
XNOR2_X1 U979 ( .A(G125), .B(KEYINPUT48), .ZN(n1289) );
NAND2_X1 U980 ( .A1(KEYINPUT23), .A2(n1086), .ZN(n1276) );
NAND2_X1 U981 ( .A1(G217), .A2(n1290), .ZN(n1086) );
INV_X1 U982 ( .A(n1239), .ZN(n1247) );
XNOR2_X1 U983 ( .A(n1087), .B(n1291), .ZN(n1239) );
NOR2_X1 U984 ( .A1(KEYINPUT7), .A2(n1089), .ZN(n1291) );
INV_X1 U985 ( .A(G472), .ZN(n1089) );
NAND3_X1 U986 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1087) );
NAND3_X1 U987 ( .A1(n1156), .A2(n1295), .A3(KEYINPUT6), .ZN(n1294) );
XOR2_X1 U988 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND2_X1 U989 ( .A1(KEYINPUT60), .A2(n1157), .ZN(n1297) );
NAND2_X1 U990 ( .A1(n1298), .A2(n1299), .ZN(n1292) );
NAND2_X1 U991 ( .A1(KEYINPUT6), .A2(n1156), .ZN(n1299) );
XOR2_X1 U992 ( .A(n1300), .B(n1301), .Z(n1156) );
XOR2_X1 U993 ( .A(n1296), .B(n1302), .Z(n1298) );
NAND2_X1 U994 ( .A1(KEYINPUT60), .A2(n1303), .ZN(n1302) );
INV_X1 U995 ( .A(n1157), .ZN(n1303) );
XOR2_X1 U996 ( .A(G113), .B(n1304), .Z(n1157) );
NAND2_X1 U997 ( .A1(n1305), .A2(n1306), .ZN(n1296) );
NAND2_X1 U998 ( .A1(n1163), .A2(n1161), .ZN(n1306) );
XOR2_X1 U999 ( .A(KEYINPUT3), .B(n1307), .Z(n1305) );
NOR2_X1 U1000 ( .A1(n1163), .A2(n1161), .ZN(n1307) );
NAND3_X1 U1001 ( .A1(n1260), .A2(n1041), .A3(G210), .ZN(n1161) );
NOR3_X1 U1002 ( .A1(n1065), .A2(n1248), .A3(n1054), .ZN(n1175) );
INV_X1 U1003 ( .A(n1184), .ZN(n1054) );
NOR2_X1 U1004 ( .A1(n1056), .A2(n1057), .ZN(n1184) );
AND2_X1 U1005 ( .A1(G214), .A2(n1308), .ZN(n1057) );
XOR2_X1 U1006 ( .A(n1077), .B(n1309), .Z(n1056) );
NOR2_X1 U1007 ( .A1(KEYINPUT11), .A2(n1078), .ZN(n1309) );
NAND2_X1 U1008 ( .A1(n1310), .A2(n1293), .ZN(n1078) );
XNOR2_X1 U1009 ( .A(n1311), .B(n1207), .ZN(n1310) );
XOR2_X1 U1010 ( .A(n1132), .B(n1312), .Z(n1207) );
NOR2_X1 U1011 ( .A1(KEYINPUT34), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1012 ( .A(n1135), .B(n1314), .Z(n1313) );
NOR2_X1 U1013 ( .A1(n1315), .A2(n1134), .ZN(n1314) );
NAND3_X1 U1014 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1134) );
NAND2_X1 U1015 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1016 ( .A1(n1321), .A2(n1322), .ZN(n1317) );
INV_X1 U1017 ( .A(KEYINPUT20), .ZN(n1322) );
NAND2_X1 U1018 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
INV_X1 U1019 ( .A(n1319), .ZN(n1324) );
XNOR2_X1 U1020 ( .A(KEYINPUT8), .B(n1320), .ZN(n1323) );
NAND2_X1 U1021 ( .A1(KEYINPUT20), .A2(n1325), .ZN(n1316) );
NAND2_X1 U1022 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
OR3_X1 U1023 ( .A1(n1319), .A2(n1320), .A3(KEYINPUT8), .ZN(n1327) );
XNOR2_X1 U1024 ( .A(G104), .B(n1328), .ZN(n1319) );
NAND2_X1 U1025 ( .A1(KEYINPUT8), .A2(n1320), .ZN(n1326) );
XOR2_X1 U1026 ( .A(G101), .B(KEYINPUT47), .Z(n1320) );
XNOR2_X1 U1027 ( .A(KEYINPUT36), .B(KEYINPUT16), .ZN(n1315) );
AND3_X1 U1028 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1135) );
NAND2_X1 U1029 ( .A1(n1332), .A2(n1242), .ZN(n1331) );
INV_X1 U1030 ( .A(G113), .ZN(n1242) );
NAND2_X1 U1031 ( .A1(n1333), .A2(KEYINPUT62), .ZN(n1332) );
XNOR2_X1 U1032 ( .A(n1304), .B(KEYINPUT61), .ZN(n1333) );
NAND3_X1 U1033 ( .A1(KEYINPUT62), .A2(G113), .A3(n1304), .ZN(n1330) );
OR2_X1 U1034 ( .A1(n1304), .A2(KEYINPUT62), .ZN(n1329) );
XOR2_X1 U1035 ( .A(G116), .B(G119), .Z(n1304) );
XNOR2_X1 U1036 ( .A(G110), .B(n1334), .ZN(n1132) );
INV_X1 U1037 ( .A(G122), .ZN(n1334) );
NAND2_X1 U1038 ( .A1(KEYINPUT30), .A2(n1205), .ZN(n1311) );
XNOR2_X1 U1039 ( .A(n1335), .B(n1336), .ZN(n1205) );
XOR2_X1 U1040 ( .A(n1301), .B(n1337), .Z(n1336) );
AND2_X1 U1041 ( .A1(n1041), .A2(G224), .ZN(n1337) );
NOR2_X1 U1042 ( .A1(KEYINPUT33), .A2(n1259), .ZN(n1301) );
XOR2_X1 U1043 ( .A(G143), .B(G146), .Z(n1259) );
XNOR2_X1 U1044 ( .A(G128), .B(G125), .ZN(n1335) );
NAND2_X1 U1045 ( .A1(G210), .A2(n1308), .ZN(n1077) );
NAND2_X1 U1046 ( .A1(n1293), .A2(n1260), .ZN(n1308) );
INV_X1 U1047 ( .A(G237), .ZN(n1260) );
INV_X1 U1048 ( .A(n1230), .ZN(n1248) );
NAND2_X1 U1049 ( .A1(n1069), .A2(n1338), .ZN(n1230) );
NAND4_X1 U1050 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1128), .ZN(n1338) );
INV_X1 U1051 ( .A(G898), .ZN(n1128) );
NAND3_X1 U1052 ( .A1(n1234), .A2(n1041), .A3(G952), .ZN(n1069) );
NAND2_X1 U1053 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U1054 ( .A(n1225), .ZN(n1065) );
NOR2_X1 U1055 ( .A1(n1068), .A2(n1067), .ZN(n1225) );
INV_X1 U1056 ( .A(n1249), .ZN(n1067) );
NAND2_X1 U1057 ( .A1(G221), .A2(n1290), .ZN(n1249) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1293), .ZN(n1290) );
XNOR2_X1 U1059 ( .A(n1339), .B(n1168), .ZN(n1068) );
INV_X1 U1060 ( .A(G469), .ZN(n1168) );
NAND2_X1 U1061 ( .A1(n1340), .A2(n1293), .ZN(n1339) );
INV_X1 U1062 ( .A(G902), .ZN(n1293) );
XNOR2_X1 U1063 ( .A(n1167), .B(n1341), .ZN(n1340) );
XOR2_X1 U1064 ( .A(KEYINPUT9), .B(KEYINPUT39), .Z(n1341) );
XNOR2_X1 U1065 ( .A(n1342), .B(n1343), .ZN(n1167) );
XNOR2_X1 U1066 ( .A(n1163), .B(n1344), .ZN(n1343) );
XNOR2_X1 U1067 ( .A(n1111), .B(G110), .ZN(n1344) );
INV_X1 U1068 ( .A(G140), .ZN(n1111) );
INV_X1 U1069 ( .A(G101), .ZN(n1163) );
XNOR2_X1 U1070 ( .A(n1104), .B(n1345), .ZN(n1342) );
XOR2_X1 U1071 ( .A(n1346), .B(n1347), .Z(n1345) );
NAND2_X1 U1072 ( .A1(G227), .A2(n1041), .ZN(n1347) );
INV_X1 U1073 ( .A(G953), .ZN(n1041) );
NAND2_X1 U1074 ( .A1(n1348), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1075 ( .A1(n1350), .A2(n1253), .ZN(n1349) );
XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n1328), .ZN(n1350) );
XOR2_X1 U1077 ( .A(KEYINPUT44), .B(n1351), .Z(n1348) );
NOR2_X1 U1078 ( .A1(n1253), .A2(n1352), .ZN(n1351) );
XNOR2_X1 U1079 ( .A(KEYINPUT37), .B(n1328), .ZN(n1352) );
INV_X1 U1080 ( .A(G107), .ZN(n1328) );
INV_X1 U1081 ( .A(G104), .ZN(n1253) );
XNOR2_X1 U1082 ( .A(n1300), .B(n1353), .ZN(n1104) );
XOR2_X1 U1083 ( .A(G146), .B(n1354), .Z(n1353) );
NOR2_X1 U1084 ( .A1(G143), .A2(KEYINPUT45), .ZN(n1354) );
XOR2_X1 U1085 ( .A(n1355), .B(n1356), .Z(n1300) );
XOR2_X1 U1086 ( .A(KEYINPUT63), .B(G137), .Z(n1356) );
XNOR2_X1 U1087 ( .A(G131), .B(n1268), .ZN(n1355) );
XOR2_X1 U1088 ( .A(G134), .B(G128), .Z(n1268) );
endmodule


