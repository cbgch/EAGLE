//Key = 1001010101110001100101001110011000000101100000000011011001100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391;

XNOR2_X1 U757 ( .A(G107), .B(n1056), .ZN(G9) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U759 ( .A1(G953), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
XOR2_X1 U760 ( .A(KEYINPUT7), .B(n1062), .Z(n1061) );
NOR3_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR4_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1065) );
NOR2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR3_X1 U769 ( .A1(n1082), .A2(n1083), .A3(n1067), .ZN(n1064) );
XOR2_X1 U770 ( .A(n1084), .B(KEYINPUT41), .Z(n1083) );
NAND2_X1 U771 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U772 ( .A1(n1087), .A2(n1082), .ZN(n1063) );
OR3_X1 U773 ( .A1(n1073), .A2(n1079), .A3(n1069), .ZN(n1082) );
INV_X1 U774 ( .A(n1088), .ZN(n1079) );
INV_X1 U775 ( .A(n1089), .ZN(n1073) );
NOR2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NOR2_X1 U777 ( .A1(n1092), .A2(n1068), .ZN(n1091) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR3_X1 U779 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1057) );
AND4_X1 U780 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1059) );
NOR4_X1 U781 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1098) );
XNOR2_X1 U782 ( .A(G469), .B(n1103), .ZN(n1102) );
XNOR2_X1 U783 ( .A(G472), .B(n1104), .ZN(n1099) );
NOR2_X1 U784 ( .A1(n1105), .A2(KEYINPUT13), .ZN(n1104) );
NOR3_X1 U785 ( .A1(n1106), .A2(n1107), .A3(n1085), .ZN(n1097) );
NAND3_X1 U786 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1096) );
NAND2_X1 U787 ( .A1(KEYINPUT12), .A2(n1111), .ZN(n1110) );
NAND3_X1 U788 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1109) );
INV_X1 U789 ( .A(KEYINPUT12), .ZN(n1113) );
OR2_X1 U790 ( .A1(n1114), .A2(n1112), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1115), .A2(n1111), .ZN(n1112) );
INV_X1 U792 ( .A(KEYINPUT29), .ZN(n1115) );
XNOR2_X1 U793 ( .A(n1116), .B(KEYINPUT25), .ZN(n1114) );
NAND2_X1 U794 ( .A1(G475), .A2(n1117), .ZN(n1095) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(G72) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1120) );
NAND2_X1 U799 ( .A1(n1126), .A2(n1123), .ZN(n1125) );
NAND2_X1 U800 ( .A1(G953), .A2(n1127), .ZN(n1123) );
INV_X1 U801 ( .A(n1128), .ZN(n1126) );
INV_X1 U802 ( .A(n1122), .ZN(n1124) );
XNOR2_X1 U803 ( .A(n1129), .B(n1130), .ZN(n1122) );
NOR2_X1 U804 ( .A1(n1128), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U805 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U806 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NAND3_X1 U807 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(n1138) );
AND2_X1 U809 ( .A1(n1141), .A2(KEYINPUT40), .ZN(n1140) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1143) );
INV_X1 U812 ( .A(KEYINPUT46), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1139), .B(n1144), .Z(n1142) );
NOR2_X1 U814 ( .A1(n1145), .A2(n1141), .ZN(n1144) );
XOR2_X1 U815 ( .A(G134), .B(n1146), .Z(n1141) );
NOR2_X1 U816 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1146) );
INV_X1 U817 ( .A(KEYINPUT40), .ZN(n1145) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1129) );
NAND2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(G69) );
NAND2_X1 U821 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U822 ( .A1(KEYINPUT52), .A2(n1155), .ZN(n1154) );
INV_X1 U823 ( .A(n1156), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1157), .A2(n1156), .ZN(n1153) );
NAND2_X1 U825 ( .A1(n1147), .A2(n1158), .ZN(n1156) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U827 ( .A(n1161), .B(KEYINPUT35), .ZN(n1159) );
NAND2_X1 U828 ( .A1(G953), .A2(n1162), .ZN(n1157) );
NAND2_X1 U829 ( .A1(G898), .A2(G224), .ZN(n1162) );
NAND2_X1 U830 ( .A1(n1163), .A2(n1164), .ZN(n1151) );
NAND2_X1 U831 ( .A1(G953), .A2(n1165), .ZN(n1164) );
XOR2_X1 U832 ( .A(n1166), .B(n1167), .Z(n1163) );
XNOR2_X1 U833 ( .A(n1168), .B(KEYINPUT42), .ZN(n1167) );
NAND2_X1 U834 ( .A1(KEYINPUT16), .A2(n1169), .ZN(n1168) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR4_X1 U836 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(G66) );
NOR2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U838 ( .A(KEYINPUT26), .B(n1178), .Z(n1177) );
NOR2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(n1174) );
XOR2_X1 U840 ( .A(KEYINPUT36), .B(n1178), .Z(n1180) );
NOR2_X1 U841 ( .A1(n1181), .A2(n1116), .ZN(n1178) );
AND2_X1 U842 ( .A1(KEYINPUT24), .A2(n1182), .ZN(n1173) );
NOR3_X1 U843 ( .A1(KEYINPUT24), .A2(G953), .A3(G952), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1182), .A2(n1183), .ZN(G63) );
XNOR2_X1 U845 ( .A(n1184), .B(n1185), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1186), .A2(n1181), .ZN(n1184) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1187), .ZN(G60) );
XOR2_X1 U848 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U849 ( .A1(n1190), .A2(n1181), .ZN(n1189) );
NAND2_X1 U850 ( .A1(n1191), .A2(n1192), .ZN(G6) );
NAND2_X1 U851 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U852 ( .A(KEYINPUT55), .B(n1195), .ZN(n1193) );
NAND2_X1 U853 ( .A1(n1196), .A2(G104), .ZN(n1191) );
XNOR2_X1 U854 ( .A(KEYINPUT58), .B(n1195), .ZN(n1196) );
NOR2_X1 U855 ( .A1(n1182), .A2(n1197), .ZN(G57) );
XOR2_X1 U856 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U857 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U858 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U859 ( .A1(n1204), .A2(n1181), .ZN(n1203) );
NOR2_X1 U860 ( .A1(n1205), .A2(n1206), .ZN(n1202) );
XOR2_X1 U861 ( .A(KEYINPUT17), .B(n1207), .Z(n1206) );
NOR2_X1 U862 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
AND2_X1 U863 ( .A1(n1209), .A2(n1208), .ZN(n1205) );
XOR2_X1 U864 ( .A(n1210), .B(KEYINPUT45), .Z(n1209) );
XOR2_X1 U865 ( .A(n1211), .B(n1212), .Z(n1198) );
XNOR2_X1 U866 ( .A(G101), .B(KEYINPUT47), .ZN(n1212) );
NOR2_X1 U867 ( .A1(n1182), .A2(n1213), .ZN(G54) );
XOR2_X1 U868 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U869 ( .A(n1216), .B(n1217), .Z(n1215) );
NOR2_X1 U870 ( .A1(n1218), .A2(n1181), .ZN(n1217) );
INV_X1 U871 ( .A(G469), .ZN(n1218) );
XNOR2_X1 U872 ( .A(G110), .B(n1219), .ZN(n1214) );
XNOR2_X1 U873 ( .A(KEYINPUT8), .B(n1220), .ZN(n1219) );
NOR3_X1 U874 ( .A1(n1182), .A2(n1221), .A3(n1222), .ZN(G51) );
NOR2_X1 U875 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
INV_X1 U876 ( .A(n1225), .ZN(n1224) );
XOR2_X1 U877 ( .A(KEYINPUT5), .B(n1226), .Z(n1223) );
NOR2_X1 U878 ( .A1(n1225), .A2(n1227), .ZN(n1221) );
XOR2_X1 U879 ( .A(KEYINPUT59), .B(n1226), .Z(n1227) );
XNOR2_X1 U880 ( .A(n1228), .B(n1229), .ZN(n1226) );
NOR3_X1 U881 ( .A1(n1181), .A2(KEYINPUT1), .A3(n1230), .ZN(n1229) );
NAND2_X1 U882 ( .A1(G902), .A2(n1060), .ZN(n1181) );
NAND4_X1 U883 ( .A1(n1149), .A2(n1160), .A3(n1231), .A4(n1232), .ZN(n1060) );
XNOR2_X1 U884 ( .A(KEYINPUT37), .B(n1150), .ZN(n1231) );
AND4_X1 U885 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1160) );
AND4_X1 U886 ( .A1(n1237), .A2(n1056), .A3(n1238), .A4(n1239), .ZN(n1236) );
NAND3_X1 U887 ( .A1(n1090), .A2(n1240), .A3(n1080), .ZN(n1056) );
NOR2_X1 U888 ( .A1(n1241), .A2(n1242), .ZN(n1235) );
NOR2_X1 U889 ( .A1(n1243), .A2(n1195), .ZN(n1242) );
NAND3_X1 U890 ( .A1(n1090), .A2(n1240), .A3(n1081), .ZN(n1195) );
INV_X1 U891 ( .A(KEYINPUT50), .ZN(n1243) );
NOR3_X1 U892 ( .A1(KEYINPUT50), .A2(n1244), .A3(n1245), .ZN(n1241) );
AND3_X1 U893 ( .A1(n1081), .A2(n1246), .A3(n1240), .ZN(n1244) );
INV_X1 U894 ( .A(n1067), .ZN(n1246) );
NAND3_X1 U895 ( .A1(n1089), .A2(n1075), .A3(n1247), .ZN(n1233) );
AND4_X1 U896 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1149) );
NOR3_X1 U897 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
NAND4_X1 U898 ( .A1(n1093), .A2(n1081), .A3(n1255), .A4(n1256), .ZN(n1250) );
NAND2_X1 U899 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
NAND2_X1 U900 ( .A1(n1259), .A2(n1075), .ZN(n1258) );
NAND2_X1 U901 ( .A1(n1088), .A2(n1260), .ZN(n1257) );
NOR2_X1 U902 ( .A1(n1147), .A2(G952), .ZN(n1182) );
XNOR2_X1 U903 ( .A(G146), .B(n1248), .ZN(G48) );
NAND3_X1 U904 ( .A1(n1261), .A2(n1260), .A3(n1081), .ZN(n1248) );
XNOR2_X1 U905 ( .A(G143), .B(n1249), .ZN(G45) );
NAND4_X1 U906 ( .A1(n1262), .A2(n1260), .A3(n1101), .A4(n1263), .ZN(n1249) );
XNOR2_X1 U907 ( .A(G140), .B(n1264), .ZN(G42) );
NAND4_X1 U908 ( .A1(n1265), .A2(n1256), .A3(n1259), .A4(n1266), .ZN(n1264) );
AND2_X1 U909 ( .A1(n1081), .A2(n1093), .ZN(n1266) );
XNOR2_X1 U910 ( .A(KEYINPUT33), .B(n1267), .ZN(n1265) );
NAND2_X1 U911 ( .A1(n1268), .A2(n1269), .ZN(G39) );
NAND2_X1 U912 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
INV_X1 U913 ( .A(n1272), .ZN(n1271) );
NAND2_X1 U914 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U915 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U916 ( .A1(n1252), .A2(n1277), .ZN(n1273) );
NAND2_X1 U917 ( .A1(KEYINPUT10), .A2(n1276), .ZN(n1277) );
INV_X1 U918 ( .A(KEYINPUT4), .ZN(n1276) );
NAND3_X1 U919 ( .A1(KEYINPUT10), .A2(n1252), .A3(n1272), .ZN(n1268) );
XOR2_X1 U920 ( .A(G137), .B(KEYINPUT19), .Z(n1272) );
INV_X1 U921 ( .A(n1275), .ZN(n1252) );
NAND3_X1 U922 ( .A1(n1259), .A2(n1261), .A3(n1089), .ZN(n1275) );
XNOR2_X1 U923 ( .A(G134), .B(n1150), .ZN(G36) );
NAND3_X1 U924 ( .A1(n1259), .A2(n1080), .A3(n1262), .ZN(n1150) );
XNOR2_X1 U925 ( .A(n1136), .B(n1254), .ZN(G33) );
AND3_X1 U926 ( .A1(n1262), .A2(n1259), .A3(n1081), .ZN(n1254) );
INV_X1 U927 ( .A(n1068), .ZN(n1259) );
NAND2_X1 U928 ( .A1(n1086), .A2(n1278), .ZN(n1068) );
AND3_X1 U929 ( .A1(n1075), .A2(n1256), .A3(n1094), .ZN(n1262) );
XOR2_X1 U930 ( .A(G128), .B(n1253), .Z(G30) );
AND3_X1 U931 ( .A1(n1080), .A2(n1260), .A3(n1261), .ZN(n1253) );
NOR4_X1 U932 ( .A1(n1267), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1261) );
INV_X1 U933 ( .A(n1256), .ZN(n1281) );
XNOR2_X1 U934 ( .A(G101), .B(n1282), .ZN(G3) );
NAND3_X1 U935 ( .A1(n1247), .A2(n1089), .A3(n1283), .ZN(n1282) );
XNOR2_X1 U936 ( .A(n1075), .B(KEYINPUT21), .ZN(n1283) );
INV_X1 U937 ( .A(n1267), .ZN(n1075) );
XNOR2_X1 U938 ( .A(G125), .B(n1284), .ZN(G27) );
NAND4_X1 U939 ( .A1(n1093), .A2(n1081), .A3(n1285), .A4(n1088), .ZN(n1284) );
NOR2_X1 U940 ( .A1(n1286), .A2(n1245), .ZN(n1285) );
XOR2_X1 U941 ( .A(n1256), .B(KEYINPUT11), .Z(n1286) );
NAND2_X1 U942 ( .A1(n1069), .A2(n1287), .ZN(n1256) );
NAND3_X1 U943 ( .A1(G902), .A2(n1288), .A3(n1128), .ZN(n1287) );
NOR2_X1 U944 ( .A1(G900), .A2(n1147), .ZN(n1128) );
XNOR2_X1 U945 ( .A(G122), .B(n1289), .ZN(G24) );
NOR2_X1 U946 ( .A1(n1161), .A2(KEYINPUT49), .ZN(n1289) );
INV_X1 U947 ( .A(n1232), .ZN(n1161) );
NAND3_X1 U948 ( .A1(n1088), .A2(n1090), .A3(n1290), .ZN(n1232) );
NOR3_X1 U949 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1290) );
NOR2_X1 U950 ( .A1(n1245), .A2(n1067), .ZN(n1090) );
NAND2_X1 U951 ( .A1(n1294), .A2(n1280), .ZN(n1067) );
INV_X1 U952 ( .A(n1260), .ZN(n1245) );
XNOR2_X1 U953 ( .A(n1295), .B(n1237), .ZN(G21) );
NAND4_X1 U954 ( .A1(n1088), .A2(n1260), .A3(n1089), .A4(n1296), .ZN(n1237) );
NOR3_X1 U955 ( .A1(n1279), .A2(n1293), .A3(n1280), .ZN(n1296) );
INV_X1 U956 ( .A(n1297), .ZN(n1280) );
NAND2_X1 U957 ( .A1(KEYINPUT62), .A2(n1298), .ZN(n1295) );
XNOR2_X1 U958 ( .A(G116), .B(n1239), .ZN(G18) );
NAND3_X1 U959 ( .A1(n1088), .A2(n1080), .A3(n1247), .ZN(n1239) );
NOR2_X1 U960 ( .A1(n1263), .A2(n1291), .ZN(n1080) );
INV_X1 U961 ( .A(n1101), .ZN(n1291) );
XNOR2_X1 U962 ( .A(G113), .B(n1238), .ZN(G15) );
NAND3_X1 U963 ( .A1(n1081), .A2(n1088), .A3(n1247), .ZN(n1238) );
AND3_X1 U964 ( .A1(n1260), .A2(n1299), .A3(n1094), .ZN(n1247) );
AND2_X1 U965 ( .A1(n1294), .A2(n1297), .ZN(n1094) );
NOR2_X1 U966 ( .A1(n1076), .A2(n1106), .ZN(n1088) );
INV_X1 U967 ( .A(n1077), .ZN(n1106) );
NOR2_X1 U968 ( .A1(n1101), .A2(n1292), .ZN(n1081) );
INV_X1 U969 ( .A(n1263), .ZN(n1292) );
XNOR2_X1 U970 ( .A(G110), .B(n1234), .ZN(G12) );
NAND4_X1 U971 ( .A1(n1093), .A2(n1089), .A3(n1240), .A4(n1260), .ZN(n1234) );
NOR2_X1 U972 ( .A1(n1086), .A2(n1085), .ZN(n1260) );
INV_X1 U973 ( .A(n1278), .ZN(n1085) );
NAND2_X1 U974 ( .A1(G214), .A2(n1300), .ZN(n1278) );
XOR2_X1 U975 ( .A(n1100), .B(KEYINPUT9), .Z(n1086) );
XOR2_X1 U976 ( .A(n1301), .B(n1230), .Z(n1100) );
NAND2_X1 U977 ( .A1(G210), .A2(n1300), .ZN(n1230) );
NAND2_X1 U978 ( .A1(n1302), .A2(n1119), .ZN(n1300) );
NAND2_X1 U979 ( .A1(n1303), .A2(n1119), .ZN(n1301) );
XNOR2_X1 U980 ( .A(n1225), .B(n1304), .ZN(n1303) );
XNOR2_X1 U981 ( .A(KEYINPUT51), .B(n1228), .ZN(n1304) );
XOR2_X1 U982 ( .A(n1166), .B(n1305), .Z(n1228) );
NOR2_X1 U983 ( .A1(KEYINPUT32), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U984 ( .A(n1170), .B(n1171), .ZN(n1306) );
XOR2_X1 U985 ( .A(n1307), .B(n1308), .Z(n1171) );
NOR2_X1 U986 ( .A1(G101), .A2(KEYINPUT22), .ZN(n1308) );
XOR2_X1 U987 ( .A(G104), .B(n1309), .Z(n1170) );
XNOR2_X1 U988 ( .A(n1310), .B(G107), .ZN(n1309) );
XOR2_X1 U989 ( .A(n1311), .B(G122), .Z(n1166) );
NAND2_X1 U990 ( .A1(KEYINPUT63), .A2(n1312), .ZN(n1311) );
XOR2_X1 U991 ( .A(n1313), .B(n1314), .Z(n1225) );
INV_X1 U992 ( .A(n1210), .ZN(n1314) );
XNOR2_X1 U993 ( .A(G125), .B(n1315), .ZN(n1313) );
AND2_X1 U994 ( .A1(n1147), .A2(G224), .ZN(n1315) );
NOR2_X1 U995 ( .A1(n1267), .A2(n1293), .ZN(n1240) );
INV_X1 U996 ( .A(n1299), .ZN(n1293) );
NAND2_X1 U997 ( .A1(n1069), .A2(n1316), .ZN(n1299) );
NAND4_X1 U998 ( .A1(G953), .A2(G902), .A3(n1288), .A4(n1165), .ZN(n1316) );
INV_X1 U999 ( .A(G898), .ZN(n1165) );
NAND3_X1 U1000 ( .A1(n1288), .A2(n1147), .A3(G952), .ZN(n1069) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1288) );
NAND2_X1 U1002 ( .A1(n1077), .A2(n1076), .ZN(n1267) );
NAND2_X1 U1003 ( .A1(n1317), .A2(n1318), .ZN(n1076) );
NAND2_X1 U1004 ( .A1(n1319), .A2(n1103), .ZN(n1318) );
XOR2_X1 U1005 ( .A(n1320), .B(KEYINPUT6), .Z(n1317) );
OR2_X1 U1006 ( .A1(n1103), .A2(n1319), .ZN(n1320) );
XOR2_X1 U1007 ( .A(G469), .B(KEYINPUT2), .Z(n1319) );
NAND2_X1 U1008 ( .A1(n1321), .A2(n1119), .ZN(n1103) );
XOR2_X1 U1009 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1010 ( .A(n1324), .B(n1216), .Z(n1323) );
XOR2_X1 U1011 ( .A(n1325), .B(n1326), .Z(n1216) );
XOR2_X1 U1012 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1013 ( .A(G101), .B(n1329), .Z(n1328) );
NOR2_X1 U1014 ( .A1(G953), .A2(n1127), .ZN(n1329) );
INV_X1 U1015 ( .A(G227), .ZN(n1127) );
XOR2_X1 U1016 ( .A(KEYINPUT20), .B(G107), .Z(n1327) );
XNOR2_X1 U1017 ( .A(n1330), .B(n1331), .ZN(n1325) );
XOR2_X1 U1018 ( .A(n1139), .B(n1332), .Z(n1330) );
NOR2_X1 U1019 ( .A1(KEYINPUT27), .A2(n1194), .ZN(n1332) );
XOR2_X1 U1020 ( .A(n1333), .B(G128), .Z(n1139) );
NAND2_X1 U1021 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1022 ( .A1(G143), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1023 ( .A(KEYINPUT39), .B(n1337), .Z(n1334) );
NOR2_X1 U1024 ( .A1(G143), .A2(n1336), .ZN(n1337) );
NAND2_X1 U1025 ( .A1(KEYINPUT53), .A2(n1220), .ZN(n1324) );
XNOR2_X1 U1026 ( .A(KEYINPUT14), .B(n1312), .ZN(n1322) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1338), .ZN(n1077) );
NOR2_X1 U1028 ( .A1(n1101), .A2(n1263), .ZN(n1089) );
NAND2_X1 U1029 ( .A1(n1339), .A2(n1340), .ZN(n1263) );
NAND2_X1 U1030 ( .A1(G475), .A2(n1341), .ZN(n1340) );
NAND3_X1 U1031 ( .A1(n1118), .A2(n1119), .A3(KEYINPUT15), .ZN(n1341) );
NAND2_X1 U1032 ( .A1(n1107), .A2(KEYINPUT15), .ZN(n1339) );
AND3_X1 U1033 ( .A1(n1190), .A2(n1119), .A3(n1118), .ZN(n1107) );
XNOR2_X1 U1034 ( .A(n1188), .B(KEYINPUT38), .ZN(n1118) );
XOR2_X1 U1035 ( .A(n1342), .B(n1343), .Z(n1188) );
XNOR2_X1 U1036 ( .A(n1310), .B(n1344), .ZN(n1343) );
XNOR2_X1 U1037 ( .A(n1136), .B(G122), .ZN(n1344) );
XNOR2_X1 U1038 ( .A(n1345), .B(n1346), .ZN(n1342) );
XOR2_X1 U1039 ( .A(n1347), .B(n1348), .Z(n1346) );
NOR2_X1 U1040 ( .A1(KEYINPUT34), .A2(n1194), .ZN(n1348) );
INV_X1 U1041 ( .A(G104), .ZN(n1194) );
NOR2_X1 U1042 ( .A1(n1349), .A2(n1350), .ZN(n1347) );
XOR2_X1 U1043 ( .A(n1351), .B(KEYINPUT57), .Z(n1350) );
NAND2_X1 U1044 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND3_X1 U1045 ( .A1(n1302), .A2(n1147), .A3(G214), .ZN(n1353) );
XOR2_X1 U1046 ( .A(KEYINPUT54), .B(G143), .Z(n1352) );
AND4_X1 U1047 ( .A1(n1147), .A2(n1302), .A3(G143), .A4(G214), .ZN(n1349) );
INV_X1 U1048 ( .A(G475), .ZN(n1190) );
XOR2_X1 U1049 ( .A(n1354), .B(n1186), .Z(n1101) );
INV_X1 U1050 ( .A(G478), .ZN(n1186) );
NAND2_X1 U1051 ( .A1(n1355), .A2(n1185), .ZN(n1354) );
XOR2_X1 U1052 ( .A(n1356), .B(n1357), .Z(n1185) );
XOR2_X1 U1053 ( .A(G107), .B(n1358), .Z(n1357) );
XNOR2_X1 U1054 ( .A(n1359), .B(G122), .ZN(n1358) );
XOR2_X1 U1055 ( .A(n1360), .B(n1361), .Z(n1356) );
XOR2_X1 U1056 ( .A(n1362), .B(n1363), .Z(n1360) );
NOR2_X1 U1057 ( .A1(KEYINPUT28), .A2(G116), .ZN(n1363) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1364), .ZN(n1362) );
XNOR2_X1 U1059 ( .A(G902), .B(KEYINPUT48), .ZN(n1355) );
NOR2_X1 U1060 ( .A1(n1297), .A2(n1279), .ZN(n1093) );
XOR2_X1 U1061 ( .A(n1294), .B(KEYINPUT43), .Z(n1279) );
XOR2_X1 U1062 ( .A(n1111), .B(n1116), .Z(n1294) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1338), .ZN(n1116) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1119), .ZN(n1338) );
NOR2_X1 U1065 ( .A1(n1176), .A2(G902), .ZN(n1111) );
INV_X1 U1066 ( .A(n1179), .ZN(n1176) );
XNOR2_X1 U1067 ( .A(n1365), .B(n1366), .ZN(n1179) );
XNOR2_X1 U1068 ( .A(n1298), .B(n1367), .ZN(n1366) );
XNOR2_X1 U1069 ( .A(n1368), .B(G128), .ZN(n1367) );
XOR2_X1 U1070 ( .A(n1369), .B(n1345), .Z(n1365) );
XOR2_X1 U1071 ( .A(G146), .B(n1133), .Z(n1345) );
XNOR2_X1 U1072 ( .A(G125), .B(n1220), .ZN(n1133) );
INV_X1 U1073 ( .A(G140), .ZN(n1220) );
XNOR2_X1 U1074 ( .A(n1370), .B(n1312), .ZN(n1369) );
INV_X1 U1075 ( .A(G110), .ZN(n1312) );
NAND2_X1 U1076 ( .A1(G221), .A2(n1364), .ZN(n1370) );
AND2_X1 U1077 ( .A1(G234), .A2(n1147), .ZN(n1364) );
XNOR2_X1 U1078 ( .A(n1371), .B(n1372), .ZN(n1297) );
NOR2_X1 U1079 ( .A1(KEYINPUT44), .A2(n1204), .ZN(n1372) );
INV_X1 U1080 ( .A(G472), .ZN(n1204) );
XNOR2_X1 U1081 ( .A(n1105), .B(KEYINPUT60), .ZN(n1371) );
AND2_X1 U1082 ( .A1(n1373), .A2(n1119), .ZN(n1105) );
INV_X1 U1083 ( .A(G902), .ZN(n1119) );
XOR2_X1 U1084 ( .A(n1374), .B(n1375), .Z(n1373) );
XNOR2_X1 U1085 ( .A(n1376), .B(n1211), .ZN(n1375) );
NAND3_X1 U1086 ( .A1(n1302), .A2(n1147), .A3(G210), .ZN(n1211) );
INV_X1 U1087 ( .A(G953), .ZN(n1147) );
INV_X1 U1088 ( .A(G237), .ZN(n1302) );
NOR2_X1 U1089 ( .A1(KEYINPUT18), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1090 ( .A(n1378), .B(n1379), .Z(n1377) );
XOR2_X1 U1091 ( .A(KEYINPUT61), .B(n1200), .Z(n1379) );
XNOR2_X1 U1092 ( .A(n1380), .B(n1307), .ZN(n1200) );
XNOR2_X1 U1093 ( .A(G116), .B(n1298), .ZN(n1307) );
INV_X1 U1094 ( .A(G119), .ZN(n1298) );
NAND2_X1 U1095 ( .A1(KEYINPUT30), .A2(n1310), .ZN(n1380) );
INV_X1 U1096 ( .A(G113), .ZN(n1310) );
XNOR2_X1 U1097 ( .A(n1208), .B(n1210), .ZN(n1378) );
XOR2_X1 U1098 ( .A(n1361), .B(n1381), .Z(n1210) );
NOR2_X1 U1099 ( .A1(KEYINPUT31), .A2(n1336), .ZN(n1381) );
INV_X1 U1100 ( .A(G146), .ZN(n1336) );
XOR2_X1 U1101 ( .A(G128), .B(G143), .Z(n1361) );
INV_X1 U1102 ( .A(n1331), .ZN(n1208) );
NAND2_X1 U1103 ( .A1(n1382), .A2(n1383), .ZN(n1331) );
NAND2_X1 U1104 ( .A1(n1384), .A2(n1368), .ZN(n1383) );
INV_X1 U1105 ( .A(G137), .ZN(n1368) );
NAND2_X1 U1106 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
NAND2_X1 U1107 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XNOR2_X1 U1108 ( .A(KEYINPUT23), .B(n1359), .ZN(n1388) );
XNOR2_X1 U1109 ( .A(KEYINPUT0), .B(G131), .ZN(n1387) );
NAND2_X1 U1110 ( .A1(n1389), .A2(n1136), .ZN(n1385) );
INV_X1 U1111 ( .A(G131), .ZN(n1136) );
XNOR2_X1 U1112 ( .A(KEYINPUT23), .B(G134), .ZN(n1389) );
NAND2_X1 U1113 ( .A1(G137), .A2(n1390), .ZN(n1382) );
XNOR2_X1 U1114 ( .A(G131), .B(n1391), .ZN(n1390) );
AND2_X1 U1115 ( .A1(n1359), .A2(KEYINPUT0), .ZN(n1391) );
INV_X1 U1116 ( .A(G134), .ZN(n1359) );
NAND2_X1 U1117 ( .A1(KEYINPUT3), .A2(G101), .ZN(n1374) );
endmodule


