//Key = 0100010000011001000110000011011100001100111111010001100011110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321;

XNOR2_X1 U724 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U725 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR4_X1 U726 ( .A1(n1017), .A2(n1018), .A3(G953), .A4(n1019), .ZN(n1016) );
NAND3_X1 U727 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1017) );
NAND2_X1 U728 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NAND2_X1 U729 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND3_X1 U730 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NAND2_X1 U731 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NAND2_X1 U732 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U733 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U734 ( .A1(n1036), .A2(n1037), .ZN(n1030) );
NAND2_X1 U735 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U736 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND3_X1 U737 ( .A1(n1032), .A2(n1042), .A3(n1036), .ZN(n1025) );
NAND2_X1 U738 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U739 ( .A1(n1029), .A2(n1045), .ZN(n1044) );
NAND2_X1 U740 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U741 ( .A1(n1027), .A2(n1048), .ZN(n1043) );
NAND2_X1 U742 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U743 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U744 ( .A(n1053), .ZN(n1032) );
INV_X1 U745 ( .A(n1054), .ZN(n1023) );
NOR3_X1 U746 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n1015) );
AND4_X1 U747 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1019) );
NOR3_X1 U748 ( .A1(n1059), .A2(n1053), .A3(n1060), .ZN(n1058) );
XNOR2_X1 U749 ( .A(KEYINPUT3), .B(n1061), .ZN(n1059) );
XOR2_X1 U750 ( .A(n1062), .B(n1063), .Z(n1055) );
NAND2_X1 U751 ( .A1(KEYINPUT29), .A2(n1064), .ZN(n1063) );
XOR2_X1 U752 ( .A(n1065), .B(n1066), .Z(G72) );
NOR2_X1 U753 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U754 ( .A1(G227), .A2(G900), .ZN(n1067) );
NOR2_X1 U755 ( .A1(KEYINPUT16), .A2(n1069), .ZN(n1065) );
XOR2_X1 U756 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U757 ( .A1(KEYINPUT41), .A2(n1072), .ZN(n1071) );
NAND2_X1 U758 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U759 ( .A1(n1075), .A2(G953), .ZN(n1074) );
XNOR2_X1 U760 ( .A(G900), .B(KEYINPUT17), .ZN(n1075) );
XOR2_X1 U761 ( .A(n1076), .B(n1077), .Z(n1073) );
XOR2_X1 U762 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U763 ( .A1(G140), .A2(KEYINPUT7), .ZN(n1078) );
XOR2_X1 U764 ( .A(n1080), .B(n1081), .Z(n1076) );
XNOR2_X1 U765 ( .A(G125), .B(n1082), .ZN(n1081) );
NAND2_X1 U766 ( .A1(KEYINPUT52), .A2(n1083), .ZN(n1080) );
NAND2_X1 U767 ( .A1(n1068), .A2(n1084), .ZN(n1070) );
NAND2_X1 U768 ( .A1(n1085), .A2(n1022), .ZN(n1084) );
XNOR2_X1 U769 ( .A(n1018), .B(KEYINPUT9), .ZN(n1085) );
NAND2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(G69) );
NAND2_X1 U771 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U772 ( .A(KEYINPUT30), .B(n1090), .Z(n1086) );
NOR2_X1 U773 ( .A1(n1088), .A2(n1089), .ZN(n1090) );
NAND2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
OR2_X1 U775 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U776 ( .A(n1095), .B(KEYINPUT34), .Z(n1091) );
NAND2_X1 U777 ( .A1(n1094), .A2(n1093), .ZN(n1095) );
NAND2_X1 U778 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND2_X1 U779 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XOR2_X1 U780 ( .A(n1099), .B(n1100), .Z(n1096) );
XOR2_X1 U781 ( .A(n1101), .B(n1102), .Z(n1099) );
NOR2_X1 U782 ( .A1(KEYINPUT50), .A2(n1103), .ZN(n1102) );
NOR2_X1 U783 ( .A1(G953), .A2(n1020), .ZN(n1094) );
NAND2_X1 U784 ( .A1(G953), .A2(n1104), .ZN(n1088) );
NAND2_X1 U785 ( .A1(G898), .A2(G224), .ZN(n1104) );
NOR2_X1 U786 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U787 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U789 ( .A1(n1111), .A2(KEYINPUT58), .ZN(n1107) );
XNOR2_X1 U790 ( .A(n1112), .B(n1113), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1114), .ZN(G63) );
XNOR2_X1 U792 ( .A(n1115), .B(n1116), .ZN(n1114) );
AND2_X1 U793 ( .A1(G478), .A2(n1109), .ZN(n1116) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1117), .ZN(G60) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U796 ( .A1(KEYINPUT10), .A2(n1120), .ZN(n1119) );
NAND2_X1 U797 ( .A1(n1109), .A2(G475), .ZN(n1118) );
NAND3_X1 U798 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(G6) );
OR2_X1 U799 ( .A1(n1124), .A2(KEYINPUT56), .ZN(n1123) );
NAND3_X1 U800 ( .A1(KEYINPUT56), .A2(n1124), .A3(n1125), .ZN(n1122) );
NAND2_X1 U801 ( .A1(G104), .A2(n1126), .ZN(n1121) );
NAND2_X1 U802 ( .A1(n1127), .A2(KEYINPUT56), .ZN(n1126) );
XNOR2_X1 U803 ( .A(n1124), .B(KEYINPUT59), .ZN(n1127) );
INV_X1 U804 ( .A(n1128), .ZN(n1124) );
NOR2_X1 U805 ( .A1(n1105), .A2(n1129), .ZN(G57) );
XOR2_X1 U806 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U807 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U808 ( .A1(KEYINPUT26), .A2(n1134), .ZN(n1132) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(n1130) );
XOR2_X1 U810 ( .A(G101), .B(n1137), .Z(n1136) );
AND2_X1 U811 ( .A1(G472), .A2(n1109), .ZN(n1137) );
NAND2_X1 U812 ( .A1(KEYINPUT19), .A2(n1138), .ZN(n1135) );
XNOR2_X1 U813 ( .A(KEYINPUT57), .B(n1139), .ZN(n1138) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(G54) );
XOR2_X1 U815 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U816 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U817 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U818 ( .A(n1148), .B(n1149), .Z(n1142) );
XNOR2_X1 U819 ( .A(KEYINPUT55), .B(n1082), .ZN(n1149) );
AND2_X1 U820 ( .A1(G469), .A2(n1109), .ZN(n1148) );
INV_X1 U821 ( .A(n1150), .ZN(n1109) );
XOR2_X1 U822 ( .A(n1151), .B(KEYINPUT20), .Z(n1140) );
NAND2_X1 U823 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U824 ( .A(KEYINPUT51), .B(G952), .Z(n1153) );
XNOR2_X1 U825 ( .A(KEYINPUT60), .B(n1068), .ZN(n1152) );
NOR2_X1 U826 ( .A1(n1105), .A2(n1154), .ZN(G51) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U828 ( .A1(n1064), .A2(n1150), .ZN(n1156) );
NAND2_X1 U829 ( .A1(G902), .A2(n1157), .ZN(n1150) );
NAND3_X1 U830 ( .A1(n1020), .A2(n1158), .A3(n1022), .ZN(n1157) );
AND4_X1 U831 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1022) );
AND4_X1 U832 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
AND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1020) );
AND4_X1 U834 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1128), .ZN(n1168) );
NAND3_X1 U835 ( .A1(n1027), .A2(n1172), .A3(n1173), .ZN(n1128) );
NOR4_X1 U836 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1167) );
INV_X1 U837 ( .A(n1178), .ZN(n1177) );
NOR4_X1 U838 ( .A1(n1179), .A2(n1180), .A3(n1035), .A4(n1046), .ZN(n1176) );
INV_X1 U839 ( .A(n1181), .ZN(n1046) );
NOR2_X1 U840 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
INV_X1 U841 ( .A(KEYINPUT0), .ZN(n1183) );
NOR3_X1 U842 ( .A1(n1053), .A2(n1184), .A3(n1185), .ZN(n1182) );
NOR2_X1 U843 ( .A1(KEYINPUT0), .A2(n1186), .ZN(n1179) );
INV_X1 U844 ( .A(n1014), .ZN(n1175) );
NAND3_X1 U845 ( .A1(n1027), .A2(n1172), .A3(n1187), .ZN(n1014) );
NOR3_X1 U846 ( .A1(n1188), .A2(n1047), .A3(n1189), .ZN(n1174) );
XNOR2_X1 U847 ( .A(KEYINPUT40), .B(n1038), .ZN(n1189) );
INV_X1 U848 ( .A(n1190), .ZN(n1047) );
NAND3_X1 U849 ( .A1(n1191), .A2(n1192), .A3(n1036), .ZN(n1188) );
XNOR2_X1 U850 ( .A(KEYINPUT24), .B(n1049), .ZN(n1191) );
NOR2_X1 U851 ( .A1(KEYINPUT18), .A2(n1193), .ZN(n1155) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U853 ( .A1(KEYINPUT28), .A2(n1196), .ZN(n1195) );
NOR2_X1 U854 ( .A1(n1197), .A2(G952), .ZN(n1105) );
XNOR2_X1 U855 ( .A(KEYINPUT60), .B(G953), .ZN(n1197) );
XNOR2_X1 U856 ( .A(G146), .B(n1161), .ZN(G48) );
NAND3_X1 U857 ( .A1(n1173), .A2(n1184), .A3(n1198), .ZN(n1161) );
XNOR2_X1 U858 ( .A(n1018), .B(n1199), .ZN(G45) );
NAND2_X1 U859 ( .A1(KEYINPUT12), .A2(G143), .ZN(n1199) );
INV_X1 U860 ( .A(n1158), .ZN(n1018) );
NAND4_X1 U861 ( .A1(n1200), .A2(n1181), .A3(n1201), .A4(n1184), .ZN(n1158) );
XNOR2_X1 U862 ( .A(G140), .B(n1159), .ZN(G42) );
NAND4_X1 U863 ( .A1(n1029), .A2(n1201), .A3(n1190), .A4(n1173), .ZN(n1159) );
XNOR2_X1 U864 ( .A(G137), .B(n1160), .ZN(G39) );
NAND3_X1 U865 ( .A1(n1198), .A2(n1036), .A3(n1029), .ZN(n1160) );
XNOR2_X1 U866 ( .A(G134), .B(n1166), .ZN(G36) );
NAND2_X1 U867 ( .A1(n1202), .A2(n1187), .ZN(n1166) );
XNOR2_X1 U868 ( .A(G131), .B(n1165), .ZN(G33) );
NAND2_X1 U869 ( .A1(n1202), .A2(n1173), .ZN(n1165) );
AND3_X1 U870 ( .A1(n1029), .A2(n1201), .A3(n1181), .ZN(n1202) );
NOR2_X1 U871 ( .A1(n1203), .A2(n1051), .ZN(n1029) );
XNOR2_X1 U872 ( .A(G128), .B(n1164), .ZN(G30) );
NAND3_X1 U873 ( .A1(n1187), .A2(n1184), .A3(n1198), .ZN(n1164) );
AND3_X1 U874 ( .A1(n1204), .A2(n1205), .A3(n1201), .ZN(n1198) );
NOR2_X1 U875 ( .A1(n1038), .A2(n1206), .ZN(n1201) );
XOR2_X1 U876 ( .A(n1171), .B(n1207), .Z(G3) );
NOR2_X1 U877 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1207) );
NAND3_X1 U878 ( .A1(n1036), .A2(n1172), .A3(n1181), .ZN(n1171) );
XNOR2_X1 U879 ( .A(G125), .B(n1163), .ZN(G27) );
NAND3_X1 U880 ( .A1(n1190), .A2(n1173), .A3(n1208), .ZN(n1163) );
NOR3_X1 U881 ( .A1(n1053), .A2(n1206), .A3(n1049), .ZN(n1208) );
AND2_X1 U882 ( .A1(n1054), .A2(n1209), .ZN(n1206) );
NAND4_X1 U883 ( .A1(G953), .A2(G902), .A3(n1210), .A4(n1211), .ZN(n1209) );
INV_X1 U884 ( .A(G900), .ZN(n1211) );
XNOR2_X1 U885 ( .A(G122), .B(n1178), .ZN(G24) );
NAND3_X1 U886 ( .A1(n1186), .A2(n1027), .A3(n1200), .ZN(n1178) );
AND2_X1 U887 ( .A1(n1212), .A2(n1213), .ZN(n1200) );
XNOR2_X1 U888 ( .A(KEYINPUT48), .B(n1214), .ZN(n1212) );
NOR2_X1 U889 ( .A1(n1205), .A2(n1204), .ZN(n1027) );
XOR2_X1 U890 ( .A(n1170), .B(n1215), .Z(G21) );
XNOR2_X1 U891 ( .A(KEYINPUT31), .B(n1216), .ZN(n1215) );
NAND4_X1 U892 ( .A1(n1186), .A2(n1036), .A3(n1204), .A4(n1205), .ZN(n1170) );
NAND2_X1 U893 ( .A1(n1217), .A2(n1218), .ZN(G18) );
NAND2_X1 U894 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U895 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
OR2_X1 U896 ( .A1(n1223), .A2(KEYINPUT33), .ZN(n1222) );
NAND2_X1 U897 ( .A1(n1224), .A2(n1223), .ZN(n1221) );
OR2_X1 U898 ( .A1(KEYINPUT33), .A2(KEYINPUT62), .ZN(n1224) );
NAND3_X1 U899 ( .A1(n1223), .A2(n1225), .A3(G116), .ZN(n1217) );
INV_X1 U900 ( .A(KEYINPUT62), .ZN(n1225) );
NAND3_X1 U901 ( .A1(n1181), .A2(n1187), .A3(n1186), .ZN(n1223) );
INV_X1 U902 ( .A(n1035), .ZN(n1187) );
NAND2_X1 U903 ( .A1(n1214), .A2(n1213), .ZN(n1035) );
XNOR2_X1 U904 ( .A(n1226), .B(KEYINPUT49), .ZN(n1213) );
XNOR2_X1 U905 ( .A(G113), .B(n1169), .ZN(G15) );
NAND3_X1 U906 ( .A1(n1181), .A2(n1173), .A3(n1186), .ZN(n1169) );
NOR3_X1 U907 ( .A1(n1049), .A2(n1185), .A3(n1053), .ZN(n1186) );
NAND2_X1 U908 ( .A1(n1041), .A2(n1227), .ZN(n1053) );
INV_X1 U909 ( .A(n1034), .ZN(n1173) );
NAND2_X1 U910 ( .A1(n1226), .A2(n1228), .ZN(n1034) );
NOR2_X1 U911 ( .A1(n1204), .A2(n1057), .ZN(n1181) );
INV_X1 U912 ( .A(n1205), .ZN(n1057) );
XOR2_X1 U913 ( .A(n1229), .B(n1230), .Z(G12) );
AND3_X1 U914 ( .A1(n1190), .A2(n1172), .A3(n1036), .ZN(n1230) );
INV_X1 U915 ( .A(n1060), .ZN(n1036) );
NAND2_X1 U916 ( .A1(n1214), .A2(n1226), .ZN(n1060) );
XOR2_X1 U917 ( .A(n1231), .B(G478), .Z(n1226) );
NAND2_X1 U918 ( .A1(n1115), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U919 ( .A(n1233), .B(n1234), .ZN(n1115) );
XOR2_X1 U920 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U921 ( .A(G128), .B(n1237), .ZN(n1236) );
INV_X1 U922 ( .A(G122), .ZN(n1237) );
XOR2_X1 U923 ( .A(G143), .B(G134), .Z(n1235) );
XOR2_X1 U924 ( .A(n1238), .B(n1239), .Z(n1233) );
XNOR2_X1 U925 ( .A(n1220), .B(G107), .ZN(n1239) );
INV_X1 U926 ( .A(G116), .ZN(n1220) );
NAND2_X1 U927 ( .A1(G217), .A2(n1240), .ZN(n1238) );
INV_X1 U928 ( .A(n1228), .ZN(n1214) );
XNOR2_X1 U929 ( .A(n1241), .B(G475), .ZN(n1228) );
OR2_X1 U930 ( .A1(n1120), .A2(G902), .ZN(n1241) );
XNOR2_X1 U931 ( .A(G122), .B(n1242), .ZN(n1120) );
XOR2_X1 U932 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U933 ( .A(n1245), .B(n1246), .Z(n1244) );
XNOR2_X1 U934 ( .A(n1247), .B(n1248), .ZN(n1246) );
NOR4_X1 U935 ( .A1(KEYINPUT2), .A2(G953), .A3(G237), .A4(n1249), .ZN(n1248) );
INV_X1 U936 ( .A(G214), .ZN(n1249) );
XNOR2_X1 U937 ( .A(n1250), .B(n1251), .ZN(n1245) );
NAND2_X1 U938 ( .A1(KEYINPUT43), .A2(n1252), .ZN(n1251) );
INV_X1 U939 ( .A(G113), .ZN(n1252) );
NAND2_X1 U940 ( .A1(KEYINPUT1), .A2(n1253), .ZN(n1250) );
XOR2_X1 U941 ( .A(n1254), .B(n1255), .Z(n1243) );
XNOR2_X1 U942 ( .A(n1083), .B(G104), .ZN(n1255) );
INV_X1 U943 ( .A(G131), .ZN(n1083) );
XOR2_X1 U944 ( .A(KEYINPUT4), .B(KEYINPUT11), .Z(n1254) );
NOR3_X1 U945 ( .A1(n1049), .A2(n1185), .A3(n1038), .ZN(n1172) );
OR2_X1 U946 ( .A1(n1041), .A2(n1040), .ZN(n1038) );
INV_X1 U947 ( .A(n1227), .ZN(n1040) );
NAND2_X1 U948 ( .A1(G221), .A2(n1256), .ZN(n1227) );
XOR2_X1 U949 ( .A(n1257), .B(G469), .Z(n1041) );
NAND2_X1 U950 ( .A1(n1258), .A2(n1232), .ZN(n1257) );
XOR2_X1 U951 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U952 ( .A(n1147), .B(n1144), .Z(n1260) );
XOR2_X1 U953 ( .A(n1261), .B(KEYINPUT61), .Z(n1144) );
XNOR2_X1 U954 ( .A(n1262), .B(n1263), .ZN(n1147) );
XOR2_X1 U955 ( .A(G140), .B(G110), .Z(n1263) );
NAND2_X1 U956 ( .A1(G227), .A2(n1068), .ZN(n1262) );
XNOR2_X1 U957 ( .A(n1264), .B(n1082), .ZN(n1259) );
NAND2_X1 U958 ( .A1(n1265), .A2(n1266), .ZN(n1082) );
NAND2_X1 U959 ( .A1(G128), .A2(n1247), .ZN(n1266) );
XOR2_X1 U960 ( .A(KEYINPUT63), .B(n1267), .Z(n1265) );
NOR2_X1 U961 ( .A1(G128), .A2(n1247), .ZN(n1267) );
XNOR2_X1 U962 ( .A(KEYINPUT25), .B(n1268), .ZN(n1264) );
NOR2_X1 U963 ( .A1(KEYINPUT35), .A2(n1146), .ZN(n1268) );
XOR2_X1 U964 ( .A(n1269), .B(G101), .Z(n1146) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U966 ( .A1(G107), .A2(n1125), .ZN(n1271) );
XOR2_X1 U967 ( .A(n1272), .B(KEYINPUT23), .Z(n1270) );
NAND2_X1 U968 ( .A1(G104), .A2(n1273), .ZN(n1272) );
INV_X1 U969 ( .A(n1192), .ZN(n1185) );
NAND2_X1 U970 ( .A1(n1274), .A2(n1054), .ZN(n1192) );
NAND3_X1 U971 ( .A1(n1210), .A2(n1068), .A3(G952), .ZN(n1054) );
XOR2_X1 U972 ( .A(KEYINPUT45), .B(n1275), .Z(n1274) );
AND4_X1 U973 ( .A1(n1098), .A2(n1210), .A3(G902), .A4(G953), .ZN(n1275) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1210) );
INV_X1 U975 ( .A(G898), .ZN(n1098) );
INV_X1 U976 ( .A(n1184), .ZN(n1049) );
NOR2_X1 U977 ( .A1(n1052), .A2(n1051), .ZN(n1184) );
INV_X1 U978 ( .A(n1056), .ZN(n1051) );
NAND2_X1 U979 ( .A1(G214), .A2(n1276), .ZN(n1056) );
INV_X1 U980 ( .A(n1203), .ZN(n1052) );
XNOR2_X1 U981 ( .A(n1062), .B(n1277), .ZN(n1203) );
NOR2_X1 U982 ( .A1(KEYINPUT21), .A2(n1064), .ZN(n1277) );
NAND2_X1 U983 ( .A1(G210), .A2(n1276), .ZN(n1064) );
NAND2_X1 U984 ( .A1(n1278), .A2(n1232), .ZN(n1276) );
INV_X1 U985 ( .A(G237), .ZN(n1278) );
NAND2_X1 U986 ( .A1(n1279), .A2(n1232), .ZN(n1062) );
XOR2_X1 U987 ( .A(n1280), .B(n1194), .Z(n1279) );
XOR2_X1 U988 ( .A(n1281), .B(n1282), .Z(n1194) );
XOR2_X1 U989 ( .A(n1103), .B(n1100), .Z(n1282) );
XNOR2_X1 U990 ( .A(n1283), .B(n1284), .ZN(n1100) );
XNOR2_X1 U991 ( .A(G113), .B(KEYINPUT39), .ZN(n1283) );
XOR2_X1 U992 ( .A(G110), .B(G122), .Z(n1103) );
XOR2_X1 U993 ( .A(n1285), .B(n1286), .Z(n1281) );
XOR2_X1 U994 ( .A(G125), .B(n1287), .Z(n1286) );
AND2_X1 U995 ( .A1(n1068), .A2(G224), .ZN(n1287) );
NAND2_X1 U996 ( .A1(KEYINPUT36), .A2(n1101), .ZN(n1285) );
XOR2_X1 U997 ( .A(n1288), .B(n1289), .Z(n1101) );
XOR2_X1 U998 ( .A(KEYINPUT13), .B(G101), .Z(n1289) );
NAND2_X1 U999 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
NAND2_X1 U1000 ( .A1(KEYINPUT5), .A2(n1292), .ZN(n1291) );
INV_X1 U1001 ( .A(n1293), .ZN(n1292) );
NAND2_X1 U1002 ( .A1(KEYINPUT53), .A2(n1293), .ZN(n1290) );
XOR2_X1 U1003 ( .A(n1294), .B(n1125), .Z(n1293) );
INV_X1 U1004 ( .A(G104), .ZN(n1125) );
NAND2_X1 U1005 ( .A1(KEYINPUT42), .A2(n1273), .ZN(n1294) );
INV_X1 U1006 ( .A(G107), .ZN(n1273) );
NAND2_X1 U1007 ( .A1(KEYINPUT44), .A2(n1196), .ZN(n1280) );
NOR2_X1 U1008 ( .A1(n1205), .A2(n1061), .ZN(n1190) );
INV_X1 U1009 ( .A(n1204), .ZN(n1061) );
XNOR2_X1 U1010 ( .A(n1295), .B(n1110), .ZN(n1204) );
AND2_X1 U1011 ( .A1(G217), .A2(n1256), .ZN(n1110) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1232), .ZN(n1256) );
NAND2_X1 U1013 ( .A1(n1296), .A2(n1232), .ZN(n1295) );
XNOR2_X1 U1014 ( .A(n1113), .B(n1297), .ZN(n1296) );
INV_X1 U1015 ( .A(n1112), .ZN(n1297) );
XNOR2_X1 U1016 ( .A(n1298), .B(n1299), .ZN(n1112) );
XNOR2_X1 U1017 ( .A(G110), .B(n1300), .ZN(n1299) );
NAND2_X1 U1018 ( .A1(KEYINPUT47), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1019 ( .A(G146), .B(n1253), .Z(n1301) );
XOR2_X1 U1020 ( .A(G125), .B(G140), .Z(n1253) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1240), .ZN(n1298) );
AND2_X1 U1022 ( .A1(G234), .A2(n1068), .ZN(n1240) );
XNOR2_X1 U1023 ( .A(n1216), .B(n1302), .ZN(n1113) );
XOR2_X1 U1024 ( .A(G137), .B(G128), .Z(n1302) );
XNOR2_X1 U1025 ( .A(n1303), .B(G472), .ZN(n1205) );
NAND2_X1 U1026 ( .A1(n1304), .A2(n1232), .ZN(n1303) );
INV_X1 U1027 ( .A(G902), .ZN(n1232) );
XOR2_X1 U1028 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1029 ( .A(n1134), .B(n1307), .Z(n1306) );
NOR2_X1 U1030 ( .A1(KEYINPUT32), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1031 ( .A(n1133), .B(n1139), .ZN(n1308) );
INV_X1 U1032 ( .A(n1261), .ZN(n1139) );
XOR2_X1 U1033 ( .A(G131), .B(n1079), .Z(n1261) );
XOR2_X1 U1034 ( .A(G134), .B(G137), .Z(n1079) );
XOR2_X1 U1035 ( .A(n1309), .B(n1310), .Z(n1133) );
XNOR2_X1 U1036 ( .A(G113), .B(n1196), .ZN(n1310) );
NAND3_X1 U1037 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1196) );
NAND2_X1 U1038 ( .A1(G128), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1039 ( .A1(n1315), .A2(n1247), .ZN(n1314) );
NAND2_X1 U1040 ( .A1(KEYINPUT46), .A2(n1316), .ZN(n1312) );
OR3_X1 U1041 ( .A1(n1315), .A2(KEYINPUT46), .A3(n1316), .ZN(n1311) );
INV_X1 U1042 ( .A(n1247), .ZN(n1316) );
XOR2_X1 U1043 ( .A(G143), .B(G146), .Z(n1247) );
XOR2_X1 U1044 ( .A(n1317), .B(G128), .Z(n1315) );
XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(KEYINPUT27), .ZN(n1317) );
NAND3_X1 U1046 ( .A1(n1318), .A2(n1319), .A3(KEYINPUT37), .ZN(n1309) );
OR2_X1 U1047 ( .A1(n1284), .A2(KEYINPUT14), .ZN(n1319) );
XNOR2_X1 U1048 ( .A(G116), .B(n1216), .ZN(n1284) );
NAND3_X1 U1049 ( .A1(G116), .A2(n1216), .A3(KEYINPUT14), .ZN(n1318) );
INV_X1 U1050 ( .A(G119), .ZN(n1216) );
AND3_X1 U1051 ( .A1(G210), .A2(n1068), .A3(n1320), .ZN(n1134) );
XNOR2_X1 U1052 ( .A(G237), .B(KEYINPUT8), .ZN(n1320) );
INV_X1 U1053 ( .A(G953), .ZN(n1068) );
XNOR2_X1 U1054 ( .A(G101), .B(KEYINPUT38), .ZN(n1305) );
NOR2_X1 U1055 ( .A1(KEYINPUT22), .A2(n1321), .ZN(n1229) );
XOR2_X1 U1056 ( .A(KEYINPUT15), .B(G110), .Z(n1321) );
endmodule


