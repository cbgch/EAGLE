//Key = 0101000001000010001111101101100110000101111011101100001011001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372;

XNOR2_X1 U754 ( .A(G107), .B(n1051), .ZN(G9) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U758 ( .A(KEYINPUT30), .ZN(n1059) );
NOR4_X1 U759 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1063), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1062), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U764 ( .A1(n1061), .A2(KEYINPUT30), .A3(n1060), .ZN(n1068) );
NOR3_X1 U765 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1065) );
XOR2_X1 U766 ( .A(KEYINPUT48), .B(n1073), .Z(n1070) );
NAND3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1073), .A2(n1077), .ZN(n1076) );
NAND2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND2_X1 U771 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1083) );
OR2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U776 ( .A(n1093), .B(KEYINPUT35), .Z(n1078) );
NAND3_X1 U777 ( .A1(n1071), .A2(n1072), .A3(n1094), .ZN(n1093) );
INV_X1 U778 ( .A(n1063), .ZN(n1094) );
NAND3_X1 U779 ( .A1(n1089), .A2(n1085), .A3(n1082), .ZN(n1063) );
INV_X1 U780 ( .A(n1095), .ZN(n1082) );
NOR3_X1 U781 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1052) );
INV_X1 U782 ( .A(n1074), .ZN(n1096) );
NAND4_X1 U783 ( .A1(n1097), .A2(n1085), .A3(n1098), .A4(n1099), .ZN(n1074) );
AND4_X1 U784 ( .A1(n1060), .A2(n1072), .A3(n1100), .A4(n1101), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1102), .B(n1103), .Z(n1100) );
XOR2_X1 U786 ( .A(KEYINPUT54), .B(G475), .Z(n1103) );
XOR2_X1 U787 ( .A(n1104), .B(n1105), .Z(n1098) );
XNOR2_X1 U788 ( .A(n1061), .B(KEYINPUT12), .ZN(n1097) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(G72) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1075), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1106) );
NAND2_X1 U793 ( .A1(n1113), .A2(n1075), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND3_X1 U795 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1114) );
XNOR2_X1 U796 ( .A(n1119), .B(KEYINPUT45), .ZN(n1118) );
NAND3_X1 U797 ( .A1(G900), .A2(n1115), .A3(G953), .ZN(n1111) );
XNOR2_X1 U798 ( .A(n1120), .B(n1121), .ZN(n1115) );
XNOR2_X1 U799 ( .A(n1122), .B(n1123), .ZN(n1121) );
XNOR2_X1 U800 ( .A(G131), .B(n1124), .ZN(n1120) );
NOR2_X1 U801 ( .A1(KEYINPUT0), .A2(n1125), .ZN(n1124) );
XOR2_X1 U802 ( .A(G140), .B(G125), .Z(n1125) );
XOR2_X1 U803 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U804 ( .A1(n1128), .A2(n1075), .ZN(n1127) );
AND2_X1 U805 ( .A1(G224), .A2(G898), .ZN(n1128) );
NAND2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1131), .A2(n1075), .ZN(n1130) );
XNOR2_X1 U808 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND3_X1 U809 ( .A1(n1132), .A2(n1134), .A3(G953), .ZN(n1129) );
INV_X1 U810 ( .A(n1135), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XOR2_X1 U812 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XNOR2_X1 U815 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U816 ( .A1(n1145), .A2(n1141), .ZN(n1144) );
INV_X1 U817 ( .A(G478), .ZN(n1145) );
NOR2_X1 U818 ( .A1(n1136), .A2(n1146), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
AND2_X1 U820 ( .A1(n1150), .A2(KEYINPUT7), .ZN(n1149) );
NOR2_X1 U821 ( .A1(KEYINPUT7), .A2(n1151), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1152), .A2(n1102), .ZN(n1151) );
NOR2_X1 U823 ( .A1(n1153), .A2(n1150), .ZN(n1152) );
AND2_X1 U824 ( .A1(n1055), .A2(G475), .ZN(n1153) );
NOR3_X1 U825 ( .A1(n1141), .A2(n1154), .A3(n1155), .ZN(n1147) );
INV_X1 U826 ( .A(G475), .ZN(n1155) );
NOR2_X1 U827 ( .A1(KEYINPUT7), .A2(n1150), .ZN(n1154) );
XOR2_X1 U828 ( .A(G104), .B(n1156), .Z(G6) );
NOR2_X1 U829 ( .A1(n1136), .A2(n1157), .ZN(G57) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U831 ( .A(G101), .B(n1160), .Z(n1159) );
NOR2_X1 U832 ( .A1(KEYINPUT59), .A2(n1161), .ZN(n1158) );
XOR2_X1 U833 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U834 ( .A(n1164), .B(n1165), .Z(n1162) );
NOR2_X1 U835 ( .A1(n1166), .A2(n1141), .ZN(n1165) );
INV_X1 U836 ( .A(G472), .ZN(n1166) );
NAND2_X1 U837 ( .A1(KEYINPUT56), .A2(n1167), .ZN(n1164) );
NOR2_X1 U838 ( .A1(n1136), .A2(n1168), .ZN(G54) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U841 ( .A1(n1173), .A2(KEYINPUT3), .ZN(n1171) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U843 ( .A1(G110), .A2(KEYINPUT5), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1169) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1141), .ZN(n1179) );
INV_X1 U847 ( .A(G469), .ZN(n1180) );
NAND2_X1 U848 ( .A1(KEYINPUT60), .A2(n1181), .ZN(n1176) );
NOR2_X1 U849 ( .A1(n1136), .A2(n1182), .ZN(G51) );
XOR2_X1 U850 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U851 ( .A(n1132), .B(n1185), .Z(n1184) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1183) );
XOR2_X1 U853 ( .A(G125), .B(n1188), .Z(n1187) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1141), .ZN(n1186) );
NAND2_X1 U855 ( .A1(G902), .A2(n1055), .ZN(n1141) );
NAND4_X1 U856 ( .A1(n1116), .A2(n1133), .A3(n1119), .A4(n1117), .ZN(n1055) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1117) );
AND4_X1 U858 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1119) );
NAND3_X1 U859 ( .A1(n1089), .A2(n1196), .A3(n1197), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1069), .ZN(n1192) );
AND4_X1 U861 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1133) );
AND4_X1 U862 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1051), .ZN(n1202) );
NAND3_X1 U863 ( .A1(n1206), .A2(n1191), .A3(n1085), .ZN(n1051) );
NOR2_X1 U864 ( .A1(n1207), .A2(n1156), .ZN(n1201) );
AND3_X1 U865 ( .A1(n1085), .A2(n1206), .A3(n1208), .ZN(n1156) );
INV_X1 U866 ( .A(n1209), .ZN(n1207) );
NAND3_X1 U867 ( .A1(n1206), .A2(n1210), .A3(n1091), .ZN(n1200) );
XOR2_X1 U868 ( .A(KEYINPUT51), .B(n1089), .Z(n1210) );
NAND2_X1 U869 ( .A1(n1069), .A2(n1211), .ZN(n1199) );
XNOR2_X1 U870 ( .A(KEYINPUT2), .B(n1212), .ZN(n1211) );
AND3_X1 U871 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1116) );
AND2_X1 U872 ( .A1(G953), .A2(n1216), .ZN(n1136) );
XOR2_X1 U873 ( .A(KEYINPUT14), .B(G952), .Z(n1216) );
XNOR2_X1 U874 ( .A(G146), .B(n1217), .ZN(G48) );
NAND2_X1 U875 ( .A1(n1069), .A2(n1218), .ZN(n1217) );
XOR2_X1 U876 ( .A(KEYINPUT38), .B(n1198), .Z(n1218) );
AND3_X1 U877 ( .A1(n1219), .A2(n1208), .A3(n1197), .ZN(n1198) );
NAND2_X1 U878 ( .A1(n1220), .A2(n1221), .ZN(G45) );
OR2_X1 U879 ( .A1(n1194), .A2(G143), .ZN(n1221) );
XOR2_X1 U880 ( .A(n1222), .B(KEYINPUT8), .Z(n1220) );
NAND2_X1 U881 ( .A1(G143), .A2(n1194), .ZN(n1222) );
NAND4_X1 U882 ( .A1(n1223), .A2(n1224), .A3(n1069), .A4(n1225), .ZN(n1194) );
NOR2_X1 U883 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U884 ( .A(n1174), .B(n1195), .Z(G42) );
NAND3_X1 U885 ( .A1(n1091), .A2(n1208), .A3(n1196), .ZN(n1195) );
XOR2_X1 U886 ( .A(n1228), .B(n1229), .Z(G39) );
NAND3_X1 U887 ( .A1(n1196), .A2(n1230), .A3(n1089), .ZN(n1229) );
XOR2_X1 U888 ( .A(KEYINPUT10), .B(n1197), .Z(n1230) );
XNOR2_X1 U889 ( .A(G134), .B(n1213), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1092), .A2(n1191), .A3(n1196), .ZN(n1213) );
NAND2_X1 U891 ( .A1(n1231), .A2(n1232), .ZN(G33) );
NAND2_X1 U892 ( .A1(G131), .A2(n1215), .ZN(n1232) );
XOR2_X1 U893 ( .A(KEYINPUT40), .B(n1233), .Z(n1231) );
NOR2_X1 U894 ( .A1(G131), .A2(n1215), .ZN(n1233) );
NAND3_X1 U895 ( .A1(n1092), .A2(n1208), .A3(n1196), .ZN(n1215) );
AND2_X1 U896 ( .A1(n1219), .A2(n1073), .ZN(n1196) );
NOR2_X1 U897 ( .A1(n1061), .A2(n1234), .ZN(n1073) );
NAND3_X1 U898 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(G30) );
NAND2_X1 U899 ( .A1(G128), .A2(n1238), .ZN(n1237) );
NAND2_X1 U900 ( .A1(KEYINPUT26), .A2(n1239), .ZN(n1236) );
NAND2_X1 U901 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
INV_X1 U902 ( .A(n1238), .ZN(n1241) );
XNOR2_X1 U903 ( .A(KEYINPUT13), .B(G128), .ZN(n1240) );
NAND2_X1 U904 ( .A1(n1242), .A2(n1243), .ZN(n1235) );
INV_X1 U905 ( .A(KEYINPUT26), .ZN(n1243) );
NAND2_X1 U906 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
OR3_X1 U907 ( .A1(n1238), .A2(G128), .A3(KEYINPUT13), .ZN(n1245) );
NAND2_X1 U908 ( .A1(n1246), .A2(n1190), .ZN(n1238) );
AND3_X1 U909 ( .A1(n1219), .A2(n1069), .A3(n1197), .ZN(n1190) );
INV_X1 U910 ( .A(n1226), .ZN(n1219) );
NAND3_X1 U911 ( .A1(n1072), .A2(n1247), .A3(n1071), .ZN(n1226) );
XOR2_X1 U912 ( .A(n1088), .B(KEYINPUT24), .Z(n1246) );
NAND2_X1 U913 ( .A1(KEYINPUT13), .A2(G128), .ZN(n1244) );
XOR2_X1 U914 ( .A(n1248), .B(n1209), .Z(G3) );
NAND2_X1 U915 ( .A1(n1249), .A2(n1092), .ZN(n1209) );
XNOR2_X1 U916 ( .A(G125), .B(n1214), .ZN(G27) );
NAND3_X1 U917 ( .A1(n1091), .A2(n1080), .A3(n1250), .ZN(n1214) );
AND3_X1 U918 ( .A1(n1208), .A2(n1247), .A3(n1069), .ZN(n1250) );
NAND2_X1 U919 ( .A1(n1251), .A2(n1095), .ZN(n1247) );
NAND2_X1 U920 ( .A1(n1252), .A2(n1110), .ZN(n1251) );
INV_X1 U921 ( .A(G900), .ZN(n1110) );
XOR2_X1 U922 ( .A(n1205), .B(n1253), .Z(G24) );
NAND2_X1 U923 ( .A1(KEYINPUT44), .A2(G122), .ZN(n1253) );
NAND4_X1 U924 ( .A1(n1254), .A2(n1085), .A3(n1223), .A4(n1224), .ZN(n1205) );
INV_X1 U925 ( .A(n1255), .ZN(n1224) );
INV_X1 U926 ( .A(n1101), .ZN(n1223) );
NOR2_X1 U927 ( .A1(n1256), .A2(n1257), .ZN(n1085) );
XOR2_X1 U928 ( .A(n1258), .B(n1204), .Z(G21) );
NAND3_X1 U929 ( .A1(n1089), .A2(n1254), .A3(n1197), .ZN(n1204) );
AND2_X1 U930 ( .A1(n1257), .A2(n1256), .ZN(n1197) );
INV_X1 U931 ( .A(n1259), .ZN(n1257) );
XOR2_X1 U932 ( .A(n1203), .B(n1260), .Z(G18) );
NAND2_X1 U933 ( .A1(KEYINPUT32), .A2(G116), .ZN(n1260) );
NAND3_X1 U934 ( .A1(n1092), .A2(n1191), .A3(n1254), .ZN(n1203) );
AND3_X1 U935 ( .A1(n1069), .A2(n1261), .A3(n1080), .ZN(n1254) );
INV_X1 U936 ( .A(n1088), .ZN(n1191) );
NAND2_X1 U937 ( .A1(n1262), .A2(n1255), .ZN(n1088) );
XOR2_X1 U938 ( .A(n1101), .B(KEYINPUT37), .Z(n1262) );
XOR2_X1 U939 ( .A(G113), .B(n1263), .Z(G15) );
NOR2_X1 U940 ( .A1(n1264), .A2(n1212), .ZN(n1263) );
NAND4_X1 U941 ( .A1(n1092), .A2(n1080), .A3(n1208), .A4(n1261), .ZN(n1212) );
INV_X1 U942 ( .A(n1087), .ZN(n1208) );
NAND2_X1 U943 ( .A1(n1265), .A2(n1101), .ZN(n1087) );
XOR2_X1 U944 ( .A(n1255), .B(KEYINPUT28), .Z(n1265) );
INV_X1 U945 ( .A(n1062), .ZN(n1080) );
NAND2_X1 U946 ( .A1(n1266), .A2(n1072), .ZN(n1062) );
INV_X1 U947 ( .A(n1227), .ZN(n1092) );
NAND2_X1 U948 ( .A1(n1259), .A2(n1256), .ZN(n1227) );
XNOR2_X1 U949 ( .A(G110), .B(n1267), .ZN(G12) );
NAND2_X1 U950 ( .A1(n1249), .A2(n1091), .ZN(n1267) );
NOR2_X1 U951 ( .A1(n1256), .A2(n1259), .ZN(n1091) );
XOR2_X1 U952 ( .A(n1140), .B(n1268), .Z(n1259) );
NOR2_X1 U953 ( .A1(G902), .A2(n1269), .ZN(n1268) );
XOR2_X1 U954 ( .A(KEYINPUT42), .B(n1270), .Z(n1269) );
INV_X1 U955 ( .A(n1138), .ZN(n1270) );
XOR2_X1 U956 ( .A(n1271), .B(n1272), .Z(n1138) );
XOR2_X1 U957 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR3_X1 U958 ( .A1(n1275), .A2(KEYINPUT50), .A3(n1276), .ZN(n1274) );
NOR4_X1 U959 ( .A1(G953), .A2(n1228), .A3(n1277), .A4(n1278), .ZN(n1276) );
NOR2_X1 U960 ( .A1(n1279), .A2(n1280), .ZN(n1275) );
XOR2_X1 U961 ( .A(n1228), .B(KEYINPUT63), .Z(n1280) );
NOR3_X1 U962 ( .A1(n1278), .A2(G953), .A3(n1277), .ZN(n1279) );
INV_X1 U963 ( .A(G221), .ZN(n1277) );
INV_X1 U964 ( .A(G234), .ZN(n1278) );
NOR2_X1 U965 ( .A1(n1281), .A2(n1282), .ZN(n1273) );
XOR2_X1 U966 ( .A(KEYINPUT47), .B(n1283), .Z(n1282) );
NOR2_X1 U967 ( .A1(G110), .A2(n1284), .ZN(n1283) );
INV_X1 U968 ( .A(n1285), .ZN(n1284) );
NOR2_X1 U969 ( .A1(n1285), .A2(n1286), .ZN(n1281) );
XOR2_X1 U970 ( .A(KEYINPUT19), .B(G110), .Z(n1286) );
XNOR2_X1 U971 ( .A(G128), .B(n1287), .ZN(n1285) );
NOR2_X1 U972 ( .A1(KEYINPUT29), .A2(n1258), .ZN(n1287) );
INV_X1 U973 ( .A(G119), .ZN(n1258) );
NAND2_X1 U974 ( .A1(n1288), .A2(KEYINPUT62), .ZN(n1271) );
XOR2_X1 U975 ( .A(n1289), .B(n1290), .Z(n1288) );
NAND2_X1 U976 ( .A1(KEYINPUT22), .A2(n1174), .ZN(n1289) );
NAND2_X1 U977 ( .A1(G217), .A2(n1291), .ZN(n1140) );
XNOR2_X1 U978 ( .A(n1292), .B(G472), .ZN(n1256) );
NAND2_X1 U979 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U980 ( .A(n1295), .B(n1296), .Z(n1293) );
XOR2_X1 U981 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U982 ( .A(n1248), .B(KEYINPUT34), .Z(n1298) );
NAND2_X1 U983 ( .A1(n1299), .A2(n1160), .ZN(n1297) );
AND3_X1 U984 ( .A1(n1300), .A2(n1075), .A3(G210), .ZN(n1160) );
XNOR2_X1 U985 ( .A(KEYINPUT55), .B(KEYINPUT53), .ZN(n1299) );
XNOR2_X1 U986 ( .A(n1163), .B(n1167), .ZN(n1295) );
XNOR2_X1 U987 ( .A(n1301), .B(G113), .ZN(n1167) );
XNOR2_X1 U988 ( .A(n1302), .B(n1303), .ZN(n1163) );
XOR2_X1 U989 ( .A(KEYINPUT52), .B(n1304), .Z(n1303) );
AND2_X1 U990 ( .A1(n1089), .A2(n1206), .ZN(n1249) );
AND4_X1 U991 ( .A1(n1071), .A2(n1069), .A3(n1261), .A4(n1072), .ZN(n1206) );
NAND2_X1 U992 ( .A1(G221), .A2(n1291), .ZN(n1072) );
NAND2_X1 U993 ( .A1(G234), .A2(n1294), .ZN(n1291) );
NAND2_X1 U994 ( .A1(n1095), .A2(n1305), .ZN(n1261) );
NAND2_X1 U995 ( .A1(n1252), .A2(n1135), .ZN(n1305) );
XNOR2_X1 U996 ( .A(G898), .B(KEYINPUT43), .ZN(n1135) );
AND3_X1 U997 ( .A1(G902), .A2(n1306), .A3(G953), .ZN(n1252) );
NAND3_X1 U998 ( .A1(n1306), .A2(n1075), .A3(G952), .ZN(n1095) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1306) );
INV_X1 U1000 ( .A(n1264), .ZN(n1069) );
NAND2_X1 U1001 ( .A1(n1307), .A2(n1061), .ZN(n1264) );
XOR2_X1 U1002 ( .A(n1308), .B(n1189), .Z(n1061) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1309), .ZN(n1189) );
NAND3_X1 U1004 ( .A1(n1310), .A2(n1294), .A3(n1311), .ZN(n1308) );
XOR2_X1 U1005 ( .A(KEYINPUT1), .B(n1312), .Z(n1311) );
NOR2_X1 U1006 ( .A1(n1313), .A2(n1132), .ZN(n1312) );
NAND2_X1 U1007 ( .A1(n1313), .A2(n1132), .ZN(n1310) );
XNOR2_X1 U1008 ( .A(n1314), .B(n1315), .ZN(n1132) );
XOR2_X1 U1009 ( .A(n1301), .B(n1316), .Z(n1315) );
XNOR2_X1 U1010 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U1011 ( .A1(KEYINPUT15), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U1012 ( .A(G116), .B(n1320), .ZN(n1301) );
XOR2_X1 U1013 ( .A(KEYINPUT20), .B(G119), .Z(n1320) );
XOR2_X1 U1014 ( .A(n1248), .B(n1321), .Z(n1314) );
XOR2_X1 U1015 ( .A(KEYINPUT39), .B(G110), .Z(n1321) );
AND2_X1 U1016 ( .A1(n1322), .A2(n1323), .ZN(n1313) );
NAND2_X1 U1017 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1018 ( .A(n1326), .B(n1185), .Z(n1324) );
INV_X1 U1019 ( .A(n1302), .ZN(n1185) );
NAND2_X1 U1020 ( .A1(n1188), .A2(n1327), .ZN(n1322) );
XOR2_X1 U1021 ( .A(n1302), .B(n1326), .Z(n1327) );
AND2_X1 U1022 ( .A1(KEYINPUT9), .A2(G125), .ZN(n1326) );
XNOR2_X1 U1023 ( .A(G146), .B(n1328), .ZN(n1302) );
INV_X1 U1024 ( .A(n1325), .ZN(n1188) );
NAND2_X1 U1025 ( .A1(G224), .A2(n1075), .ZN(n1325) );
XOR2_X1 U1026 ( .A(KEYINPUT49), .B(n1234), .Z(n1307) );
INV_X1 U1027 ( .A(n1060), .ZN(n1234) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1309), .ZN(n1060) );
NAND2_X1 U1029 ( .A1(n1329), .A2(n1294), .ZN(n1309) );
XOR2_X1 U1030 ( .A(KEYINPUT46), .B(G237), .Z(n1329) );
INV_X1 U1031 ( .A(n1266), .ZN(n1071) );
XNOR2_X1 U1032 ( .A(n1330), .B(n1105), .ZN(n1266) );
XOR2_X1 U1033 ( .A(G469), .B(KEYINPUT6), .Z(n1105) );
NAND2_X1 U1034 ( .A1(KEYINPUT31), .A2(n1104), .ZN(n1330) );
NAND2_X1 U1035 ( .A1(n1331), .A2(n1294), .ZN(n1104) );
INV_X1 U1036 ( .A(G902), .ZN(n1294) );
XOR2_X1 U1037 ( .A(n1332), .B(KEYINPUT33), .Z(n1331) );
NAND2_X1 U1038 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NAND2_X1 U1039 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
XOR2_X1 U1040 ( .A(KEYINPUT41), .B(n1337), .Z(n1333) );
NOR2_X1 U1041 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
XNOR2_X1 U1042 ( .A(n1178), .B(n1338), .ZN(n1335) );
NAND2_X1 U1043 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1044 ( .A1(G110), .A2(n1174), .ZN(n1340) );
XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n1341), .Z(n1339) );
NOR2_X1 U1046 ( .A1(G110), .A2(n1174), .ZN(n1341) );
INV_X1 U1047 ( .A(G140), .ZN(n1174) );
NOR2_X1 U1048 ( .A1(n1109), .A2(G953), .ZN(n1178) );
INV_X1 U1049 ( .A(G227), .ZN(n1109) );
XOR2_X1 U1050 ( .A(n1304), .B(n1181), .Z(n1336) );
XNOR2_X1 U1051 ( .A(n1342), .B(n1343), .ZN(n1181) );
XOR2_X1 U1052 ( .A(n1123), .B(n1319), .Z(n1343) );
XOR2_X1 U1053 ( .A(G104), .B(G107), .Z(n1319) );
XNOR2_X1 U1054 ( .A(n1344), .B(n1328), .ZN(n1123) );
XOR2_X1 U1055 ( .A(G143), .B(G128), .Z(n1328) );
XNOR2_X1 U1056 ( .A(KEYINPUT4), .B(n1345), .ZN(n1344) );
NOR2_X1 U1057 ( .A1(KEYINPUT11), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1058 ( .A(KEYINPUT27), .B(G146), .Z(n1346) );
XOR2_X1 U1059 ( .A(n1248), .B(KEYINPUT17), .Z(n1342) );
INV_X1 U1060 ( .A(G101), .ZN(n1248) );
INV_X1 U1061 ( .A(n1172), .ZN(n1304) );
XNOR2_X1 U1062 ( .A(G131), .B(n1347), .ZN(n1172) );
NOR2_X1 U1063 ( .A1(KEYINPUT36), .A2(n1122), .ZN(n1347) );
XOR2_X1 U1064 ( .A(G134), .B(n1228), .Z(n1122) );
INV_X1 U1065 ( .A(G137), .ZN(n1228) );
AND2_X1 U1066 ( .A1(n1348), .A2(n1101), .ZN(n1089) );
XOR2_X1 U1067 ( .A(n1349), .B(G478), .Z(n1101) );
NAND2_X1 U1068 ( .A1(n1350), .A2(n1143), .ZN(n1349) );
NAND2_X1 U1069 ( .A1(n1351), .A2(n1352), .ZN(n1143) );
NAND2_X1 U1070 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1071 ( .A(n1355), .B(KEYINPUT58), .Z(n1351) );
OR2_X1 U1072 ( .A1(n1354), .A2(n1353), .ZN(n1355) );
XOR2_X1 U1073 ( .A(n1356), .B(n1357), .Z(n1353) );
XOR2_X1 U1074 ( .A(G116), .B(n1358), .Z(n1357) );
XOR2_X1 U1075 ( .A(G134), .B(G122), .Z(n1358) );
XOR2_X1 U1076 ( .A(n1359), .B(G107), .Z(n1356) );
NAND2_X1 U1077 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1078 ( .A1(G128), .A2(n1362), .ZN(n1361) );
XOR2_X1 U1079 ( .A(KEYINPUT21), .B(n1363), .Z(n1360) );
NOR2_X1 U1080 ( .A1(G128), .A2(n1362), .ZN(n1363) );
INV_X1 U1081 ( .A(G143), .ZN(n1362) );
NAND3_X1 U1082 ( .A1(G234), .A2(n1075), .A3(G217), .ZN(n1354) );
XOR2_X1 U1083 ( .A(KEYINPUT25), .B(G902), .Z(n1350) );
XOR2_X1 U1084 ( .A(n1255), .B(KEYINPUT61), .Z(n1348) );
XOR2_X1 U1085 ( .A(n1364), .B(G475), .Z(n1255) );
NAND2_X1 U1086 ( .A1(KEYINPUT18), .A2(n1102), .ZN(n1364) );
NOR2_X1 U1087 ( .A1(n1150), .A2(G902), .ZN(n1102) );
XOR2_X1 U1088 ( .A(n1365), .B(n1366), .Z(n1150) );
XOR2_X1 U1089 ( .A(n1317), .B(n1367), .Z(n1366) );
XOR2_X1 U1090 ( .A(n1368), .B(n1290), .Z(n1367) );
XOR2_X1 U1091 ( .A(G125), .B(G146), .Z(n1290) );
NOR2_X1 U1092 ( .A1(G104), .A2(KEYINPUT16), .ZN(n1368) );
XOR2_X1 U1093 ( .A(G113), .B(G122), .Z(n1317) );
XOR2_X1 U1094 ( .A(n1369), .B(n1370), .Z(n1365) );
XOR2_X1 U1095 ( .A(G143), .B(G140), .Z(n1370) );
XNOR2_X1 U1096 ( .A(G131), .B(n1371), .ZN(n1369) );
NOR2_X1 U1097 ( .A1(n1372), .A2(KEYINPUT23), .ZN(n1371) );
AND3_X1 U1098 ( .A1(G214), .A2(n1075), .A3(n1300), .ZN(n1372) );
INV_X1 U1099 ( .A(G237), .ZN(n1300) );
INV_X1 U1100 ( .A(G953), .ZN(n1075) );
endmodule


