//Key = 1101111010001110101011011110010001100011101011000100000000111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327;

XNOR2_X1 U737 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U748 ( .A1(KEYINPUT30), .A2(n1037), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
XNOR2_X1 U752 ( .A(KEYINPUT63), .B(n1044), .ZN(n1042) );
AND3_X1 U753 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1027) );
NOR3_X1 U754 ( .A1(n1030), .A2(n1048), .A3(n1039), .ZN(n1023) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR3_X1 U756 ( .A1(n1051), .A2(n1034), .A3(n1052), .ZN(n1050) );
NOR3_X1 U757 ( .A1(n1053), .A2(KEYINPUT19), .A3(n1054), .ZN(n1049) );
XOR2_X1 U758 ( .A(KEYINPUT28), .B(n1055), .Z(n1018) );
NOR2_X1 U759 ( .A1(n1026), .A2(n1056), .ZN(n1055) );
XOR2_X1 U760 ( .A(KEYINPUT61), .B(n1057), .Z(n1056) );
NOR4_X1 U761 ( .A1(n1034), .A2(n1039), .A3(n1058), .A4(n1022), .ZN(n1057) );
NAND4_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1017) );
NAND3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(KEYINPUT19), .ZN(n1060) );
OR4_X1 U764 ( .A1(n1022), .A2(n1030), .A3(n1054), .A4(n1039), .ZN(n1064) );
XOR2_X1 U765 ( .A(n1034), .B(KEYINPUT62), .Z(n1054) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(KEYINPUT30), .ZN(n1059) );
OR4_X1 U767 ( .A1(n1022), .A2(n1030), .A3(n1037), .A4(n1034), .ZN(n1066) );
INV_X1 U768 ( .A(n1067), .ZN(n1037) );
INV_X1 U769 ( .A(n1068), .ZN(n1030) );
NOR3_X1 U770 ( .A1(n1069), .A2(G953), .A3(G952), .ZN(n1015) );
INV_X1 U771 ( .A(n1061), .ZN(n1069) );
NAND4_X1 U772 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1061) );
NOR4_X1 U773 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
XOR2_X1 U774 ( .A(n1078), .B(n1079), .Z(n1076) );
NOR2_X1 U775 ( .A1(G472), .A2(KEYINPUT43), .ZN(n1079) );
NOR3_X1 U776 ( .A1(n1026), .A2(n1080), .A3(n1081), .ZN(n1072) );
AND3_X1 U777 ( .A1(KEYINPUT45), .A2(n1082), .A3(G475), .ZN(n1081) );
NOR2_X1 U778 ( .A1(KEYINPUT45), .A2(G475), .ZN(n1080) );
INV_X1 U779 ( .A(n1065), .ZN(n1026) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U782 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U783 ( .A(n1089), .B(n1090), .ZN(n1088) );
XOR2_X1 U784 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U785 ( .A1(KEYINPUT52), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U786 ( .A(n1094), .B(G125), .ZN(n1093) );
XNOR2_X1 U787 ( .A(G128), .B(n1095), .ZN(n1087) );
XNOR2_X1 U788 ( .A(KEYINPUT36), .B(n1096), .ZN(n1095) );
NOR2_X1 U789 ( .A1(G900), .A2(n1062), .ZN(n1085) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1083) );
NAND2_X1 U791 ( .A1(n1099), .A2(G953), .ZN(n1098) );
XOR2_X1 U792 ( .A(n1100), .B(KEYINPUT7), .Z(n1099) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND3_X1 U794 ( .A1(KEYINPUT21), .A2(n1101), .A3(n1062), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U796 ( .A(n1104), .ZN(n1103) );
XOR2_X1 U797 ( .A(n1105), .B(KEYINPUT24), .Z(n1102) );
XOR2_X1 U798 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1062), .ZN(n1109) );
AND2_X1 U801 ( .A1(G224), .A2(G898), .ZN(n1110) );
NAND2_X1 U802 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U803 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U804 ( .A(n1114), .B(n1115), .Z(n1111) );
XOR2_X1 U805 ( .A(n1116), .B(G110), .Z(n1115) );
XOR2_X1 U806 ( .A(n1117), .B(KEYINPUT3), .Z(n1114) );
XNOR2_X1 U807 ( .A(KEYINPUT38), .B(KEYINPUT35), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1062), .A2(n1118), .ZN(n1106) );
NOR3_X1 U809 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(G66) );
AND3_X1 U810 ( .A1(KEYINPUT15), .A2(G953), .A3(G952), .ZN(n1121) );
NOR2_X1 U811 ( .A1(KEYINPUT15), .A2(n1122), .ZN(n1120) );
INV_X1 U812 ( .A(n1123), .ZN(n1122) );
XOR2_X1 U813 ( .A(n1124), .B(n1125), .Z(n1119) );
NAND3_X1 U814 ( .A1(n1126), .A2(n1127), .A3(KEYINPUT1), .ZN(n1124) );
NOR2_X1 U815 ( .A1(n1123), .A2(n1128), .ZN(G63) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U817 ( .A(KEYINPUT18), .B(n1131), .Z(n1130) );
AND2_X1 U818 ( .A1(G478), .A2(n1126), .ZN(n1131) );
NOR2_X1 U819 ( .A1(n1123), .A2(n1132), .ZN(G60) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U821 ( .A1(G475), .A2(n1126), .ZN(n1133) );
XNOR2_X1 U822 ( .A(G104), .B(n1135), .ZN(G6) );
NAND4_X1 U823 ( .A1(n1136), .A2(n1047), .A3(n1137), .A4(n1063), .ZN(n1135) );
NOR2_X1 U824 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XNOR2_X1 U825 ( .A(n1041), .B(KEYINPUT27), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1123), .A2(n1140), .ZN(G57) );
XOR2_X1 U827 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U828 ( .A(n1143), .B(n1144), .ZN(n1142) );
XOR2_X1 U829 ( .A(n1145), .B(n1146), .Z(n1141) );
AND2_X1 U830 ( .A1(G472), .A2(n1126), .ZN(n1146) );
NOR2_X1 U831 ( .A1(n1123), .A2(n1147), .ZN(G54) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U833 ( .A(n1144), .B(n1150), .ZN(n1149) );
XOR2_X1 U834 ( .A(KEYINPUT51), .B(n1151), .Z(n1148) );
AND2_X1 U835 ( .A1(G469), .A2(n1126), .ZN(n1151) );
NOR2_X1 U836 ( .A1(n1152), .A2(n1153), .ZN(G51) );
XNOR2_X1 U837 ( .A(n1123), .B(KEYINPUT14), .ZN(n1153) );
NOR2_X1 U838 ( .A1(n1062), .A2(G952), .ZN(n1123) );
NOR2_X1 U839 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
XOR2_X1 U840 ( .A(KEYINPUT31), .B(n1156), .Z(n1155) );
NOR2_X1 U841 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
AND2_X1 U842 ( .A1(n1158), .A2(n1157), .ZN(n1154) );
XOR2_X1 U843 ( .A(n1159), .B(n1160), .Z(n1157) );
XOR2_X1 U844 ( .A(KEYINPUT55), .B(n1161), .Z(n1160) );
NOR2_X1 U845 ( .A1(G125), .A2(KEYINPUT46), .ZN(n1161) );
NAND2_X1 U846 ( .A1(n1126), .A2(n1162), .ZN(n1158) );
AND2_X1 U847 ( .A1(n1163), .A2(n1020), .ZN(n1126) );
OR3_X1 U848 ( .A1(n1118), .A2(n1104), .A3(n1105), .ZN(n1020) );
NAND4_X1 U849 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1105) );
NAND4_X1 U850 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1104) );
NAND2_X1 U851 ( .A1(n1136), .A2(n1172), .ZN(n1171) );
NAND2_X1 U852 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U853 ( .A1(n1175), .A2(n1036), .ZN(n1174) );
NAND2_X1 U854 ( .A1(KEYINPUT58), .A2(n1176), .ZN(n1173) );
OR3_X1 U855 ( .A1(n1177), .A2(KEYINPUT58), .A3(n1136), .ZN(n1170) );
NAND4_X1 U856 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1118) );
AND4_X1 U857 ( .A1(n1014), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1181) );
NAND3_X1 U858 ( .A1(n1045), .A2(n1047), .A3(n1185), .ZN(n1014) );
NAND2_X1 U859 ( .A1(n1185), .A2(n1186), .ZN(n1180) );
NAND2_X1 U860 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U861 ( .A1(n1189), .A2(n1068), .ZN(n1188) );
XNOR2_X1 U862 ( .A(n1067), .B(KEYINPUT59), .ZN(n1189) );
NAND2_X1 U863 ( .A1(n1136), .A2(n1047), .ZN(n1187) );
NAND2_X1 U864 ( .A1(n1190), .A2(n1191), .ZN(n1178) );
XNOR2_X1 U865 ( .A(KEYINPUT9), .B(n1192), .ZN(n1163) );
XOR2_X1 U866 ( .A(n1193), .B(n1194), .Z(G48) );
XOR2_X1 U867 ( .A(KEYINPUT11), .B(G146), .Z(n1194) );
NOR2_X1 U868 ( .A1(n1058), .A2(n1177), .ZN(n1193) );
INV_X1 U869 ( .A(n1136), .ZN(n1058) );
NAND2_X1 U870 ( .A1(n1195), .A2(n1196), .ZN(G45) );
NAND2_X1 U871 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U872 ( .A(KEYINPUT47), .B(n1168), .ZN(n1197) );
NAND2_X1 U873 ( .A1(n1199), .A2(G143), .ZN(n1195) );
XNOR2_X1 U874 ( .A(KEYINPUT6), .B(n1168), .ZN(n1199) );
NAND4_X1 U875 ( .A1(n1200), .A2(n1067), .A3(n1201), .A4(n1202), .ZN(n1168) );
XNOR2_X1 U876 ( .A(G140), .B(n1203), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1204), .A2(n1065), .A3(n1205), .ZN(n1203) );
XNOR2_X1 U878 ( .A(n1041), .B(KEYINPUT0), .ZN(n1205) );
XNOR2_X1 U879 ( .A(G137), .B(n1169), .ZN(G39) );
NAND2_X1 U880 ( .A1(n1206), .A2(n1175), .ZN(n1169) );
XNOR2_X1 U881 ( .A(G134), .B(n1165), .ZN(G36) );
NAND3_X1 U882 ( .A1(n1175), .A2(n1045), .A3(n1067), .ZN(n1165) );
XNOR2_X1 U883 ( .A(n1166), .B(n1207), .ZN(G33) );
NOR2_X1 U884 ( .A1(KEYINPUT32), .A2(n1208), .ZN(n1207) );
INV_X1 U885 ( .A(G131), .ZN(n1208) );
NAND3_X1 U886 ( .A1(n1175), .A2(n1136), .A3(n1067), .ZN(n1166) );
AND3_X1 U887 ( .A1(n1041), .A2(n1209), .A3(n1065), .ZN(n1175) );
NOR2_X1 U888 ( .A1(n1052), .A2(n1210), .ZN(n1065) );
INV_X1 U889 ( .A(n1051), .ZN(n1210) );
XNOR2_X1 U890 ( .A(G128), .B(n1164), .ZN(G30) );
NAND2_X1 U891 ( .A1(n1176), .A2(n1045), .ZN(n1164) );
INV_X1 U892 ( .A(n1177), .ZN(n1176) );
NAND3_X1 U893 ( .A1(n1211), .A2(n1077), .A3(n1200), .ZN(n1177) );
AND3_X1 U894 ( .A1(n1063), .A2(n1209), .A3(n1041), .ZN(n1200) );
XNOR2_X1 U895 ( .A(G101), .B(n1212), .ZN(G3) );
NAND2_X1 U896 ( .A1(n1213), .A2(n1067), .ZN(n1212) );
XNOR2_X1 U897 ( .A(G125), .B(n1167), .ZN(G27) );
NAND3_X1 U898 ( .A1(n1063), .A2(n1046), .A3(n1204), .ZN(n1167) );
AND3_X1 U899 ( .A1(n1036), .A2(n1209), .A3(n1136), .ZN(n1204) );
NAND2_X1 U900 ( .A1(n1022), .A2(n1214), .ZN(n1209) );
NAND4_X1 U901 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1216), .ZN(n1214) );
INV_X1 U902 ( .A(G900), .ZN(n1216) );
XNOR2_X1 U903 ( .A(G122), .B(n1217), .ZN(G24) );
NAND4_X1 U904 ( .A1(n1218), .A2(n1190), .A3(n1046), .A4(n1219), .ZN(n1217) );
NOR3_X1 U905 ( .A1(n1071), .A2(n1220), .A3(n1039), .ZN(n1190) );
XNOR2_X1 U906 ( .A(n1063), .B(KEYINPUT49), .ZN(n1218) );
INV_X1 U907 ( .A(n1053), .ZN(n1063) );
XNOR2_X1 U908 ( .A(G119), .B(n1179), .ZN(G21) );
NAND2_X1 U909 ( .A1(n1206), .A2(n1191), .ZN(n1179) );
AND3_X1 U910 ( .A1(n1211), .A2(n1077), .A3(n1068), .ZN(n1206) );
XNOR2_X1 U911 ( .A(G116), .B(n1184), .ZN(G18) );
NAND3_X1 U912 ( .A1(n1067), .A2(n1045), .A3(n1191), .ZN(n1184) );
NOR2_X1 U913 ( .A1(n1202), .A2(n1071), .ZN(n1045) );
INV_X1 U914 ( .A(n1201), .ZN(n1071) );
XNOR2_X1 U915 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1067), .A2(n1136), .A3(n1191), .ZN(n1183) );
NOR3_X1 U917 ( .A1(n1034), .A2(n1138), .A3(n1053), .ZN(n1191) );
INV_X1 U918 ( .A(n1046), .ZN(n1034) );
NAND2_X1 U919 ( .A1(n1221), .A2(n1222), .ZN(n1046) );
OR2_X1 U920 ( .A1(n1223), .A2(KEYINPUT63), .ZN(n1222) );
NAND3_X1 U921 ( .A1(n1070), .A2(n1043), .A3(KEYINPUT63), .ZN(n1221) );
NOR2_X1 U922 ( .A1(n1201), .A2(n1220), .ZN(n1136) );
NOR2_X1 U923 ( .A1(n1224), .A2(n1077), .ZN(n1067) );
XNOR2_X1 U924 ( .A(G110), .B(n1182), .ZN(G12) );
NAND2_X1 U925 ( .A1(n1213), .A2(n1036), .ZN(n1182) );
NAND2_X1 U926 ( .A1(n1225), .A2(n1226), .ZN(n1036) );
OR2_X1 U927 ( .A1(n1039), .A2(KEYINPUT60), .ZN(n1226) );
INV_X1 U928 ( .A(n1047), .ZN(n1039) );
NOR2_X1 U929 ( .A1(n1077), .A2(n1211), .ZN(n1047) );
INV_X1 U930 ( .A(n1224), .ZN(n1211) );
NAND3_X1 U931 ( .A1(n1077), .A2(n1224), .A3(KEYINPUT60), .ZN(n1225) );
NAND3_X1 U932 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1224) );
NAND2_X1 U933 ( .A1(G472), .A2(n1230), .ZN(n1229) );
NAND2_X1 U934 ( .A1(n1231), .A2(n1078), .ZN(n1230) );
INV_X1 U935 ( .A(n1232), .ZN(n1231) );
NAND3_X1 U936 ( .A1(KEYINPUT39), .A2(n1232), .A3(n1078), .ZN(n1228) );
XNOR2_X1 U937 ( .A(n1233), .B(G472), .ZN(n1232) );
XNOR2_X1 U938 ( .A(KEYINPUT41), .B(KEYINPUT13), .ZN(n1233) );
OR2_X1 U939 ( .A1(n1078), .A2(KEYINPUT39), .ZN(n1227) );
NAND2_X1 U940 ( .A1(n1234), .A2(n1192), .ZN(n1078) );
XOR2_X1 U941 ( .A(n1235), .B(n1145), .Z(n1234) );
XNOR2_X1 U942 ( .A(n1236), .B(n1237), .ZN(n1145) );
NAND2_X1 U943 ( .A1(n1238), .A2(G210), .ZN(n1236) );
NAND3_X1 U944 ( .A1(n1239), .A2(n1240), .A3(KEYINPUT16), .ZN(n1235) );
NAND2_X1 U945 ( .A1(n1143), .A2(n1241), .ZN(n1240) );
INV_X1 U946 ( .A(n1144), .ZN(n1241) );
NAND2_X1 U947 ( .A1(n1242), .A2(n1144), .ZN(n1239) );
XNOR2_X1 U948 ( .A(n1143), .B(KEYINPUT53), .ZN(n1242) );
XNOR2_X1 U949 ( .A(n1243), .B(n1244), .ZN(n1143) );
XNOR2_X1 U950 ( .A(n1245), .B(G113), .ZN(n1244) );
XOR2_X1 U951 ( .A(n1246), .B(n1247), .Z(n1243) );
XNOR2_X1 U952 ( .A(n1248), .B(n1127), .ZN(n1077) );
AND2_X1 U953 ( .A1(G217), .A2(n1249), .ZN(n1127) );
NAND2_X1 U954 ( .A1(n1125), .A2(n1192), .ZN(n1248) );
XNOR2_X1 U955 ( .A(n1250), .B(n1251), .ZN(n1125) );
XNOR2_X1 U956 ( .A(n1096), .B(n1252), .ZN(n1251) );
NOR2_X1 U957 ( .A1(KEYINPUT10), .A2(n1253), .ZN(n1252) );
XOR2_X1 U958 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U959 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U960 ( .A1(KEYINPUT17), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U961 ( .A(G119), .B(KEYINPUT4), .ZN(n1258) );
XNOR2_X1 U962 ( .A(G125), .B(n1259), .ZN(n1254) );
XOR2_X1 U963 ( .A(KEYINPUT2), .B(G146), .Z(n1259) );
NAND2_X1 U964 ( .A1(n1260), .A2(G221), .ZN(n1250) );
AND2_X1 U965 ( .A1(n1068), .A2(n1185), .ZN(n1213) );
NOR3_X1 U966 ( .A1(n1053), .A2(n1138), .A3(n1223), .ZN(n1185) );
INV_X1 U967 ( .A(n1041), .ZN(n1223) );
NOR2_X1 U968 ( .A1(n1070), .A2(n1075), .ZN(n1041) );
INV_X1 U969 ( .A(n1043), .ZN(n1075) );
NAND2_X1 U970 ( .A1(G221), .A2(n1249), .ZN(n1043) );
NAND2_X1 U971 ( .A1(G234), .A2(n1192), .ZN(n1249) );
INV_X1 U972 ( .A(n1044), .ZN(n1070) );
XNOR2_X1 U973 ( .A(n1261), .B(G469), .ZN(n1044) );
NAND2_X1 U974 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U975 ( .A(n1264), .B(n1150), .ZN(n1263) );
XOR2_X1 U976 ( .A(n1265), .B(n1266), .Z(n1150) );
XOR2_X1 U977 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U978 ( .A(KEYINPUT40), .B(n1237), .ZN(n1268) );
AND2_X1 U979 ( .A1(n1062), .A2(G227), .ZN(n1267) );
XNOR2_X1 U980 ( .A(n1269), .B(n1270), .ZN(n1265) );
XNOR2_X1 U981 ( .A(n1256), .B(n1271), .ZN(n1269) );
XNOR2_X1 U982 ( .A(G140), .B(n1272), .ZN(n1256) );
NAND2_X1 U983 ( .A1(KEYINPUT42), .A2(n1144), .ZN(n1264) );
XNOR2_X1 U984 ( .A(n1091), .B(n1273), .ZN(n1144) );
NOR2_X1 U985 ( .A1(KEYINPUT22), .A2(n1096), .ZN(n1273) );
INV_X1 U986 ( .A(G137), .ZN(n1096) );
XNOR2_X1 U987 ( .A(G131), .B(G134), .ZN(n1091) );
XNOR2_X1 U988 ( .A(G902), .B(KEYINPUT57), .ZN(n1262) );
INV_X1 U989 ( .A(n1219), .ZN(n1138) );
NAND2_X1 U990 ( .A1(n1022), .A2(n1274), .ZN(n1219) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1113), .ZN(n1274) );
INV_X1 U992 ( .A(G898), .ZN(n1113) );
NAND3_X1 U993 ( .A1(n1215), .A2(n1062), .A3(G952), .ZN(n1022) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1215) );
NAND2_X1 U995 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
NAND2_X1 U996 ( .A1(G214), .A2(n1275), .ZN(n1051) );
XNOR2_X1 U997 ( .A(n1276), .B(n1162), .ZN(n1052) );
AND2_X1 U998 ( .A1(G210), .A2(n1275), .ZN(n1162) );
NAND2_X1 U999 ( .A1(n1277), .A2(n1192), .ZN(n1275) );
INV_X1 U1000 ( .A(G237), .ZN(n1277) );
NAND2_X1 U1001 ( .A1(n1278), .A2(n1192), .ZN(n1276) );
XNOR2_X1 U1002 ( .A(G125), .B(n1159), .ZN(n1278) );
XOR2_X1 U1003 ( .A(n1279), .B(n1280), .Z(n1159) );
XOR2_X1 U1004 ( .A(n1246), .B(n1281), .Z(n1280) );
NAND2_X1 U1005 ( .A1(G224), .A2(n1062), .ZN(n1281) );
NAND2_X1 U1006 ( .A1(KEYINPUT8), .A2(n1271), .ZN(n1246) );
INV_X1 U1007 ( .A(n1089), .ZN(n1271) );
XOR2_X1 U1008 ( .A(G143), .B(G146), .Z(n1089) );
XOR2_X1 U1009 ( .A(n1116), .B(n1272), .Z(n1279) );
XNOR2_X1 U1010 ( .A(G110), .B(n1245), .ZN(n1272) );
INV_X1 U1011 ( .A(G128), .ZN(n1245) );
XNOR2_X1 U1012 ( .A(n1282), .B(n1283), .ZN(n1116) );
XOR2_X1 U1013 ( .A(n1284), .B(n1285), .Z(n1283) );
NAND2_X1 U1014 ( .A1(KEYINPUT33), .A2(n1247), .ZN(n1285) );
XOR2_X1 U1015 ( .A(G116), .B(G119), .Z(n1247) );
NAND3_X1 U1016 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1284) );
OR2_X1 U1017 ( .A1(n1237), .A2(n1289), .ZN(n1288) );
NAND3_X1 U1018 ( .A1(n1289), .A2(n1237), .A3(KEYINPUT5), .ZN(n1287) );
INV_X1 U1019 ( .A(G101), .ZN(n1237) );
NOR2_X1 U1020 ( .A1(KEYINPUT37), .A2(n1270), .ZN(n1289) );
OR2_X1 U1021 ( .A1(n1290), .A2(KEYINPUT5), .ZN(n1286) );
INV_X1 U1022 ( .A(n1270), .ZN(n1290) );
XNOR2_X1 U1023 ( .A(G107), .B(G104), .ZN(n1270) );
NOR2_X1 U1024 ( .A1(n1201), .A2(n1202), .ZN(n1068) );
INV_X1 U1025 ( .A(n1220), .ZN(n1202) );
NOR2_X1 U1026 ( .A1(n1074), .A2(n1291), .ZN(n1220) );
AND2_X1 U1027 ( .A1(G475), .A2(n1082), .ZN(n1291) );
NOR2_X1 U1028 ( .A1(n1082), .A2(G475), .ZN(n1074) );
OR2_X1 U1029 ( .A1(n1134), .A2(G902), .ZN(n1082) );
XNOR2_X1 U1030 ( .A(n1292), .B(n1293), .ZN(n1134) );
XOR2_X1 U1031 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1032 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1033 ( .A(n1298), .B(KEYINPUT44), .Z(n1297) );
NAND2_X1 U1034 ( .A1(G104), .A2(n1282), .ZN(n1298) );
NOR2_X1 U1035 ( .A1(G104), .A2(n1282), .ZN(n1296) );
XOR2_X1 U1036 ( .A(G113), .B(G122), .Z(n1282) );
AND2_X1 U1037 ( .A1(G214), .A2(n1238), .ZN(n1294) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1238) );
XOR2_X1 U1039 ( .A(n1299), .B(n1300), .Z(n1292) );
XNOR2_X1 U1040 ( .A(n1198), .B(G131), .ZN(n1300) );
INV_X1 U1041 ( .A(G143), .ZN(n1198) );
NAND2_X1 U1042 ( .A1(n1301), .A2(KEYINPUT29), .ZN(n1299) );
XOR2_X1 U1043 ( .A(n1302), .B(G146), .Z(n1301) );
NAND4_X1 U1044 ( .A1(KEYINPUT20), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1302) );
NAND3_X1 U1045 ( .A1(n1306), .A2(n1094), .A3(KEYINPUT25), .ZN(n1305) );
INV_X1 U1046 ( .A(G140), .ZN(n1094) );
INV_X1 U1047 ( .A(n1307), .ZN(n1306) );
OR2_X1 U1048 ( .A1(n1308), .A2(KEYINPUT25), .ZN(n1304) );
NAND2_X1 U1049 ( .A1(G140), .A2(n1307), .ZN(n1303) );
NAND2_X1 U1050 ( .A1(KEYINPUT23), .A2(n1308), .ZN(n1307) );
INV_X1 U1051 ( .A(G125), .ZN(n1308) );
XNOR2_X1 U1052 ( .A(n1309), .B(G478), .ZN(n1201) );
NAND2_X1 U1053 ( .A1(n1129), .A2(n1192), .ZN(n1309) );
INV_X1 U1054 ( .A(G902), .ZN(n1192) );
NAND2_X1 U1055 ( .A1(n1310), .A2(n1311), .ZN(n1129) );
NAND2_X1 U1056 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1057 ( .A1(n1314), .A2(n1315), .ZN(n1310) );
XOR2_X1 U1058 ( .A(n1316), .B(n1312), .Z(n1315) );
XNOR2_X1 U1059 ( .A(n1317), .B(n1318), .ZN(n1312) );
NOR3_X1 U1060 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1318) );
AND2_X1 U1061 ( .A1(KEYINPUT48), .A2(n1322), .ZN(n1321) );
NOR3_X1 U1062 ( .A1(KEYINPUT48), .A2(G134), .A3(n1323), .ZN(n1320) );
AND2_X1 U1063 ( .A1(n1323), .A2(G134), .ZN(n1319) );
OR2_X1 U1064 ( .A1(KEYINPUT50), .A2(n1322), .ZN(n1323) );
XNOR2_X1 U1065 ( .A(n1324), .B(n1325), .ZN(n1322) );
NOR2_X1 U1066 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1325) );
XNOR2_X1 U1067 ( .A(G128), .B(KEYINPUT54), .ZN(n1324) );
NAND2_X1 U1068 ( .A1(n1326), .A2(KEYINPUT26), .ZN(n1317) );
XNOR2_X1 U1069 ( .A(G107), .B(n1327), .ZN(n1326) );
XOR2_X1 U1070 ( .A(G122), .B(G116), .Z(n1327) );
XNOR2_X1 U1071 ( .A(KEYINPUT34), .B(KEYINPUT12), .ZN(n1316) );
INV_X1 U1072 ( .A(n1313), .ZN(n1314) );
NAND2_X1 U1073 ( .A1(G217), .A2(n1260), .ZN(n1313) );
AND2_X1 U1074 ( .A1(G234), .A2(n1062), .ZN(n1260) );
INV_X1 U1075 ( .A(G953), .ZN(n1062) );
endmodule


