//Key = 1001111000000001010101110011011001100100001011100110111000111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307;

NAND2_X1 U725 ( .A1(n995), .A2(n996), .ZN(G9) );
NAND2_X1 U726 ( .A1(n997), .A2(n998), .ZN(n996) );
XOR2_X1 U727 ( .A(n999), .B(KEYINPUT50), .Z(n997) );
XOR2_X1 U728 ( .A(KEYINPUT22), .B(n1000), .Z(n995) );
NOR2_X1 U729 ( .A1(n1001), .A2(n998), .ZN(n1000) );
XOR2_X1 U730 ( .A(n999), .B(KEYINPUT33), .Z(n1001) );
INV_X1 U731 ( .A(G107), .ZN(n999) );
NOR2_X1 U732 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR3_X1 U733 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NAND3_X1 U734 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
NAND2_X1 U735 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U736 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND3_X1 U737 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND2_X1 U738 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NAND2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1017) );
NAND2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
OR2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U745 ( .A1(n1025), .A2(n1031), .A3(n1019), .ZN(n1012) );
NAND2_X1 U746 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U747 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
OR2_X1 U748 ( .A1(n1037), .A2(n1014), .ZN(n1035) );
NAND3_X1 U749 ( .A1(n1038), .A2(n1039), .A3(n1037), .ZN(n1034) );
NAND2_X1 U750 ( .A1(n1014), .A2(n1040), .ZN(n1032) );
INV_X1 U751 ( .A(n1041), .ZN(n1010) );
NOR3_X1 U752 ( .A1(n1042), .A2(G953), .A3(G952), .ZN(n1002) );
INV_X1 U753 ( .A(n1007), .ZN(n1042) );
NAND3_X1 U754 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1007) );
NOR3_X1 U755 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
XNOR2_X1 U756 ( .A(n1049), .B(n1050), .ZN(n1048) );
NOR2_X1 U757 ( .A1(G472), .A2(KEYINPUT14), .ZN(n1050) );
XNOR2_X1 U758 ( .A(n1051), .B(n1052), .ZN(n1047) );
NOR2_X1 U759 ( .A1(n1053), .A2(KEYINPUT9), .ZN(n1052) );
XOR2_X1 U760 ( .A(n1054), .B(n1055), .Z(n1044) );
XOR2_X1 U761 ( .A(KEYINPUT35), .B(n1056), .Z(n1055) );
NAND2_X1 U762 ( .A1(KEYINPUT5), .A2(G475), .ZN(n1054) );
XOR2_X1 U763 ( .A(n1057), .B(KEYINPUT54), .Z(n1043) );
NAND3_X1 U764 ( .A1(n1058), .A2(n1037), .A3(n1019), .ZN(n1057) );
XOR2_X1 U765 ( .A(n1059), .B(n1060), .Z(n1058) );
NAND2_X1 U766 ( .A1(KEYINPUT46), .A2(n1061), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(G72) );
NAND2_X1 U768 ( .A1(n1064), .A2(n1008), .ZN(n1063) );
XNOR2_X1 U769 ( .A(n1065), .B(n1066), .ZN(n1064) );
NOR2_X1 U770 ( .A1(n1067), .A2(KEYINPUT24), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1068), .A2(G953), .ZN(n1062) );
XOR2_X1 U772 ( .A(n1065), .B(n1069), .Z(n1068) );
AND2_X1 U773 ( .A1(G227), .A2(G900), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1070), .A2(n1071), .ZN(n1065) );
NAND2_X1 U775 ( .A1(n1072), .A2(G953), .ZN(n1071) );
XOR2_X1 U776 ( .A(n1073), .B(KEYINPUT31), .Z(n1072) );
XOR2_X1 U777 ( .A(n1074), .B(n1075), .Z(n1070) );
XOR2_X1 U778 ( .A(KEYINPUT47), .B(n1076), .Z(n1075) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U780 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U781 ( .A(n1081), .B(KEYINPUT13), .Z(n1080) );
XOR2_X1 U782 ( .A(n1082), .B(n1083), .Z(n1074) );
XOR2_X1 U783 ( .A(n1084), .B(n1085), .Z(G69) );
XOR2_X1 U784 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U785 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U786 ( .A1(G898), .A2(G224), .ZN(n1088) );
NAND2_X1 U787 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U788 ( .A1(G953), .A2(n1091), .ZN(n1090) );
XOR2_X1 U789 ( .A(n1092), .B(n1093), .Z(n1089) );
XNOR2_X1 U790 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1096), .A2(G953), .ZN(n1084) );
NOR3_X1 U792 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(G66) );
NOR3_X1 U793 ( .A1(n1100), .A2(G953), .A3(G952), .ZN(n1099) );
AND2_X1 U794 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
INV_X1 U795 ( .A(KEYINPUT55), .ZN(n1100) );
XOR2_X1 U796 ( .A(n1102), .B(n1103), .Z(n1097) );
NOR2_X1 U797 ( .A1(KEYINPUT25), .A2(n1104), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1053), .A2(n1105), .ZN(n1102) );
INV_X1 U799 ( .A(n1106), .ZN(n1053) );
NOR2_X1 U800 ( .A1(n1101), .A2(n1107), .ZN(G63) );
XNOR2_X1 U801 ( .A(n1108), .B(n1109), .ZN(n1107) );
AND2_X1 U802 ( .A1(G478), .A2(n1105), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1101), .A2(n1110), .ZN(G60) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U805 ( .A(KEYINPUT20), .B(n1113), .Z(n1112) );
NOR2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1116), .B(KEYINPUT34), .Z(n1115) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1116), .ZN(n1111) );
NAND2_X1 U809 ( .A1(n1105), .A2(G475), .ZN(n1116) );
INV_X1 U810 ( .A(n1118), .ZN(n1105) );
XOR2_X1 U811 ( .A(n1114), .B(KEYINPUT19), .Z(n1117) );
XOR2_X1 U812 ( .A(n1119), .B(n1120), .Z(G6) );
NOR2_X1 U813 ( .A1(n1101), .A2(n1121), .ZN(G57) );
XOR2_X1 U814 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U815 ( .A(n1124), .B(n1125), .ZN(n1122) );
NOR2_X1 U816 ( .A1(n1126), .A2(n1118), .ZN(n1125) );
NOR2_X1 U817 ( .A1(n1101), .A2(n1127), .ZN(G54) );
XOR2_X1 U818 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U819 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U820 ( .A1(n1059), .A2(n1118), .ZN(n1130) );
INV_X1 U821 ( .A(G469), .ZN(n1059) );
XOR2_X1 U822 ( .A(n1132), .B(n1133), .Z(n1128) );
XNOR2_X1 U823 ( .A(n1134), .B(n1135), .ZN(n1133) );
NAND2_X1 U824 ( .A1(n1136), .A2(KEYINPUT4), .ZN(n1132) );
XNOR2_X1 U825 ( .A(G140), .B(n1137), .ZN(n1136) );
NOR2_X1 U826 ( .A1(G110), .A2(KEYINPUT38), .ZN(n1137) );
NOR2_X1 U827 ( .A1(n1101), .A2(n1138), .ZN(G51) );
XOR2_X1 U828 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U829 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U830 ( .A1(n1143), .A2(n1118), .ZN(n1141) );
NAND2_X1 U831 ( .A1(G902), .A2(n1144), .ZN(n1118) );
NAND2_X1 U832 ( .A1(n1096), .A2(n1067), .ZN(n1144) );
INV_X1 U833 ( .A(n1005), .ZN(n1067) );
NAND4_X1 U834 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1005) );
AND4_X1 U835 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NOR2_X1 U836 ( .A1(n1153), .A2(n1154), .ZN(n1147) );
NAND2_X1 U837 ( .A1(n1019), .A2(n1155), .ZN(n1145) );
XOR2_X1 U838 ( .A(KEYINPUT11), .B(n1156), .Z(n1155) );
INV_X1 U839 ( .A(n1006), .ZN(n1096) );
NAND2_X1 U840 ( .A1(n1157), .A2(n1158), .ZN(n1006) );
AND4_X1 U841 ( .A1(n998), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1158) );
NAND3_X1 U842 ( .A1(n1025), .A2(n1162), .A3(n1163), .ZN(n998) );
AND4_X1 U843 ( .A1(n1164), .A2(n1165), .A3(n1120), .A4(n1166), .ZN(n1157) );
OR3_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NAND3_X1 U845 ( .A1(n1025), .A2(n1162), .A3(n1170), .ZN(n1120) );
XOR2_X1 U846 ( .A(n1171), .B(n1172), .Z(n1139) );
NAND2_X1 U847 ( .A1(n1173), .A2(KEYINPUT37), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1082), .B(n1174), .Z(n1173) );
NOR2_X1 U849 ( .A1(G125), .A2(KEYINPUT28), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1008), .A2(G952), .ZN(n1101) );
NAND2_X1 U851 ( .A1(n1175), .A2(n1176), .ZN(G48) );
NAND2_X1 U852 ( .A1(n1177), .A2(n1146), .ZN(n1176) );
XOR2_X1 U853 ( .A(KEYINPUT42), .B(n1178), .Z(n1175) );
NOR2_X1 U854 ( .A1(n1146), .A2(n1177), .ZN(n1178) );
XOR2_X1 U855 ( .A(KEYINPUT1), .B(G146), .Z(n1177) );
NAND4_X1 U856 ( .A1(n1179), .A2(n1170), .A3(n1180), .A4(n1181), .ZN(n1146) );
NOR2_X1 U857 ( .A1(n1182), .A2(n1027), .ZN(n1180) );
XOR2_X1 U858 ( .A(n1183), .B(n1184), .Z(G45) );
NAND2_X1 U859 ( .A1(KEYINPUT26), .A2(n1154), .ZN(n1184) );
NOR3_X1 U860 ( .A1(n1167), .A2(n1027), .A3(n1185), .ZN(n1154) );
XOR2_X1 U861 ( .A(G140), .B(n1153), .Z(G42) );
AND3_X1 U862 ( .A1(n1019), .A2(n1040), .A3(n1186), .ZN(n1153) );
NAND2_X1 U863 ( .A1(n1187), .A2(n1188), .ZN(G39) );
NAND2_X1 U864 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U865 ( .A(KEYINPUT61), .B(n1191), .Z(n1187) );
NOR2_X1 U866 ( .A1(n1189), .A2(n1190), .ZN(n1191) );
INV_X1 U867 ( .A(G137), .ZN(n1190) );
INV_X1 U868 ( .A(n1152), .ZN(n1189) );
NAND4_X1 U869 ( .A1(n1179), .A2(n1181), .A3(n1192), .A4(n1014), .ZN(n1152) );
NOR2_X1 U870 ( .A1(n1182), .A2(n1193), .ZN(n1192) );
INV_X1 U871 ( .A(n1194), .ZN(n1179) );
XOR2_X1 U872 ( .A(n1195), .B(n1196), .Z(G36) );
NAND2_X1 U873 ( .A1(n1156), .A2(n1019), .ZN(n1196) );
NOR2_X1 U874 ( .A1(n1185), .A2(n1039), .ZN(n1156) );
INV_X1 U875 ( .A(n1163), .ZN(n1039) );
XOR2_X1 U876 ( .A(n1081), .B(n1151), .Z(G33) );
OR3_X1 U877 ( .A1(n1038), .A2(n1193), .A3(n1185), .ZN(n1151) );
NAND3_X1 U878 ( .A1(n1040), .A2(n1197), .A3(n1198), .ZN(n1185) );
INV_X1 U879 ( .A(n1182), .ZN(n1040) );
XOR2_X1 U880 ( .A(n1199), .B(KEYINPUT41), .Z(n1182) );
INV_X1 U881 ( .A(n1019), .ZN(n1193) );
NOR2_X1 U882 ( .A1(n1029), .A2(n1200), .ZN(n1019) );
XOR2_X1 U883 ( .A(n1150), .B(n1201), .Z(G30) );
NOR2_X1 U884 ( .A1(G128), .A2(KEYINPUT10), .ZN(n1201) );
NAND4_X1 U885 ( .A1(n1202), .A2(n1203), .A3(n1163), .A4(n1204), .ZN(n1150) );
NOR2_X1 U886 ( .A1(n1024), .A2(n1194), .ZN(n1204) );
XNOR2_X1 U887 ( .A(G101), .B(n1165), .ZN(G3) );
NAND3_X1 U888 ( .A1(n1014), .A2(n1162), .A3(n1198), .ZN(n1165) );
XNOR2_X1 U889 ( .A(G125), .B(n1149), .ZN(G27) );
NAND3_X1 U890 ( .A1(n1016), .A2(n1203), .A3(n1186), .ZN(n1149) );
NOR3_X1 U891 ( .A1(n1038), .A2(n1181), .A3(n1194), .ZN(n1186) );
NAND2_X1 U892 ( .A1(n1023), .A2(n1197), .ZN(n1194) );
NAND2_X1 U893 ( .A1(n1041), .A2(n1205), .ZN(n1197) );
NAND4_X1 U894 ( .A1(G902), .A2(G953), .A3(n1206), .A4(n1073), .ZN(n1205) );
INV_X1 U895 ( .A(G900), .ZN(n1073) );
XOR2_X1 U896 ( .A(G122), .B(n1207), .Z(G24) );
NOR4_X1 U897 ( .A1(KEYINPUT7), .A2(n1168), .A3(n1169), .A4(n1167), .ZN(n1207) );
NAND2_X1 U898 ( .A1(n1046), .A2(n1208), .ZN(n1167) );
INV_X1 U899 ( .A(n1025), .ZN(n1168) );
NOR2_X1 U900 ( .A1(n1023), .A2(n1181), .ZN(n1025) );
XOR2_X1 U901 ( .A(n1209), .B(n1164), .Z(G21) );
NAND4_X1 U902 ( .A1(n1210), .A2(n1181), .A3(n1023), .A4(n1014), .ZN(n1164) );
NAND2_X1 U903 ( .A1(n1211), .A2(n1212), .ZN(G18) );
NAND2_X1 U904 ( .A1(G116), .A2(n1161), .ZN(n1212) );
XOR2_X1 U905 ( .A(KEYINPUT59), .B(n1213), .Z(n1211) );
NOR2_X1 U906 ( .A1(G116), .A2(n1161), .ZN(n1213) );
NAND3_X1 U907 ( .A1(n1198), .A2(n1163), .A3(n1210), .ZN(n1161) );
NOR2_X1 U908 ( .A1(n1208), .A2(n1214), .ZN(n1163) );
XOR2_X1 U909 ( .A(G113), .B(n1215), .Z(G15) );
NOR2_X1 U910 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NOR2_X1 U911 ( .A1(KEYINPUT18), .A2(n1218), .ZN(n1217) );
INV_X1 U912 ( .A(n1160), .ZN(n1218) );
NOR2_X1 U913 ( .A1(KEYINPUT58), .A2(n1160), .ZN(n1216) );
NAND3_X1 U914 ( .A1(n1198), .A2(n1170), .A3(n1210), .ZN(n1160) );
INV_X1 U915 ( .A(n1169), .ZN(n1210) );
NAND2_X1 U916 ( .A1(n1016), .A2(n1219), .ZN(n1169) );
AND2_X1 U917 ( .A1(n1036), .A2(n1037), .ZN(n1016) );
INV_X1 U918 ( .A(n1220), .ZN(n1036) );
INV_X1 U919 ( .A(n1038), .ZN(n1170) );
NAND2_X1 U920 ( .A1(n1214), .A2(n1208), .ZN(n1038) );
INV_X1 U921 ( .A(n1021), .ZN(n1198) );
NAND2_X1 U922 ( .A1(n1181), .A2(n1221), .ZN(n1021) );
XNOR2_X1 U923 ( .A(KEYINPUT56), .B(n1023), .ZN(n1221) );
INV_X1 U924 ( .A(n1024), .ZN(n1181) );
XOR2_X1 U925 ( .A(n1159), .B(n1222), .Z(G12) );
NOR2_X1 U926 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1222) );
NAND4_X1 U927 ( .A1(n1023), .A2(n1014), .A3(n1162), .A4(n1024), .ZN(n1159) );
NAND3_X1 U928 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1024) );
NAND2_X1 U929 ( .A1(KEYINPUT63), .A2(n1049), .ZN(n1225) );
NAND3_X1 U930 ( .A1(n1226), .A2(n1227), .A3(n1126), .ZN(n1224) );
INV_X1 U931 ( .A(KEYINPUT63), .ZN(n1227) );
OR2_X1 U932 ( .A1(n1126), .A2(n1226), .ZN(n1223) );
NOR2_X1 U933 ( .A1(n1049), .A2(KEYINPUT8), .ZN(n1226) );
AND2_X1 U934 ( .A1(n1228), .A2(n1229), .ZN(n1049) );
XNOR2_X1 U935 ( .A(n1230), .B(n1123), .ZN(n1228) );
XNOR2_X1 U936 ( .A(n1231), .B(n1232), .ZN(n1123) );
XOR2_X1 U937 ( .A(G113), .B(n1134), .Z(n1232) );
XNOR2_X1 U938 ( .A(n1233), .B(n1234), .ZN(n1231) );
NOR2_X1 U939 ( .A1(KEYINPUT12), .A2(n1235), .ZN(n1234) );
XOR2_X1 U940 ( .A(n1209), .B(G116), .Z(n1235) );
NAND2_X1 U941 ( .A1(KEYINPUT44), .A2(n1124), .ZN(n1230) );
AND3_X1 U942 ( .A1(n1236), .A2(n1237), .A3(G210), .ZN(n1124) );
XOR2_X1 U943 ( .A(KEYINPUT52), .B(G953), .Z(n1236) );
INV_X1 U944 ( .A(G472), .ZN(n1126) );
AND2_X1 U945 ( .A1(n1219), .A2(n1202), .ZN(n1162) );
XOR2_X1 U946 ( .A(n1199), .B(KEYINPUT27), .Z(n1202) );
NAND2_X1 U947 ( .A1(n1220), .A2(n1037), .ZN(n1199) );
NAND2_X1 U948 ( .A1(G221), .A2(n1238), .ZN(n1037) );
XOR2_X1 U949 ( .A(n1239), .B(G469), .Z(n1220) );
NAND2_X1 U950 ( .A1(KEYINPUT53), .A2(n1061), .ZN(n1239) );
NAND2_X1 U951 ( .A1(n1240), .A2(n1229), .ZN(n1061) );
XOR2_X1 U952 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U953 ( .A(n1135), .B(n1243), .ZN(n1242) );
NOR2_X1 U954 ( .A1(KEYINPUT48), .A2(n1244), .ZN(n1243) );
XOR2_X1 U955 ( .A(n1134), .B(n1245), .Z(n1244) );
NOR2_X1 U956 ( .A1(KEYINPUT57), .A2(n1131), .ZN(n1245) );
XNOR2_X1 U957 ( .A(n1246), .B(n1233), .ZN(n1131) );
XOR2_X1 U958 ( .A(G101), .B(n1247), .Z(n1233) );
INV_X1 U959 ( .A(n1082), .ZN(n1247) );
XNOR2_X1 U960 ( .A(n1248), .B(KEYINPUT51), .ZN(n1246) );
NOR2_X1 U961 ( .A1(n1249), .A2(n1077), .ZN(n1134) );
NOR2_X1 U962 ( .A1(n1250), .A2(G131), .ZN(n1077) );
NOR2_X1 U963 ( .A1(n1081), .A2(n1079), .ZN(n1249) );
INV_X1 U964 ( .A(n1250), .ZN(n1079) );
XNOR2_X1 U965 ( .A(n1195), .B(G137), .ZN(n1250) );
INV_X1 U966 ( .A(G134), .ZN(n1195) );
INV_X1 U967 ( .A(G131), .ZN(n1081) );
NAND2_X1 U968 ( .A1(G227), .A2(n1008), .ZN(n1135) );
XOR2_X1 U969 ( .A(n1251), .B(G110), .Z(n1241) );
NAND2_X1 U970 ( .A1(n1252), .A2(KEYINPUT45), .ZN(n1251) );
XNOR2_X1 U971 ( .A(G140), .B(KEYINPUT36), .ZN(n1252) );
AND2_X1 U972 ( .A1(n1203), .A2(n1253), .ZN(n1219) );
NAND2_X1 U973 ( .A1(n1041), .A2(n1254), .ZN(n1253) );
NAND4_X1 U974 ( .A1(G902), .A2(G953), .A3(n1206), .A4(n1091), .ZN(n1254) );
INV_X1 U975 ( .A(G898), .ZN(n1091) );
NAND3_X1 U976 ( .A1(n1206), .A2(n1008), .A3(G952), .ZN(n1041) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1206) );
INV_X1 U978 ( .A(n1027), .ZN(n1203) );
NAND2_X1 U979 ( .A1(n1255), .A2(n1029), .ZN(n1027) );
XOR2_X1 U980 ( .A(n1256), .B(n1143), .Z(n1029) );
NAND2_X1 U981 ( .A1(G210), .A2(n1257), .ZN(n1143) );
NAND2_X1 U982 ( .A1(n1258), .A2(n1229), .ZN(n1256) );
XOR2_X1 U983 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U984 ( .A(n1142), .B(n1082), .Z(n1260) );
XNOR2_X1 U985 ( .A(G128), .B(n1261), .ZN(n1082) );
XNOR2_X1 U986 ( .A(n1262), .B(n1095), .ZN(n1142) );
XNOR2_X1 U987 ( .A(G110), .B(n1263), .ZN(n1095) );
NAND3_X1 U988 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1262) );
OR2_X1 U989 ( .A1(n1094), .A2(KEYINPUT30), .ZN(n1266) );
NAND3_X1 U990 ( .A1(KEYINPUT30), .A2(n1094), .A3(n1092), .ZN(n1265) );
INV_X1 U991 ( .A(n1267), .ZN(n1092) );
NAND2_X1 U992 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
NAND2_X1 U993 ( .A1(n1269), .A2(KEYINPUT30), .ZN(n1268) );
XNOR2_X1 U994 ( .A(n1094), .B(KEYINPUT0), .ZN(n1269) );
XNOR2_X1 U995 ( .A(n1270), .B(G113), .ZN(n1094) );
NAND2_X1 U996 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U997 ( .A1(G116), .A2(n1209), .ZN(n1272) );
XOR2_X1 U998 ( .A(KEYINPUT49), .B(n1273), .Z(n1271) );
NOR2_X1 U999 ( .A1(G116), .A2(n1209), .ZN(n1273) );
INV_X1 U1000 ( .A(G119), .ZN(n1209) );
XOR2_X1 U1001 ( .A(G101), .B(n1248), .Z(n1267) );
XNOR2_X1 U1002 ( .A(n1119), .B(G107), .ZN(n1248) );
INV_X1 U1003 ( .A(G104), .ZN(n1119) );
XOR2_X1 U1004 ( .A(n1274), .B(n1172), .Z(n1259) );
AND2_X1 U1005 ( .A1(n1275), .A2(G224), .ZN(n1172) );
XOR2_X1 U1006 ( .A(n1008), .B(KEYINPUT32), .Z(n1275) );
XNOR2_X1 U1007 ( .A(G125), .B(KEYINPUT62), .ZN(n1274) );
XOR2_X1 U1008 ( .A(KEYINPUT23), .B(n1200), .Z(n1255) );
INV_X1 U1009 ( .A(n1030), .ZN(n1200) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1257), .ZN(n1030) );
NAND2_X1 U1011 ( .A1(n1237), .A2(n1229), .ZN(n1257) );
NOR2_X1 U1012 ( .A1(n1046), .A2(n1208), .ZN(n1014) );
XOR2_X1 U1013 ( .A(n1056), .B(G475), .Z(n1208) );
NOR2_X1 U1014 ( .A1(n1114), .A2(G902), .ZN(n1056) );
XOR2_X1 U1015 ( .A(n1276), .B(n1277), .Z(n1114) );
XOR2_X1 U1016 ( .A(n1083), .B(n1278), .Z(n1277) );
XOR2_X1 U1017 ( .A(n1279), .B(n1261), .Z(n1278) );
XOR2_X1 U1018 ( .A(G143), .B(G146), .Z(n1261) );
NOR2_X1 U1019 ( .A1(G122), .A2(KEYINPUT39), .ZN(n1279) );
XOR2_X1 U1020 ( .A(n1280), .B(n1281), .Z(n1276) );
XOR2_X1 U1021 ( .A(G131), .B(G113), .Z(n1281) );
XOR2_X1 U1022 ( .A(n1282), .B(n1283), .Z(n1280) );
AND3_X1 U1023 ( .A1(G214), .A2(n1008), .A3(n1237), .ZN(n1283) );
INV_X1 U1024 ( .A(G237), .ZN(n1237) );
NAND2_X1 U1025 ( .A1(KEYINPUT21), .A2(n1284), .ZN(n1282) );
XOR2_X1 U1026 ( .A(KEYINPUT29), .B(G104), .Z(n1284) );
INV_X1 U1027 ( .A(n1214), .ZN(n1046) );
XOR2_X1 U1028 ( .A(n1285), .B(G478), .Z(n1214) );
NAND2_X1 U1029 ( .A1(n1108), .A2(n1229), .ZN(n1285) );
XNOR2_X1 U1030 ( .A(n1286), .B(n1287), .ZN(n1108) );
AND3_X1 U1031 ( .A1(G234), .A2(n1008), .A3(G217), .ZN(n1287) );
NAND2_X1 U1032 ( .A1(n1288), .A2(KEYINPUT17), .ZN(n1286) );
XOR2_X1 U1033 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1034 ( .A(G107), .B(n1291), .Z(n1290) );
NOR2_X1 U1035 ( .A1(KEYINPUT40), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1036 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1037 ( .A(G134), .B(G128), .Z(n1294) );
NOR2_X1 U1038 ( .A1(KEYINPUT2), .A2(n1183), .ZN(n1293) );
INV_X1 U1039 ( .A(G143), .ZN(n1183) );
NAND2_X1 U1040 ( .A1(n1295), .A2(KEYINPUT60), .ZN(n1289) );
XOR2_X1 U1041 ( .A(n1296), .B(G116), .Z(n1295) );
NAND2_X1 U1042 ( .A1(KEYINPUT6), .A2(n1263), .ZN(n1296) );
INV_X1 U1043 ( .A(G122), .ZN(n1263) );
XOR2_X1 U1044 ( .A(n1297), .B(n1051), .Z(n1023) );
NOR2_X1 U1045 ( .A1(n1104), .A2(G902), .ZN(n1051) );
XNOR2_X1 U1046 ( .A(n1298), .B(n1299), .ZN(n1104) );
XOR2_X1 U1047 ( .A(G119), .B(n1300), .Z(n1299) );
XOR2_X1 U1048 ( .A(G146), .B(G128), .Z(n1300) );
XOR2_X1 U1049 ( .A(n1301), .B(n1083), .Z(n1298) );
XOR2_X1 U1050 ( .A(G125), .B(G140), .Z(n1083) );
XNOR2_X1 U1051 ( .A(G110), .B(n1302), .ZN(n1301) );
NOR2_X1 U1052 ( .A1(KEYINPUT16), .A2(n1303), .ZN(n1302) );
NOR2_X1 U1053 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1054 ( .A(n1306), .B(KEYINPUT15), .Z(n1305) );
NAND2_X1 U1055 ( .A1(n1307), .A2(G137), .ZN(n1306) );
NOR2_X1 U1056 ( .A1(G137), .A2(n1307), .ZN(n1304) );
AND3_X1 U1057 ( .A1(G234), .A2(n1008), .A3(G221), .ZN(n1307) );
INV_X1 U1058 ( .A(G953), .ZN(n1008) );
NAND2_X1 U1059 ( .A1(KEYINPUT3), .A2(n1106), .ZN(n1297) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1238), .ZN(n1106) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1229), .ZN(n1238) );
INV_X1 U1062 ( .A(G902), .ZN(n1229) );
endmodule


