//Key = 1111011110011101111111111110011000010001110101100100100111111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330;

XNOR2_X1 U736 ( .A(n998), .B(n999), .ZN(G9) );
XNOR2_X1 U737 ( .A(KEYINPUT12), .B(n1000), .ZN(n999) );
NOR2_X1 U738 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NOR3_X1 U740 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NOR2_X1 U741 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR3_X1 U742 ( .A1(n1012), .A2(KEYINPUT44), .A3(n1013), .ZN(n1010) );
NOR3_X1 U743 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1004) );
NOR2_X1 U744 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U745 ( .A1(n1018), .A2(n1007), .ZN(n1017) );
OR3_X1 U746 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1007) );
NOR3_X1 U747 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1018) );
AND2_X1 U748 ( .A1(n1025), .A2(KEYINPUT44), .ZN(n1022) );
NOR3_X1 U749 ( .A1(n1021), .A2(n1026), .A3(n1027), .ZN(n1016) );
NOR3_X1 U750 ( .A1(n1009), .A2(n1028), .A3(n1029), .ZN(n1027) );
NOR2_X1 U751 ( .A1(n1030), .A2(n1020), .ZN(n1029) );
NOR2_X1 U752 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U753 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U754 ( .A1(n1035), .A2(n1019), .ZN(n1028) );
NOR2_X1 U755 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
AND2_X1 U756 ( .A1(n1038), .A2(KEYINPUT5), .ZN(n1036) );
INV_X1 U757 ( .A(n1025), .ZN(n1009) );
NOR2_X1 U758 ( .A1(n1025), .A2(n1039), .ZN(n1026) );
NOR3_X1 U759 ( .A1(n1019), .A2(KEYINPUT5), .A3(n1040), .ZN(n1039) );
NAND2_X1 U760 ( .A1(n1041), .A2(n1042), .ZN(n1003) );
NOR3_X1 U761 ( .A1(n1043), .A2(G952), .A3(n1005), .ZN(n1001) );
AND4_X1 U762 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1005) );
NOR4_X1 U763 ( .A1(n1048), .A2(n1049), .A3(n1034), .A4(n1050), .ZN(n1047) );
XOR2_X1 U764 ( .A(G478), .B(n1051), .Z(n1050) );
XOR2_X1 U765 ( .A(KEYINPUT37), .B(n1052), .Z(n1049) );
NOR2_X1 U766 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U767 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1048) );
XNOR2_X1 U768 ( .A(n1058), .B(KEYINPUT39), .ZN(n1057) );
NAND2_X1 U769 ( .A1(KEYINPUT28), .A2(n1059), .ZN(n1056) );
NAND2_X1 U770 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
XNOR2_X1 U771 ( .A(KEYINPUT46), .B(n1062), .ZN(n1061) );
NAND2_X1 U772 ( .A1(n1063), .A2(n1064), .ZN(n1055) );
INV_X1 U773 ( .A(KEYINPUT28), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NAND3_X1 U775 ( .A1(KEYINPUT46), .A2(n1060), .A3(n1062), .ZN(n1066) );
OR2_X1 U776 ( .A1(n1062), .A2(KEYINPUT46), .ZN(n1065) );
NOR3_X1 U777 ( .A1(n1067), .A2(n1068), .A3(n1014), .ZN(n1046) );
NOR2_X1 U778 ( .A1(G472), .A2(n1069), .ZN(n1067) );
OR2_X1 U779 ( .A1(n1062), .A2(n1060), .ZN(n1045) );
XOR2_X1 U780 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U781 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U782 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U783 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND3_X1 U784 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NAND2_X1 U785 ( .A1(G953), .A2(n1075), .ZN(n1079) );
NAND2_X1 U786 ( .A1(n1081), .A2(n1073), .ZN(n1078) );
XOR2_X1 U787 ( .A(n1082), .B(KEYINPUT10), .Z(n1076) );
NAND3_X1 U788 ( .A1(n1081), .A2(n1073), .A3(n1083), .ZN(n1082) );
INV_X1 U789 ( .A(n1080), .ZN(n1083) );
XNOR2_X1 U790 ( .A(n1084), .B(n1085), .ZN(n1080) );
XNOR2_X1 U791 ( .A(n1086), .B(n1087), .ZN(n1085) );
NOR2_X1 U792 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U793 ( .A(n1090), .B(KEYINPUT43), .Z(n1089) );
NAND3_X1 U794 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
INV_X1 U795 ( .A(n1094), .ZN(n1092) );
NOR2_X1 U796 ( .A1(n1095), .A2(n1093), .ZN(n1088) );
XOR2_X1 U797 ( .A(KEYINPUT35), .B(G131), .Z(n1093) );
NOR2_X1 U798 ( .A1(n1094), .A2(n1096), .ZN(n1095) );
NOR2_X1 U799 ( .A1(G134), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U800 ( .A(n1098), .B(n1099), .ZN(n1084) );
NAND2_X1 U801 ( .A1(KEYINPUT29), .A2(n1100), .ZN(n1099) );
NAND2_X1 U802 ( .A1(KEYINPUT2), .A2(n1101), .ZN(n1098) );
XOR2_X1 U803 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U804 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U805 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
INV_X1 U806 ( .A(n1108), .ZN(n1107) );
NAND3_X1 U807 ( .A1(G953), .A2(n1109), .A3(KEYINPUT45), .ZN(n1104) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1109) );
AND2_X1 U809 ( .A1(n1110), .A2(n1073), .ZN(n1102) );
NOR2_X1 U810 ( .A1(n1111), .A2(n1112), .ZN(G66) );
XNOR2_X1 U811 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND2_X1 U812 ( .A1(n1115), .A2(G217), .ZN(n1113) );
NOR2_X1 U813 ( .A1(n1111), .A2(n1116), .ZN(G63) );
XOR2_X1 U814 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U815 ( .A1(n1115), .A2(G478), .ZN(n1118) );
NOR2_X1 U816 ( .A1(n1111), .A2(n1119), .ZN(G60) );
XOR2_X1 U817 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND3_X1 U818 ( .A1(n1115), .A2(G475), .A3(KEYINPUT15), .ZN(n1120) );
XOR2_X1 U819 ( .A(G104), .B(n1122), .Z(G6) );
NOR2_X1 U820 ( .A1(n1111), .A2(n1123), .ZN(G57) );
XNOR2_X1 U821 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U822 ( .A(n1126), .B(n1127), .Z(n1124) );
NOR2_X1 U823 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U824 ( .A1(n1115), .A2(G472), .ZN(n1126) );
NOR2_X1 U825 ( .A1(n1111), .A2(n1130), .ZN(G54) );
XOR2_X1 U826 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U827 ( .A(n1133), .B(KEYINPUT17), .Z(n1132) );
NAND2_X1 U828 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U829 ( .A(KEYINPUT53), .B(KEYINPUT11), .Z(n1135) );
XNOR2_X1 U830 ( .A(G140), .B(n1136), .ZN(n1134) );
NAND2_X1 U831 ( .A1(n1115), .A2(G469), .ZN(n1131) );
NOR2_X1 U832 ( .A1(n1137), .A2(n1138), .ZN(G51) );
XNOR2_X1 U833 ( .A(n1111), .B(KEYINPUT24), .ZN(n1138) );
NOR2_X1 U834 ( .A1(n1073), .A2(G952), .ZN(n1111) );
NOR2_X1 U835 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
XOR2_X1 U836 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U837 ( .A1(n1115), .A2(n1060), .ZN(n1142) );
NOR2_X1 U838 ( .A1(n1143), .A2(n1042), .ZN(n1115) );
NOR2_X1 U839 ( .A1(n1081), .A2(n1110), .ZN(n1042) );
NAND4_X1 U840 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1110) );
NOR4_X1 U841 ( .A1(n1122), .A2(n998), .A3(n1148), .A4(n1149), .ZN(n1147) );
NOR2_X1 U842 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NOR2_X1 U844 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NOR2_X1 U845 ( .A1(n1040), .A2(n1156), .ZN(n1155) );
NOR3_X1 U846 ( .A1(n1157), .A2(n1158), .A3(n1020), .ZN(n1154) );
NAND3_X1 U847 ( .A1(n1159), .A2(n1151), .A3(n1160), .ZN(n1157) );
INV_X1 U848 ( .A(KEYINPUT55), .ZN(n1151) );
AND3_X1 U849 ( .A1(n1038), .A2(n1025), .A3(n1161), .ZN(n998) );
AND3_X1 U850 ( .A1(n1161), .A2(n1025), .A3(n1037), .ZN(n1122) );
NOR2_X1 U851 ( .A1(n1162), .A2(n1163), .ZN(n1146) );
NAND4_X1 U852 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1081) );
NOR4_X1 U853 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NAND2_X1 U854 ( .A1(n1172), .A2(n1173), .ZN(n1166) );
INV_X1 U855 ( .A(KEYINPUT38), .ZN(n1173) );
NAND3_X1 U856 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1165) );
NAND2_X1 U857 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
OR2_X1 U858 ( .A1(n1153), .A2(KEYINPUT19), .ZN(n1177) );
NAND3_X1 U859 ( .A1(n1179), .A2(n1180), .A3(n1037), .ZN(n1174) );
NAND2_X1 U860 ( .A1(KEYINPUT19), .A2(n1023), .ZN(n1179) );
NAND2_X1 U861 ( .A1(n1011), .A2(n1181), .ZN(n1164) );
NAND2_X1 U862 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND3_X1 U863 ( .A1(n1184), .A2(n1158), .A3(KEYINPUT38), .ZN(n1183) );
XOR2_X1 U864 ( .A(n1185), .B(KEYINPUT31), .Z(n1182) );
NAND2_X1 U865 ( .A1(KEYINPUT0), .A2(n1186), .ZN(n1141) );
NOR2_X1 U866 ( .A1(KEYINPUT0), .A2(n1186), .ZN(n1139) );
XNOR2_X1 U867 ( .A(n1187), .B(n1188), .ZN(n1186) );
XNOR2_X1 U868 ( .A(n1101), .B(n1189), .ZN(n1188) );
XOR2_X1 U869 ( .A(n1190), .B(n1106), .Z(n1187) );
NAND2_X1 U870 ( .A1(KEYINPUT41), .A2(n1191), .ZN(n1190) );
INV_X1 U871 ( .A(n1100), .ZN(n1191) );
XOR2_X1 U872 ( .A(G146), .B(n1171), .Z(G48) );
AND4_X1 U873 ( .A1(n1037), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1171) );
INV_X1 U874 ( .A(n1178), .ZN(n1037) );
XNOR2_X1 U875 ( .A(G143), .B(n1195), .ZN(G45) );
NAND2_X1 U876 ( .A1(KEYINPUT61), .A2(n1170), .ZN(n1195) );
AND3_X1 U877 ( .A1(n1023), .A2(n1193), .A3(n1196), .ZN(n1170) );
NOR3_X1 U878 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
XNOR2_X1 U879 ( .A(G140), .B(n1200), .ZN(G42) );
NAND3_X1 U880 ( .A1(n1201), .A2(n1032), .A3(n1202), .ZN(n1200) );
NOR3_X1 U881 ( .A1(n1203), .A2(n1014), .A3(n1013), .ZN(n1202) );
XNOR2_X1 U882 ( .A(n1198), .B(KEYINPUT16), .ZN(n1203) );
INV_X1 U883 ( .A(n1158), .ZN(n1032) );
NAND3_X1 U884 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(G39) );
NAND2_X1 U885 ( .A1(n1169), .A2(n1097), .ZN(n1206) );
NAND2_X1 U886 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U887 ( .A(KEYINPUT23), .ZN(n1208) );
NAND2_X1 U888 ( .A1(n1209), .A2(G137), .ZN(n1207) );
XNOR2_X1 U889 ( .A(n1210), .B(n1169), .ZN(n1209) );
NAND2_X1 U890 ( .A1(KEYINPUT23), .A2(n1211), .ZN(n1204) );
NAND2_X1 U891 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND3_X1 U892 ( .A1(G137), .A2(n1214), .A3(n1215), .ZN(n1213) );
INV_X1 U893 ( .A(n1210), .ZN(n1214) );
NAND2_X1 U894 ( .A1(n1210), .A2(n1169), .ZN(n1212) );
INV_X1 U895 ( .A(n1215), .ZN(n1169) );
NAND3_X1 U896 ( .A1(n1216), .A2(n1176), .A3(n1192), .ZN(n1215) );
XOR2_X1 U897 ( .A(KEYINPUT21), .B(KEYINPUT1), .Z(n1210) );
XNOR2_X1 U898 ( .A(n1217), .B(n1168), .ZN(G36) );
NOR3_X1 U899 ( .A1(n1218), .A2(n1040), .A3(n1153), .ZN(n1168) );
XOR2_X1 U900 ( .A(G131), .B(n1219), .Z(G33) );
NOR3_X1 U901 ( .A1(n1178), .A2(n1218), .A3(n1153), .ZN(n1219) );
INV_X1 U902 ( .A(n1176), .ZN(n1218) );
NOR4_X1 U903 ( .A1(n1158), .A2(n1013), .A3(n1198), .A4(n1014), .ZN(n1176) );
INV_X1 U904 ( .A(n1012), .ZN(n1014) );
INV_X1 U905 ( .A(n1194), .ZN(n1198) );
XOR2_X1 U906 ( .A(G128), .B(n1172), .Z(G30) );
AND2_X1 U907 ( .A1(n1184), .A2(n1193), .ZN(n1172) );
AND3_X1 U908 ( .A1(n1038), .A2(n1194), .A3(n1192), .ZN(n1184) );
XNOR2_X1 U909 ( .A(G101), .B(n1150), .ZN(G3) );
NAND3_X1 U910 ( .A1(n1023), .A2(n1161), .A3(n1216), .ZN(n1150) );
INV_X1 U911 ( .A(n1153), .ZN(n1023) );
XOR2_X1 U912 ( .A(n1220), .B(n1221), .Z(G27) );
XNOR2_X1 U913 ( .A(KEYINPUT42), .B(n1101), .ZN(n1221) );
NOR2_X1 U914 ( .A1(n1160), .A2(n1185), .ZN(n1220) );
NAND3_X1 U915 ( .A1(n1201), .A2(n1194), .A3(n1222), .ZN(n1185) );
NAND2_X1 U916 ( .A1(n1021), .A2(n1223), .ZN(n1194) );
NAND4_X1 U917 ( .A1(G902), .A2(G953), .A3(n1224), .A4(n1075), .ZN(n1223) );
INV_X1 U918 ( .A(G900), .ZN(n1075) );
NOR2_X1 U919 ( .A1(n1180), .A2(n1178), .ZN(n1201) );
INV_X1 U920 ( .A(n1024), .ZN(n1180) );
XNOR2_X1 U921 ( .A(G122), .B(n1144), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1225), .A2(n1025), .A3(n1226), .A4(n1227), .ZN(n1144) );
NOR2_X1 U923 ( .A1(n1228), .A2(n1229), .ZN(n1025) );
XNOR2_X1 U924 ( .A(G119), .B(n1145), .ZN(G21) );
NAND3_X1 U925 ( .A1(n1192), .A2(n1216), .A3(n1225), .ZN(n1145) );
INV_X1 U926 ( .A(n1156), .ZN(n1225) );
AND2_X1 U927 ( .A1(n1229), .A2(n1228), .ZN(n1192) );
XNOR2_X1 U928 ( .A(G116), .B(n1230), .ZN(G18) );
NAND4_X1 U929 ( .A1(n1231), .A2(n1159), .A3(n1038), .A4(n1232), .ZN(n1230) );
NOR2_X1 U930 ( .A1(n1153), .A2(n1019), .ZN(n1232) );
INV_X1 U931 ( .A(n1222), .ZN(n1019) );
INV_X1 U932 ( .A(n1040), .ZN(n1038) );
NAND2_X1 U933 ( .A1(n1044), .A2(n1227), .ZN(n1040) );
XNOR2_X1 U934 ( .A(KEYINPUT62), .B(n1160), .ZN(n1231) );
XOR2_X1 U935 ( .A(n1233), .B(n1163), .Z(G15) );
NOR3_X1 U936 ( .A1(n1178), .A2(n1153), .A3(n1156), .ZN(n1163) );
NAND3_X1 U937 ( .A1(n1011), .A2(n1159), .A3(n1222), .ZN(n1156) );
NOR2_X1 U938 ( .A1(n1034), .A2(n1234), .ZN(n1222) );
INV_X1 U939 ( .A(n1160), .ZN(n1011) );
NAND2_X1 U940 ( .A1(n1058), .A2(n1228), .ZN(n1153) );
NAND2_X1 U941 ( .A1(n1199), .A2(n1235), .ZN(n1178) );
XNOR2_X1 U942 ( .A(KEYINPUT27), .B(n1197), .ZN(n1235) );
INV_X1 U943 ( .A(n1226), .ZN(n1197) );
XNOR2_X1 U944 ( .A(n1044), .B(KEYINPUT33), .ZN(n1226) );
XNOR2_X1 U945 ( .A(G113), .B(KEYINPUT57), .ZN(n1233) );
XOR2_X1 U946 ( .A(G110), .B(n1162), .Z(G12) );
AND3_X1 U947 ( .A1(n1216), .A2(n1161), .A3(n1024), .ZN(n1162) );
NOR2_X1 U948 ( .A1(n1228), .A2(n1058), .ZN(n1024) );
INV_X1 U949 ( .A(n1229), .ZN(n1058) );
NAND3_X1 U950 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1229) );
NAND2_X1 U951 ( .A1(n1239), .A2(n1114), .ZN(n1238) );
OR3_X1 U952 ( .A1(n1114), .A2(n1239), .A3(G902), .ZN(n1237) );
NOR2_X1 U953 ( .A1(n1240), .A2(G234), .ZN(n1239) );
INV_X1 U954 ( .A(G217), .ZN(n1240) );
XNOR2_X1 U955 ( .A(n1241), .B(n1242), .ZN(n1114) );
XOR2_X1 U956 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U957 ( .A(n1097), .B(G125), .ZN(n1244) );
INV_X1 U958 ( .A(G137), .ZN(n1097) );
XNOR2_X1 U959 ( .A(KEYINPUT22), .B(n1086), .ZN(n1243) );
XOR2_X1 U960 ( .A(n1245), .B(n1246), .Z(n1241) );
XNOR2_X1 U961 ( .A(n1247), .B(n1248), .ZN(n1245) );
AND3_X1 U962 ( .A1(G221), .A2(n1073), .A3(G234), .ZN(n1248) );
NAND2_X1 U963 ( .A1(G217), .A2(G902), .ZN(n1236) );
NAND3_X1 U964 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1228) );
NAND2_X1 U965 ( .A1(G472), .A2(n1069), .ZN(n1251) );
NAND2_X1 U966 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
INV_X1 U967 ( .A(KEYINPUT60), .ZN(n1253) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1054), .ZN(n1252) );
XNOR2_X1 U969 ( .A(n1053), .B(KEYINPUT20), .ZN(n1254) );
NAND2_X1 U970 ( .A1(KEYINPUT60), .A2(n1255), .ZN(n1249) );
NAND2_X1 U971 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
OR2_X1 U972 ( .A1(n1053), .A2(KEYINPUT20), .ZN(n1257) );
NAND3_X1 U973 ( .A1(n1053), .A2(n1054), .A3(KEYINPUT20), .ZN(n1256) );
INV_X1 U974 ( .A(G472), .ZN(n1054) );
INV_X1 U975 ( .A(n1069), .ZN(n1053) );
NAND2_X1 U976 ( .A1(n1258), .A2(n1143), .ZN(n1069) );
XOR2_X1 U977 ( .A(n1259), .B(n1260), .Z(n1258) );
NOR2_X1 U978 ( .A1(KEYINPUT51), .A2(n1125), .ZN(n1260) );
XOR2_X1 U979 ( .A(n1261), .B(G101), .Z(n1125) );
NAND2_X1 U980 ( .A1(n1262), .A2(G210), .ZN(n1261) );
NOR2_X1 U981 ( .A1(n1129), .A2(n1263), .ZN(n1259) );
XNOR2_X1 U982 ( .A(n1128), .B(KEYINPUT30), .ZN(n1263) );
NOR2_X1 U983 ( .A1(n1264), .A2(n1265), .ZN(n1128) );
AND2_X1 U984 ( .A1(n1265), .A2(n1264), .ZN(n1129) );
XNOR2_X1 U985 ( .A(n1266), .B(n1267), .ZN(n1264) );
XNOR2_X1 U986 ( .A(G113), .B(n1268), .ZN(n1266) );
AND2_X1 U987 ( .A1(n1193), .A2(n1159), .ZN(n1161) );
NAND2_X1 U988 ( .A1(n1021), .A2(n1269), .ZN(n1159) );
NAND3_X1 U989 ( .A1(n1108), .A2(n1224), .A3(G902), .ZN(n1269) );
NOR2_X1 U990 ( .A1(n1073), .A2(G898), .ZN(n1108) );
NAND3_X1 U991 ( .A1(n1041), .A2(n1224), .A3(G952), .ZN(n1021) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1224) );
INV_X1 U993 ( .A(n1043), .ZN(n1041) );
XOR2_X1 U994 ( .A(G953), .B(KEYINPUT9), .Z(n1043) );
NOR2_X1 U995 ( .A1(n1158), .A2(n1160), .ZN(n1193) );
NAND2_X1 U996 ( .A1(n1013), .A2(n1270), .ZN(n1160) );
XNOR2_X1 U997 ( .A(KEYINPUT59), .B(n1012), .ZN(n1270) );
NAND2_X1 U998 ( .A1(G214), .A2(n1271), .ZN(n1012) );
XNOR2_X1 U999 ( .A(n1060), .B(n1272), .ZN(n1013) );
NOR2_X1 U1000 ( .A1(KEYINPUT4), .A2(n1273), .ZN(n1272) );
XOR2_X1 U1001 ( .A(n1062), .B(KEYINPUT25), .Z(n1273) );
NAND2_X1 U1002 ( .A1(n1274), .A2(n1143), .ZN(n1062) );
XOR2_X1 U1003 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U1004 ( .A(n1106), .B(n1100), .ZN(n1276) );
XOR2_X1 U1005 ( .A(G143), .B(n1246), .Z(n1100) );
XNOR2_X1 U1006 ( .A(n1277), .B(n1278), .ZN(n1106) );
XOR2_X1 U1007 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U1008 ( .A(G101), .B(n1281), .ZN(n1280) );
NAND2_X1 U1009 ( .A1(KEYINPUT6), .A2(n1267), .ZN(n1281) );
XOR2_X1 U1010 ( .A(G116), .B(KEYINPUT18), .Z(n1267) );
NOR2_X1 U1011 ( .A1(G113), .A2(KEYINPUT48), .ZN(n1279) );
XOR2_X1 U1012 ( .A(n1282), .B(n1283), .Z(n1277) );
XOR2_X1 U1013 ( .A(n1284), .B(n1247), .Z(n1282) );
XOR2_X1 U1014 ( .A(G110), .B(n1268), .Z(n1247) );
XOR2_X1 U1015 ( .A(G119), .B(KEYINPUT50), .Z(n1268) );
NAND2_X1 U1016 ( .A1(KEYINPUT8), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1017 ( .A(n1286), .B(n1287), .ZN(n1275) );
NAND2_X1 U1018 ( .A1(KEYINPUT52), .A2(n1101), .ZN(n1287) );
INV_X1 U1019 ( .A(G125), .ZN(n1101) );
NAND2_X1 U1020 ( .A1(KEYINPUT26), .A2(n1189), .ZN(n1286) );
AND2_X1 U1021 ( .A1(G224), .A2(n1073), .ZN(n1189) );
AND2_X1 U1022 ( .A1(G210), .A2(n1271), .ZN(n1060) );
NAND2_X1 U1023 ( .A1(n1288), .A2(n1143), .ZN(n1271) );
INV_X1 U1024 ( .A(G237), .ZN(n1288) );
NAND2_X1 U1025 ( .A1(n1289), .A2(n1034), .ZN(n1158) );
XNOR2_X1 U1026 ( .A(n1290), .B(G469), .ZN(n1034) );
NAND2_X1 U1027 ( .A1(n1291), .A2(n1143), .ZN(n1290) );
XNOR2_X1 U1028 ( .A(n1292), .B(n1136), .ZN(n1291) );
XNOR2_X1 U1029 ( .A(n1293), .B(n1294), .ZN(n1136) );
XNOR2_X1 U1030 ( .A(n1265), .B(n1283), .ZN(n1294) );
XNOR2_X1 U1031 ( .A(G104), .B(n1000), .ZN(n1283) );
XOR2_X1 U1032 ( .A(n1295), .B(n1296), .Z(n1265) );
XOR2_X1 U1033 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U1034 ( .A(KEYINPUT35), .B(KEYINPUT54), .ZN(n1298) );
NAND2_X1 U1035 ( .A1(n1299), .A2(n1091), .ZN(n1297) );
NAND2_X1 U1036 ( .A1(G137), .A2(n1217), .ZN(n1091) );
XNOR2_X1 U1037 ( .A(n1094), .B(KEYINPUT47), .ZN(n1299) );
NOR2_X1 U1038 ( .A1(n1217), .A2(G137), .ZN(n1094) );
INV_X1 U1039 ( .A(G134), .ZN(n1217) );
XNOR2_X1 U1040 ( .A(n1246), .B(n1300), .ZN(n1295) );
XOR2_X1 U1041 ( .A(G128), .B(G146), .Z(n1246) );
XOR2_X1 U1042 ( .A(n1301), .B(n1302), .Z(n1293) );
NOR2_X1 U1043 ( .A1(G101), .A2(KEYINPUT63), .ZN(n1302) );
XNOR2_X1 U1044 ( .A(G110), .B(n1303), .ZN(n1301) );
NOR2_X1 U1045 ( .A1(G953), .A2(n1074), .ZN(n1303) );
INV_X1 U1046 ( .A(G227), .ZN(n1074) );
NAND2_X1 U1047 ( .A1(KEYINPUT7), .A2(n1086), .ZN(n1292) );
INV_X1 U1048 ( .A(G140), .ZN(n1086) );
INV_X1 U1049 ( .A(n1234), .ZN(n1289) );
XOR2_X1 U1050 ( .A(n1068), .B(KEYINPUT14), .Z(n1234) );
INV_X1 U1051 ( .A(n1033), .ZN(n1068) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1304), .ZN(n1033) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1143), .ZN(n1304) );
INV_X1 U1054 ( .A(n1020), .ZN(n1216) );
NAND2_X1 U1055 ( .A1(n1199), .A2(n1044), .ZN(n1020) );
XOR2_X1 U1056 ( .A(n1305), .B(G475), .Z(n1044) );
NAND2_X1 U1057 ( .A1(n1121), .A2(n1143), .ZN(n1305) );
XOR2_X1 U1058 ( .A(n1306), .B(n1307), .Z(n1121) );
XOR2_X1 U1059 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1060 ( .A(n1310), .B(n1300), .Z(n1309) );
XOR2_X1 U1061 ( .A(G131), .B(G143), .Z(n1300) );
NAND2_X1 U1062 ( .A1(KEYINPUT49), .A2(G125), .ZN(n1310) );
XOR2_X1 U1063 ( .A(n1311), .B(n1312), .Z(n1308) );
NOR2_X1 U1064 ( .A1(KEYINPUT36), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1065 ( .A(G113), .B(n1285), .Z(n1313) );
NAND2_X1 U1066 ( .A1(n1262), .A2(G214), .ZN(n1311) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1262) );
XOR2_X1 U1068 ( .A(n1314), .B(n1315), .Z(n1306) );
XOR2_X1 U1069 ( .A(KEYINPUT56), .B(G146), .Z(n1315) );
XNOR2_X1 U1070 ( .A(G104), .B(G140), .ZN(n1314) );
INV_X1 U1071 ( .A(n1227), .ZN(n1199) );
XNOR2_X1 U1072 ( .A(n1316), .B(G478), .ZN(n1227) );
NAND2_X1 U1073 ( .A1(KEYINPUT13), .A2(n1051), .ZN(n1316) );
AND2_X1 U1074 ( .A1(n1143), .A2(n1117), .ZN(n1051) );
NAND2_X1 U1075 ( .A1(n1317), .A2(n1318), .ZN(n1117) );
NAND2_X1 U1076 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1077 ( .A(n1321), .B(KEYINPUT32), .Z(n1317) );
NAND2_X1 U1078 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
INV_X1 U1079 ( .A(n1320), .ZN(n1323) );
NAND3_X1 U1080 ( .A1(G234), .A2(n1073), .A3(G217), .ZN(n1320) );
INV_X1 U1081 ( .A(G953), .ZN(n1073) );
XOR2_X1 U1082 ( .A(n1319), .B(KEYINPUT40), .Z(n1322) );
XOR2_X1 U1083 ( .A(n1324), .B(n1325), .Z(n1319) );
XNOR2_X1 U1084 ( .A(n1326), .B(G134), .ZN(n1325) );
INV_X1 U1085 ( .A(G143), .ZN(n1326) );
XOR2_X1 U1086 ( .A(n1327), .B(G128), .Z(n1324) );
NAND2_X1 U1087 ( .A1(KEYINPUT3), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1088 ( .A(n1285), .B(n1329), .Z(n1328) );
XOR2_X1 U1089 ( .A(G116), .B(n1330), .Z(n1329) );
NOR2_X1 U1090 ( .A1(KEYINPUT34), .A2(n1000), .ZN(n1330) );
INV_X1 U1091 ( .A(G107), .ZN(n1000) );
XOR2_X1 U1092 ( .A(G122), .B(KEYINPUT58), .Z(n1285) );
INV_X1 U1093 ( .A(G902), .ZN(n1143) );
endmodule


