//Key = 1000111000010101001011000011111101101011000111000110001110000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300;

NAND2_X1 U706 ( .A1(n983), .A2(n984), .ZN(G9) );
NAND3_X1 U707 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
XOR2_X1 U708 ( .A(n988), .B(KEYINPUT17), .Z(n983) );
NAND2_X1 U709 ( .A1(G107), .A2(n989), .ZN(n988) );
NAND2_X1 U710 ( .A1(n987), .A2(n985), .ZN(n989) );
INV_X1 U711 ( .A(n990), .ZN(n987) );
NOR2_X1 U712 ( .A1(n991), .A2(n992), .ZN(G75) );
NOR4_X1 U713 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n992) );
NOR2_X1 U714 ( .A1(n997), .A2(n998), .ZN(n996) );
XOR2_X1 U715 ( .A(n999), .B(KEYINPUT7), .Z(n997) );
NOR3_X1 U716 ( .A1(n1000), .A2(n999), .A3(n1001), .ZN(n995) );
NAND4_X1 U717 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n999) );
NAND3_X1 U718 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n993) );
NAND3_X1 U719 ( .A1(n1009), .A2(n1010), .A3(n1002), .ZN(n1008) );
INV_X1 U720 ( .A(n1011), .ZN(n1002) );
NAND2_X1 U721 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NAND3_X1 U722 ( .A1(n1005), .A2(n1014), .A3(n1003), .ZN(n1013) );
INV_X1 U723 ( .A(n1015), .ZN(n1014) );
NAND2_X1 U724 ( .A1(n1004), .A2(n1016), .ZN(n1012) );
NAND2_X1 U725 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U726 ( .A1(n1005), .A2(n1019), .ZN(n1018) );
NAND2_X1 U727 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U728 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
INV_X1 U729 ( .A(n1024), .ZN(n1020) );
NAND2_X1 U730 ( .A1(n1003), .A2(n1025), .ZN(n1017) );
OR2_X1 U731 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR3_X1 U732 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n991) );
INV_X1 U733 ( .A(n1006), .ZN(n1028) );
NAND4_X1 U734 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1006) );
NOR4_X1 U735 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XOR2_X1 U736 ( .A(n1037), .B(n1038), .Z(n1036) );
XOR2_X1 U737 ( .A(KEYINPUT62), .B(n1039), .Z(n1035) );
XOR2_X1 U738 ( .A(n1040), .B(n1041), .Z(n1034) );
NAND2_X1 U739 ( .A1(KEYINPUT11), .A2(n1042), .ZN(n1041) );
XOR2_X1 U740 ( .A(n1043), .B(n1044), .Z(n1033) );
NAND2_X1 U741 ( .A1(KEYINPUT26), .A2(G478), .ZN(n1044) );
NOR2_X1 U742 ( .A1(n1022), .A2(n1045), .ZN(n1031) );
XNOR2_X1 U743 ( .A(n1046), .B(n1047), .ZN(n1030) );
NOR2_X1 U744 ( .A1(n1048), .A2(KEYINPUT46), .ZN(n1047) );
XOR2_X1 U745 ( .A(n1049), .B(n1050), .Z(G72) );
NOR2_X1 U746 ( .A1(n1051), .A2(KEYINPUT40), .ZN(n1050) );
NOR2_X1 U747 ( .A1(G953), .A2(n1052), .ZN(n1051) );
XOR2_X1 U748 ( .A(n1053), .B(n1054), .Z(n1049) );
NOR2_X1 U749 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U750 ( .A(n1057), .ZN(n1056) );
NOR2_X1 U751 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NAND2_X1 U752 ( .A1(n1060), .A2(n1061), .ZN(n1053) );
NAND2_X1 U753 ( .A1(n1062), .A2(n1059), .ZN(n1061) );
XOR2_X1 U754 ( .A(n1063), .B(n1064), .Z(n1060) );
XOR2_X1 U755 ( .A(n1065), .B(n1066), .Z(n1064) );
NOR2_X1 U756 ( .A1(KEYINPUT9), .A2(n1067), .ZN(n1066) );
XNOR2_X1 U757 ( .A(G140), .B(G125), .ZN(n1067) );
XOR2_X1 U758 ( .A(n1068), .B(n1069), .Z(n1063) );
NOR2_X1 U759 ( .A1(KEYINPUT53), .A2(n1070), .ZN(n1069) );
XNOR2_X1 U760 ( .A(n1071), .B(KEYINPUT35), .ZN(n1070) );
XNOR2_X1 U761 ( .A(KEYINPUT15), .B(KEYINPUT10), .ZN(n1068) );
XOR2_X1 U762 ( .A(n1072), .B(n1073), .Z(G69) );
NOR2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U764 ( .A(KEYINPUT12), .B(n1076), .Z(n1075) );
NOR2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
AND2_X1 U766 ( .A1(n1078), .A2(n1077), .ZN(n1074) );
AND2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XNOR2_X1 U769 ( .A(KEYINPUT49), .B(n1083), .ZN(n1082) );
XOR2_X1 U770 ( .A(KEYINPUT30), .B(G953), .Z(n1079) );
NAND3_X1 U771 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1078) );
NAND2_X1 U772 ( .A1(n1062), .A2(n1087), .ZN(n1086) );
INV_X1 U773 ( .A(n1088), .ZN(n1085) );
NAND2_X1 U774 ( .A1(n1057), .A2(n1089), .ZN(n1072) );
NAND2_X1 U775 ( .A1(G898), .A2(G224), .ZN(n1089) );
XOR2_X1 U776 ( .A(n1007), .B(KEYINPUT39), .Z(n1057) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(G66) );
NOR3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NOR4_X1 U779 ( .A1(n1095), .A2(n1096), .A3(n1038), .A4(n1097), .ZN(n1094) );
NOR2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
NOR3_X1 U781 ( .A1(n1096), .A2(n1100), .A3(n1038), .ZN(n1098) );
INV_X1 U782 ( .A(n994), .ZN(n1100) );
INV_X1 U783 ( .A(KEYINPUT36), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1101), .ZN(G63) );
XOR2_X1 U785 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U786 ( .A1(n1104), .A2(KEYINPUT1), .ZN(n1103) );
INV_X1 U787 ( .A(n1105), .ZN(n1104) );
NAND2_X1 U788 ( .A1(n1106), .A2(G478), .ZN(n1102) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1107), .ZN(G60) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U791 ( .A1(KEYINPUT51), .A2(n1110), .ZN(n1109) );
NAND2_X1 U792 ( .A1(n1106), .A2(G475), .ZN(n1108) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(G6) );
NOR2_X1 U794 ( .A1(G104), .A2(KEYINPUT23), .ZN(n1112) );
NAND3_X1 U795 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1111) );
AND3_X1 U796 ( .A1(n1005), .A2(n1116), .A3(n1024), .ZN(n1115) );
XOR2_X1 U797 ( .A(n998), .B(KEYINPUT33), .Z(n1113) );
NOR2_X1 U798 ( .A1(n1090), .A2(n1117), .ZN(G57) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U800 ( .A(KEYINPUT57), .B(n1120), .ZN(n1119) );
NOR2_X1 U801 ( .A1(KEYINPUT19), .A2(n1121), .ZN(n1120) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(n1121) );
AND2_X1 U803 ( .A1(G472), .A2(n1106), .ZN(n1122) );
INV_X1 U804 ( .A(n1097), .ZN(n1106) );
NOR2_X1 U805 ( .A1(n1090), .A2(n1124), .ZN(G54) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U807 ( .A(n1127), .B(n1071), .Z(n1126) );
XOR2_X1 U808 ( .A(n1128), .B(n1129), .Z(n1125) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U810 ( .A1(KEYINPUT22), .A2(n1065), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1040), .A2(n1097), .ZN(n1130) );
NAND3_X1 U812 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
OR3_X1 U814 ( .A1(n1136), .A2(n1135), .A3(n1137), .ZN(n1133) );
INV_X1 U815 ( .A(KEYINPUT56), .ZN(n1136) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U817 ( .A1(n1139), .A2(KEYINPUT56), .ZN(n1138) );
XNOR2_X1 U818 ( .A(n1135), .B(KEYINPUT61), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1140), .B(KEYINPUT29), .Z(n1135) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(G51) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U822 ( .A(n1071), .B(n1145), .ZN(n1144) );
XOR2_X1 U823 ( .A(G125), .B(n1146), .Z(n1143) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1097), .ZN(n1146) );
NAND2_X1 U825 ( .A1(G902), .A2(n994), .ZN(n1097) );
NAND3_X1 U826 ( .A1(n1081), .A2(n1083), .A3(n1052), .ZN(n994) );
AND4_X1 U827 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1052) );
NOR4_X1 U828 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1015), .A2(n1156), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n998), .A2(n1157), .ZN(n1154) );
NOR3_X1 U831 ( .A1(n1114), .A2(n1158), .A3(n1159), .ZN(n1153) );
INV_X1 U832 ( .A(KEYINPUT48), .ZN(n1159) );
NOR2_X1 U833 ( .A1(n1160), .A2(n1161), .ZN(n1152) );
NOR2_X1 U834 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
NOR2_X1 U835 ( .A1(KEYINPUT48), .A2(n1158), .ZN(n1163) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
XOR2_X1 U837 ( .A(KEYINPUT31), .B(n1166), .Z(n1165) );
AND4_X1 U838 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1081) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1015), .A2(n990), .ZN(n1172) );
NAND2_X1 U841 ( .A1(n1173), .A2(n1005), .ZN(n990) );
NOR2_X1 U842 ( .A1(n1114), .A2(n985), .ZN(n1015) );
NOR2_X1 U843 ( .A1(n1174), .A2(n998), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XNOR2_X1 U845 ( .A(n1090), .B(KEYINPUT18), .ZN(n1141) );
NOR2_X1 U846 ( .A1(n1007), .A2(G952), .ZN(n1090) );
XNOR2_X1 U847 ( .A(G146), .B(n1177), .ZN(G48) );
NAND2_X1 U848 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XNOR2_X1 U849 ( .A(G143), .B(n1180), .ZN(G45) );
NAND2_X1 U850 ( .A1(n1181), .A2(n1166), .ZN(n1180) );
XOR2_X1 U851 ( .A(n1157), .B(KEYINPUT44), .Z(n1181) );
NAND4_X1 U852 ( .A1(n1026), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1157) );
XNOR2_X1 U853 ( .A(G140), .B(n1150), .ZN(G42) );
NAND4_X1 U854 ( .A1(n1114), .A2(n1027), .A3(n1009), .A4(n1182), .ZN(n1150) );
INV_X1 U855 ( .A(n1161), .ZN(n1114) );
XNOR2_X1 U856 ( .A(G137), .B(n1148), .ZN(G39) );
NAND3_X1 U857 ( .A1(n1004), .A2(n1179), .A3(n1009), .ZN(n1148) );
XOR2_X1 U858 ( .A(n1185), .B(n1186), .Z(G36) );
XOR2_X1 U859 ( .A(n1187), .B(KEYINPUT47), .Z(n1186) );
NAND2_X1 U860 ( .A1(n1188), .A2(n985), .ZN(n1185) );
XNOR2_X1 U861 ( .A(G131), .B(n1189), .ZN(G33) );
NAND2_X1 U862 ( .A1(n1190), .A2(n1188), .ZN(n1189) );
INV_X1 U863 ( .A(n1156), .ZN(n1188) );
NAND3_X1 U864 ( .A1(n1009), .A2(n1182), .A3(n1026), .ZN(n1156) );
NOR2_X1 U865 ( .A1(n1001), .A2(n1045), .ZN(n1009) );
INV_X1 U866 ( .A(n1000), .ZN(n1045) );
XOR2_X1 U867 ( .A(n1161), .B(KEYINPUT0), .Z(n1190) );
XNOR2_X1 U868 ( .A(G128), .B(n1149), .ZN(G30) );
NAND3_X1 U869 ( .A1(n985), .A2(n1166), .A3(n1179), .ZN(n1149) );
INV_X1 U870 ( .A(n1164), .ZN(n1179) );
NAND3_X1 U871 ( .A1(n1191), .A2(n1039), .A3(n1182), .ZN(n1164) );
AND2_X1 U872 ( .A1(n1024), .A2(n1192), .ZN(n1182) );
XOR2_X1 U873 ( .A(n1169), .B(n1193), .Z(G3) );
XOR2_X1 U874 ( .A(n1194), .B(KEYINPUT2), .Z(n1193) );
NAND3_X1 U875 ( .A1(n1004), .A2(n1173), .A3(n1026), .ZN(n1169) );
XOR2_X1 U876 ( .A(G125), .B(n1195), .Z(G27) );
NOR2_X1 U877 ( .A1(n1161), .A2(n1158), .ZN(n1195) );
NAND4_X1 U878 ( .A1(n1003), .A2(n1027), .A3(n1166), .A4(n1192), .ZN(n1158) );
NAND2_X1 U879 ( .A1(n1196), .A2(n1011), .ZN(n1192) );
XOR2_X1 U880 ( .A(KEYINPUT50), .B(n1197), .Z(n1196) );
AND4_X1 U881 ( .A1(n1059), .A2(n1198), .A3(G902), .A4(n1062), .ZN(n1197) );
INV_X1 U882 ( .A(G900), .ZN(n1059) );
XOR2_X1 U883 ( .A(n1199), .B(n1168), .Z(G24) );
NAND3_X1 U884 ( .A1(n1200), .A2(n1005), .A3(n1201), .ZN(n1168) );
NOR3_X1 U885 ( .A1(n998), .A2(n1029), .A3(n1202), .ZN(n1201) );
NOR2_X1 U886 ( .A1(n1039), .A2(n1191), .ZN(n1005) );
XOR2_X1 U887 ( .A(n1203), .B(n1204), .Z(G21) );
NAND2_X1 U888 ( .A1(n1205), .A2(n1175), .ZN(n1204) );
AND4_X1 U889 ( .A1(n1200), .A2(n1004), .A3(n1191), .A4(n1039), .ZN(n1175) );
INV_X1 U890 ( .A(n1206), .ZN(n1039) );
XOR2_X1 U891 ( .A(n998), .B(KEYINPUT6), .Z(n1205) );
XOR2_X1 U892 ( .A(G116), .B(n1207), .Z(G18) );
NOR2_X1 U893 ( .A1(n1208), .A2(n998), .ZN(n1207) );
XNOR2_X1 U894 ( .A(n1176), .B(KEYINPUT58), .ZN(n1208) );
AND3_X1 U895 ( .A1(n1026), .A2(n985), .A3(n1200), .ZN(n1176) );
NOR2_X1 U896 ( .A1(n1184), .A2(n1202), .ZN(n985) );
XNOR2_X1 U897 ( .A(G113), .B(n1083), .ZN(G15) );
NAND3_X1 U898 ( .A1(n1200), .A2(n1026), .A3(n1178), .ZN(n1083) );
NOR2_X1 U899 ( .A1(n1161), .A2(n998), .ZN(n1178) );
NAND2_X1 U900 ( .A1(n1202), .A2(n1184), .ZN(n1161) );
NOR2_X1 U901 ( .A1(n1191), .A2(n1206), .ZN(n1026) );
AND2_X1 U902 ( .A1(n1003), .A2(n1116), .ZN(n1200) );
NOR2_X1 U903 ( .A1(n1209), .A2(n1022), .ZN(n1003) );
NAND3_X1 U904 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(G12) );
OR2_X1 U905 ( .A1(G110), .A2(KEYINPUT5), .ZN(n1212) );
NAND3_X1 U906 ( .A1(KEYINPUT5), .A2(G110), .A3(n1167), .ZN(n1211) );
NAND2_X1 U907 ( .A1(n1213), .A2(n1214), .ZN(n1210) );
NAND2_X1 U908 ( .A1(KEYINPUT5), .A2(n1215), .ZN(n1214) );
XOR2_X1 U909 ( .A(KEYINPUT3), .B(G110), .Z(n1215) );
INV_X1 U910 ( .A(n1167), .ZN(n1213) );
NAND3_X1 U911 ( .A1(n1004), .A2(n1173), .A3(n1027), .ZN(n1167) );
AND2_X1 U912 ( .A1(n1191), .A2(n1206), .ZN(n1027) );
XOR2_X1 U913 ( .A(n1216), .B(G472), .Z(n1206) );
NAND2_X1 U914 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U915 ( .A(n1219), .B(n1220), .Z(n1217) );
INV_X1 U916 ( .A(n1118), .ZN(n1220) );
XOR2_X1 U917 ( .A(n1221), .B(G101), .Z(n1118) );
NAND3_X1 U918 ( .A1(n1222), .A2(n1007), .A3(G210), .ZN(n1221) );
XNOR2_X1 U919 ( .A(n1123), .B(KEYINPUT4), .ZN(n1219) );
XNOR2_X1 U920 ( .A(n1223), .B(n1224), .ZN(n1123) );
XNOR2_X1 U921 ( .A(n1225), .B(n1038), .ZN(n1191) );
NAND2_X1 U922 ( .A1(G217), .A2(n1226), .ZN(n1038) );
NAND2_X1 U923 ( .A1(KEYINPUT21), .A2(n1227), .ZN(n1225) );
XOR2_X1 U924 ( .A(KEYINPUT55), .B(n1092), .Z(n1227) );
INV_X1 U925 ( .A(n1037), .ZN(n1092) );
NAND2_X1 U926 ( .A1(n1095), .A2(n1218), .ZN(n1037) );
INV_X1 U927 ( .A(n1099), .ZN(n1095) );
XOR2_X1 U928 ( .A(n1228), .B(KEYINPUT63), .Z(n1099) );
XOR2_X1 U929 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U930 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U931 ( .A(G128), .B(G125), .Z(n1232) );
XOR2_X1 U932 ( .A(KEYINPUT32), .B(G137), .Z(n1231) );
XOR2_X1 U933 ( .A(n1233), .B(n1234), .Z(n1229) );
XOR2_X1 U934 ( .A(n1235), .B(n1140), .Z(n1234) );
XNOR2_X1 U935 ( .A(n1236), .B(G140), .ZN(n1140) );
NOR2_X1 U936 ( .A1(G146), .A2(KEYINPUT60), .ZN(n1235) );
XOR2_X1 U937 ( .A(n1237), .B(G119), .Z(n1233) );
NAND3_X1 U938 ( .A1(G234), .A2(n1007), .A3(G221), .ZN(n1237) );
AND3_X1 U939 ( .A1(n1166), .A2(n1116), .A3(n1024), .ZN(n1173) );
NOR2_X1 U940 ( .A1(n1022), .A2(n1023), .ZN(n1024) );
INV_X1 U941 ( .A(n1209), .ZN(n1023) );
NAND2_X1 U942 ( .A1(n1238), .A2(n1239), .ZN(n1209) );
NAND2_X1 U943 ( .A1(KEYINPUT52), .A2(n1040), .ZN(n1239) );
XNOR2_X1 U944 ( .A(n1042), .B(n1240), .ZN(n1238) );
NOR2_X1 U945 ( .A1(KEYINPUT52), .A2(n1040), .ZN(n1240) );
INV_X1 U946 ( .A(G469), .ZN(n1040) );
AND2_X1 U947 ( .A1(n1218), .A2(n1241), .ZN(n1042) );
NAND2_X1 U948 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U949 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U950 ( .A(KEYINPUT38), .B(n1246), .Z(n1242) );
NOR2_X1 U951 ( .A1(n1245), .A2(n1244), .ZN(n1246) );
XOR2_X1 U952 ( .A(n1127), .B(n1224), .Z(n1244) );
XNOR2_X1 U953 ( .A(n1065), .B(n1071), .ZN(n1224) );
XOR2_X1 U954 ( .A(n1247), .B(n1248), .Z(n1065) );
XOR2_X1 U955 ( .A(KEYINPUT8), .B(G137), .Z(n1248) );
XOR2_X1 U956 ( .A(G131), .B(n1187), .Z(n1247) );
INV_X1 U957 ( .A(G134), .ZN(n1187) );
XNOR2_X1 U958 ( .A(n1137), .B(n1249), .ZN(n1245) );
XOR2_X1 U959 ( .A(G140), .B(n1250), .Z(n1249) );
NOR2_X1 U960 ( .A1(KEYINPUT16), .A2(G110), .ZN(n1250) );
NOR2_X1 U961 ( .A1(n1058), .A2(G953), .ZN(n1137) );
INV_X1 U962 ( .A(G227), .ZN(n1058) );
AND2_X1 U963 ( .A1(G221), .A2(n1226), .ZN(n1022) );
NAND2_X1 U964 ( .A1(G234), .A2(n1218), .ZN(n1226) );
NAND2_X1 U965 ( .A1(n1251), .A2(n1011), .ZN(n1116) );
NAND3_X1 U966 ( .A1(n1198), .A2(n1007), .A3(G952), .ZN(n1011) );
NAND4_X1 U967 ( .A1(n1062), .A2(G902), .A3(n1198), .A4(n1087), .ZN(n1251) );
INV_X1 U968 ( .A(G898), .ZN(n1087) );
NAND2_X1 U969 ( .A1(G237), .A2(G234), .ZN(n1198) );
XOR2_X1 U970 ( .A(n1007), .B(KEYINPUT43), .Z(n1062) );
INV_X1 U971 ( .A(n998), .ZN(n1166) );
NAND2_X1 U972 ( .A1(n1001), .A2(n1000), .ZN(n998) );
NAND2_X1 U973 ( .A1(n1252), .A2(G214), .ZN(n1000) );
XOR2_X1 U974 ( .A(n1253), .B(KEYINPUT37), .Z(n1252) );
XNOR2_X1 U975 ( .A(n1046), .B(n1048), .ZN(n1001) );
INV_X1 U976 ( .A(n1147), .ZN(n1048) );
NAND2_X1 U977 ( .A1(G210), .A2(n1253), .ZN(n1147) );
NAND2_X1 U978 ( .A1(n1218), .A2(n1222), .ZN(n1253) );
INV_X1 U979 ( .A(G237), .ZN(n1222) );
NAND2_X1 U980 ( .A1(n1254), .A2(n1218), .ZN(n1046) );
XOR2_X1 U981 ( .A(n1145), .B(n1255), .Z(n1254) );
XOR2_X1 U982 ( .A(KEYINPUT25), .B(n1256), .Z(n1255) );
NOR2_X1 U983 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NOR2_X1 U984 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NOR2_X1 U985 ( .A1(n1071), .A2(n1261), .ZN(n1260) );
NOR2_X1 U986 ( .A1(G125), .A2(n1262), .ZN(n1259) );
AND2_X1 U987 ( .A1(n1071), .A2(KEYINPUT24), .ZN(n1262) );
NOR4_X1 U988 ( .A1(KEYINPUT24), .A2(G125), .A3(n1261), .A4(n1071), .ZN(n1257) );
XOR2_X1 U989 ( .A(G146), .B(n1263), .Z(n1071) );
INV_X1 U990 ( .A(KEYINPUT28), .ZN(n1261) );
XOR2_X1 U991 ( .A(n1264), .B(n1265), .Z(n1145) );
NOR2_X1 U992 ( .A1(n1088), .A2(n1266), .ZN(n1265) );
XOR2_X1 U993 ( .A(n1084), .B(KEYINPUT45), .Z(n1266) );
NAND2_X1 U994 ( .A1(n1267), .A2(n1268), .ZN(n1084) );
NOR2_X1 U995 ( .A1(n1268), .A2(n1267), .ZN(n1088) );
XNOR2_X1 U996 ( .A(n1223), .B(n1127), .ZN(n1267) );
XOR2_X1 U997 ( .A(n1194), .B(n1269), .Z(n1127) );
XOR2_X1 U998 ( .A(G107), .B(G104), .Z(n1269) );
INV_X1 U999 ( .A(G101), .ZN(n1194) );
XOR2_X1 U1000 ( .A(n1270), .B(n1271), .Z(n1223) );
INV_X1 U1001 ( .A(n1272), .ZN(n1271) );
XOR2_X1 U1002 ( .A(n1203), .B(n1273), .Z(n1270) );
INV_X1 U1003 ( .A(G119), .ZN(n1203) );
XOR2_X1 U1004 ( .A(n1199), .B(n1236), .Z(n1268) );
INV_X1 U1005 ( .A(G110), .ZN(n1236) );
INV_X1 U1006 ( .A(G122), .ZN(n1199) );
NAND2_X1 U1007 ( .A1(G224), .A2(n1007), .ZN(n1264) );
NOR2_X1 U1008 ( .A1(n1183), .A2(n1184), .ZN(n1004) );
INV_X1 U1009 ( .A(n1029), .ZN(n1184) );
XOR2_X1 U1010 ( .A(n1274), .B(n1275), .Z(n1029) );
XOR2_X1 U1011 ( .A(KEYINPUT14), .B(G475), .Z(n1275) );
OR2_X1 U1012 ( .A1(n1110), .A2(G902), .ZN(n1274) );
XNOR2_X1 U1013 ( .A(n1276), .B(G122), .ZN(n1110) );
XOR2_X1 U1014 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1015 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1016 ( .A(G143), .B(G131), .Z(n1280) );
XOR2_X1 U1017 ( .A(KEYINPUT20), .B(G146), .Z(n1279) );
XOR2_X1 U1018 ( .A(n1281), .B(n1282), .Z(n1277) );
XOR2_X1 U1019 ( .A(G104), .B(n1283), .Z(n1282) );
NOR2_X1 U1020 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U1021 ( .A(n1286), .B(KEYINPUT54), .Z(n1285) );
NAND2_X1 U1022 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NOR2_X1 U1023 ( .A1(n1288), .A2(n1287), .ZN(n1284) );
XOR2_X1 U1024 ( .A(KEYINPUT32), .B(G140), .Z(n1287) );
XOR2_X1 U1025 ( .A(KEYINPUT34), .B(G125), .Z(n1288) );
XOR2_X1 U1026 ( .A(n1272), .B(n1289), .Z(n1281) );
NOR4_X1 U1027 ( .A1(KEYINPUT59), .A2(G953), .A3(G237), .A4(n1290), .ZN(n1289) );
INV_X1 U1028 ( .A(G214), .ZN(n1290) );
XNOR2_X1 U1029 ( .A(G113), .B(KEYINPUT13), .ZN(n1272) );
INV_X1 U1030 ( .A(n1202), .ZN(n1183) );
XOR2_X1 U1031 ( .A(n1043), .B(G478), .Z(n1202) );
NAND2_X1 U1032 ( .A1(n1218), .A2(n1105), .ZN(n1043) );
NAND2_X1 U1033 ( .A1(n1291), .A2(n1292), .ZN(n1105) );
NAND4_X1 U1034 ( .A1(G217), .A2(G234), .A3(n1293), .A4(n1007), .ZN(n1292) );
INV_X1 U1035 ( .A(n1294), .ZN(n1293) );
XOR2_X1 U1036 ( .A(n1295), .B(KEYINPUT42), .Z(n1291) );
NAND2_X1 U1037 ( .A1(n1294), .A2(n1296), .ZN(n1295) );
NAND3_X1 U1038 ( .A1(G234), .A2(n1007), .A3(G217), .ZN(n1296) );
INV_X1 U1039 ( .A(G953), .ZN(n1007) );
XNOR2_X1 U1040 ( .A(n1263), .B(n1297), .ZN(n1294) );
XOR2_X1 U1041 ( .A(G134), .B(n1298), .Z(n1297) );
NOR2_X1 U1042 ( .A1(KEYINPUT41), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1043 ( .A(n1300), .B(n1273), .Z(n1299) );
XOR2_X1 U1044 ( .A(G116), .B(KEYINPUT27), .Z(n1273) );
XOR2_X1 U1045 ( .A(n986), .B(G122), .Z(n1300) );
INV_X1 U1046 ( .A(G107), .ZN(n986) );
XOR2_X1 U1047 ( .A(G128), .B(G143), .Z(n1263) );
INV_X1 U1048 ( .A(G902), .ZN(n1218) );
endmodule


