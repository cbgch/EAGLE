//Key = 1110000101000100000010001111100110001100100100110111000010101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;

XNOR2_X1 U744 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
INV_X1 U748 ( .A(n1030), .ZN(n1029) );
NOR2_X1 U749 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
NOR2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
INV_X1 U751 ( .A(n1035), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
NOR2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
NOR2_X1 U754 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR3_X1 U755 ( .A1(n1042), .A2(KEYINPUT11), .A3(n1043), .ZN(n1040) );
NAND3_X1 U756 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1024) );
NAND3_X1 U757 ( .A1(n1047), .A2(n1048), .A3(n1035), .ZN(n1046) );
NAND3_X1 U758 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND2_X1 U759 ( .A1(KEYINPUT11), .A2(n1030), .ZN(n1051) );
NOR3_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1030) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1050) );
NAND3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U767 ( .A1(KEYINPUT50), .A2(n1068), .ZN(n1064) );
OR4_X1 U768 ( .A1(n1069), .A2(KEYINPUT50), .A3(n1053), .A4(n1055), .ZN(n1049) );
INV_X1 U769 ( .A(n1054), .ZN(n1055) );
NOR3_X1 U770 ( .A1(n1070), .A2(G953), .A3(n1071), .ZN(n1022) );
INV_X1 U771 ( .A(n1044), .ZN(n1071) );
NAND4_X1 U772 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1044) );
NOR4_X1 U773 ( .A1(n1076), .A2(n1066), .A3(n1077), .A4(n1078), .ZN(n1075) );
XOR2_X1 U774 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U775 ( .A1(n1081), .A2(KEYINPUT6), .ZN(n1080) );
XNOR2_X1 U776 ( .A(n1082), .B(n1083), .ZN(n1077) );
NAND2_X1 U777 ( .A1(KEYINPUT61), .A2(n1084), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1074) );
XNOR2_X1 U779 ( .A(KEYINPUT15), .B(n1087), .ZN(n1086) );
XNOR2_X1 U780 ( .A(KEYINPUT29), .B(n1088), .ZN(n1085) );
XNOR2_X1 U781 ( .A(n1089), .B(n1090), .ZN(n1072) );
NAND2_X1 U782 ( .A1(KEYINPUT58), .A2(G469), .ZN(n1089) );
XNOR2_X1 U783 ( .A(KEYINPUT53), .B(n1027), .ZN(n1070) );
INV_X1 U784 ( .A(G952), .ZN(n1027) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(G72) );
XOR2_X1 U786 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1097), .A2(G953), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1098), .B(n1099), .Z(n1095) );
XOR2_X1 U790 ( .A(n1100), .B(n1101), .Z(n1098) );
NAND2_X1 U791 ( .A1(n1102), .A2(n1045), .ZN(n1093) );
NAND3_X1 U792 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1045), .ZN(n1091) );
AND2_X1 U794 ( .A1(G227), .A2(G900), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U796 ( .A1(n1109), .A2(n1045), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U798 ( .A1(n1112), .A2(KEYINPUT60), .ZN(n1107) );
XOR2_X1 U799 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U801 ( .A(n1117), .B(n1118), .ZN(n1116) );
XOR2_X1 U802 ( .A(n1119), .B(KEYINPUT46), .Z(n1118) );
NOR2_X1 U803 ( .A1(G898), .A2(n1045), .ZN(n1115) );
NAND2_X1 U804 ( .A1(n1045), .A2(n1120), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U806 ( .A(n1123), .B(n1124), .Z(n1122) );
AND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND3_X1 U808 ( .A1(n1127), .A2(n1128), .A3(KEYINPUT2), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1121), .A2(n1129), .ZN(G63) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U811 ( .A(KEYINPUT56), .B(n1132), .Z(n1131) );
AND2_X1 U812 ( .A1(G478), .A2(n1127), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1133), .ZN(G60) );
XOR2_X1 U814 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U815 ( .A1(n1127), .A2(G475), .A3(KEYINPUT27), .ZN(n1134) );
XOR2_X1 U816 ( .A(G104), .B(n1136), .Z(G6) );
NOR2_X1 U817 ( .A1(KEYINPUT34), .A2(n1137), .ZN(n1136) );
NOR2_X1 U818 ( .A1(n1121), .A2(n1138), .ZN(G57) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U820 ( .A1(n1084), .A2(n1141), .ZN(n1139) );
INV_X1 U821 ( .A(G472), .ZN(n1084) );
NOR2_X1 U822 ( .A1(n1142), .A2(n1143), .ZN(G54) );
XOR2_X1 U823 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U824 ( .A(n1099), .B(n1146), .Z(n1145) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U826 ( .A1(KEYINPUT9), .A2(n1149), .ZN(n1147) );
XNOR2_X1 U827 ( .A(n1150), .B(n1151), .ZN(n1099) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1144) );
XNOR2_X1 U829 ( .A(G110), .B(n1154), .ZN(n1153) );
AND2_X1 U830 ( .A1(G469), .A2(n1127), .ZN(n1154) );
NAND2_X1 U831 ( .A1(KEYINPUT13), .A2(n1155), .ZN(n1152) );
NAND2_X1 U832 ( .A1(G227), .A2(n1045), .ZN(n1155) );
XNOR2_X1 U833 ( .A(n1121), .B(KEYINPUT43), .ZN(n1142) );
NOR2_X1 U834 ( .A1(n1121), .A2(n1156), .ZN(G51) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(n1158) );
AND3_X1 U837 ( .A1(n1127), .A2(n1161), .A3(G210), .ZN(n1160) );
INV_X1 U838 ( .A(n1141), .ZN(n1127) );
NAND2_X1 U839 ( .A1(G902), .A2(n1025), .ZN(n1141) );
NAND4_X1 U840 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1105), .ZN(n1025) );
AND4_X1 U841 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1105) );
NOR3_X1 U842 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1168) );
NOR4_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1052), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
INV_X1 U845 ( .A(KEYINPUT18), .ZN(n1176) );
NOR3_X1 U846 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1175) );
NOR2_X1 U847 ( .A1(KEYINPUT18), .A2(n1180), .ZN(n1172) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1058), .ZN(n1169) );
INV_X1 U849 ( .A(n1120), .ZN(n1164) );
NAND2_X1 U850 ( .A1(n1182), .A2(n1183), .ZN(n1120) );
AND4_X1 U851 ( .A1(n1184), .A2(n1021), .A3(n1185), .A4(n1186), .ZN(n1183) );
NAND3_X1 U852 ( .A1(n1061), .A2(n1187), .A3(n1041), .ZN(n1021) );
NOR4_X1 U853 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1182) );
INV_X1 U854 ( .A(n1137), .ZN(n1191) );
NAND3_X1 U855 ( .A1(n1041), .A2(n1187), .A3(n1192), .ZN(n1137) );
NOR3_X1 U856 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1190) );
XNOR2_X1 U857 ( .A(n1068), .B(KEYINPUT5), .ZN(n1195) );
NOR4_X1 U858 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1053), .ZN(n1189) );
INV_X1 U859 ( .A(n1062), .ZN(n1053) );
INV_X1 U860 ( .A(n1037), .ZN(n1197) );
XNOR2_X1 U861 ( .A(n1041), .B(KEYINPUT38), .ZN(n1196) );
XOR2_X1 U862 ( .A(n1104), .B(KEYINPUT45), .Z(n1163) );
NAND2_X1 U863 ( .A1(n1199), .A2(n1060), .ZN(n1104) );
XOR2_X1 U864 ( .A(n1200), .B(KEYINPUT37), .Z(n1199) );
XOR2_X1 U865 ( .A(n1103), .B(KEYINPUT42), .Z(n1162) );
XNOR2_X1 U866 ( .A(G128), .B(n1201), .ZN(n1157) );
NOR2_X1 U867 ( .A1(KEYINPUT30), .A2(n1202), .ZN(n1201) );
XOR2_X1 U868 ( .A(n1203), .B(n1117), .Z(n1202) );
XOR2_X1 U869 ( .A(G110), .B(G122), .Z(n1117) );
AND2_X1 U870 ( .A1(n1204), .A2(G953), .ZN(n1121) );
XNOR2_X1 U871 ( .A(G952), .B(KEYINPUT54), .ZN(n1204) );
XNOR2_X1 U872 ( .A(n1205), .B(n1170), .ZN(G48) );
AND3_X1 U873 ( .A1(n1192), .A2(n1068), .A3(n1206), .ZN(n1170) );
XNOR2_X1 U874 ( .A(G143), .B(n1167), .ZN(G45) );
NAND4_X1 U875 ( .A1(n1180), .A2(n1068), .A3(n1207), .A4(n1208), .ZN(n1167) );
NAND2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(G42) );
NAND2_X1 U877 ( .A1(KEYINPUT62), .A2(G140), .ZN(n1210) );
XOR2_X1 U878 ( .A(n1211), .B(n1212), .Z(n1209) );
NOR2_X1 U879 ( .A1(n1052), .A2(n1200), .ZN(n1212) );
NAND4_X1 U880 ( .A1(n1192), .A2(n1041), .A3(n1037), .A4(n1177), .ZN(n1200) );
NOR2_X1 U881 ( .A1(G140), .A2(KEYINPUT62), .ZN(n1211) );
XNOR2_X1 U882 ( .A(n1165), .B(n1213), .ZN(G39) );
NOR2_X1 U883 ( .A1(KEYINPUT3), .A2(n1214), .ZN(n1213) );
NAND3_X1 U884 ( .A1(n1060), .A2(n1062), .A3(n1206), .ZN(n1165) );
XNOR2_X1 U885 ( .A(n1215), .B(n1216), .ZN(G36) );
NOR3_X1 U886 ( .A1(n1181), .A2(n1174), .A3(n1052), .ZN(n1216) );
INV_X1 U887 ( .A(n1061), .ZN(n1174) );
XNOR2_X1 U888 ( .A(G131), .B(n1217), .ZN(G33) );
NOR2_X1 U889 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR3_X1 U890 ( .A1(n1220), .A2(n1181), .A3(n1058), .ZN(n1219) );
NAND2_X1 U891 ( .A1(n1060), .A2(n1192), .ZN(n1058) );
INV_X1 U892 ( .A(n1052), .ZN(n1060) );
INV_X1 U893 ( .A(KEYINPUT40), .ZN(n1220) );
NOR3_X1 U894 ( .A1(KEYINPUT40), .A2(n1221), .A3(n1052), .ZN(n1218) );
NAND2_X1 U895 ( .A1(n1067), .A2(n1222), .ZN(n1052) );
AND2_X1 U896 ( .A1(n1192), .A2(n1180), .ZN(n1221) );
INV_X1 U897 ( .A(n1181), .ZN(n1180) );
NAND3_X1 U898 ( .A1(n1041), .A2(n1177), .A3(n1036), .ZN(n1181) );
INV_X1 U899 ( .A(n1179), .ZN(n1036) );
XNOR2_X1 U900 ( .A(n1223), .B(n1224), .ZN(G30) );
NAND2_X1 U901 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
OR2_X1 U902 ( .A1(n1103), .A2(KEYINPUT48), .ZN(n1226) );
NAND3_X1 U903 ( .A1(n1061), .A2(n1068), .A3(n1206), .ZN(n1103) );
NAND4_X1 U904 ( .A1(n1061), .A2(n1069), .A3(n1206), .A4(KEYINPUT48), .ZN(n1225) );
AND4_X1 U905 ( .A1(n1041), .A2(n1227), .A3(n1228), .A4(n1177), .ZN(n1206) );
XOR2_X1 U906 ( .A(G101), .B(n1188), .Z(G3) );
AND3_X1 U907 ( .A1(n1229), .A2(n1041), .A3(n1062), .ZN(n1188) );
XNOR2_X1 U908 ( .A(G125), .B(n1166), .ZN(G27) );
NAND3_X1 U909 ( .A1(n1192), .A2(n1035), .A3(n1230), .ZN(n1166) );
AND3_X1 U910 ( .A1(n1037), .A2(n1177), .A3(n1068), .ZN(n1230) );
NAND2_X1 U911 ( .A1(n1054), .A2(n1231), .ZN(n1177) );
NAND4_X1 U912 ( .A1(n1097), .A2(G953), .A3(G902), .A4(n1232), .ZN(n1231) );
XNOR2_X1 U913 ( .A(G900), .B(KEYINPUT52), .ZN(n1097) );
XNOR2_X1 U914 ( .A(G122), .B(n1186), .ZN(G24) );
NAND4_X1 U915 ( .A1(n1035), .A2(n1187), .A3(n1207), .A4(n1208), .ZN(n1186) );
NOR2_X1 U916 ( .A1(n1198), .A2(n1039), .ZN(n1187) );
INV_X1 U917 ( .A(n1047), .ZN(n1039) );
NAND2_X1 U918 ( .A1(n1233), .A2(n1234), .ZN(n1047) );
OR3_X1 U919 ( .A1(n1228), .A2(n1227), .A3(KEYINPUT55), .ZN(n1234) );
NAND2_X1 U920 ( .A1(KEYINPUT55), .A2(n1037), .ZN(n1233) );
NAND2_X1 U921 ( .A1(n1235), .A2(n1236), .ZN(G21) );
OR2_X1 U922 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U923 ( .A(n1239), .B(KEYINPUT35), .Z(n1235) );
NAND2_X1 U924 ( .A1(n1238), .A2(n1237), .ZN(n1239) );
NOR2_X1 U925 ( .A1(n1193), .A2(n1198), .ZN(n1238) );
NAND4_X1 U926 ( .A1(n1062), .A2(n1035), .A3(n1227), .A4(n1228), .ZN(n1193) );
XNOR2_X1 U927 ( .A(G116), .B(n1184), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1229), .A2(n1061), .A3(n1035), .ZN(n1184) );
NOR2_X1 U929 ( .A1(n1208), .A2(n1087), .ZN(n1061) );
INV_X1 U930 ( .A(n1207), .ZN(n1087) );
XNOR2_X1 U931 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U932 ( .A1(n1035), .A2(n1229), .A3(n1192), .ZN(n1185) );
NOR2_X1 U933 ( .A1(n1207), .A2(n1088), .ZN(n1192) );
INV_X1 U934 ( .A(n1208), .ZN(n1088) );
NOR2_X1 U935 ( .A1(n1179), .A2(n1198), .ZN(n1229) );
INV_X1 U936 ( .A(n1240), .ZN(n1198) );
NAND2_X1 U937 ( .A1(n1073), .A2(n1228), .ZN(n1179) );
NOR2_X1 U938 ( .A1(n1043), .A2(n1076), .ZN(n1035) );
INV_X1 U939 ( .A(n1042), .ZN(n1076) );
XOR2_X1 U940 ( .A(n1241), .B(G110), .Z(G12) );
NAND2_X1 U941 ( .A1(KEYINPUT63), .A2(n1242), .ZN(n1241) );
NAND4_X1 U942 ( .A1(n1062), .A2(n1041), .A3(n1240), .A4(n1037), .ZN(n1242) );
NOR2_X1 U943 ( .A1(n1228), .A2(n1073), .ZN(n1037) );
INV_X1 U944 ( .A(n1227), .ZN(n1073) );
XNOR2_X1 U945 ( .A(n1243), .B(n1128), .ZN(n1227) );
AND2_X1 U946 ( .A1(G217), .A2(n1244), .ZN(n1128) );
NAND3_X1 U947 ( .A1(n1126), .A2(n1245), .A3(n1125), .ZN(n1243) );
NAND2_X1 U948 ( .A1(n1246), .A2(n1247), .ZN(n1125) );
XNOR2_X1 U949 ( .A(n1248), .B(n1101), .ZN(n1246) );
NAND2_X1 U950 ( .A1(n1249), .A2(n1250), .ZN(n1126) );
XNOR2_X1 U951 ( .A(n1251), .B(n1101), .ZN(n1250) );
XNOR2_X1 U952 ( .A(G125), .B(n1149), .ZN(n1101) );
INV_X1 U953 ( .A(n1248), .ZN(n1251) );
XNOR2_X1 U954 ( .A(n1252), .B(KEYINPUT12), .ZN(n1248) );
NAND2_X1 U955 ( .A1(KEYINPUT24), .A2(G146), .ZN(n1252) );
XOR2_X1 U956 ( .A(n1247), .B(KEYINPUT32), .Z(n1249) );
XOR2_X1 U957 ( .A(n1253), .B(n1254), .Z(n1247) );
XNOR2_X1 U958 ( .A(n1255), .B(n1237), .ZN(n1253) );
INV_X1 U959 ( .A(G119), .ZN(n1237) );
NAND2_X1 U960 ( .A1(KEYINPUT47), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U961 ( .A(n1214), .B(n1257), .ZN(n1256) );
AND3_X1 U962 ( .A1(G221), .A2(n1045), .A3(G234), .ZN(n1257) );
XNOR2_X1 U963 ( .A(n1083), .B(G472), .ZN(n1228) );
NAND2_X1 U964 ( .A1(n1258), .A2(n1245), .ZN(n1083) );
XNOR2_X1 U965 ( .A(n1140), .B(n1259), .ZN(n1258) );
XOR2_X1 U966 ( .A(KEYINPUT41), .B(KEYINPUT22), .Z(n1259) );
XNOR2_X1 U967 ( .A(n1260), .B(n1261), .ZN(n1140) );
XOR2_X1 U968 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U969 ( .A(n1264), .B(G101), .Z(n1263) );
XNOR2_X1 U970 ( .A(G113), .B(G119), .ZN(n1262) );
XNOR2_X1 U971 ( .A(n1265), .B(n1150), .ZN(n1260) );
XOR2_X1 U972 ( .A(n1266), .B(n1267), .Z(n1265) );
AND3_X1 U973 ( .A1(G210), .A2(n1045), .A3(n1268), .ZN(n1267) );
NOR2_X1 U974 ( .A1(n1069), .A2(n1194), .ZN(n1240) );
AND2_X1 U975 ( .A1(n1054), .A2(n1269), .ZN(n1194) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1232), .A4(n1111), .ZN(n1269) );
INV_X1 U977 ( .A(G898), .ZN(n1111) );
NAND3_X1 U978 ( .A1(n1232), .A2(n1045), .A3(G952), .ZN(n1054) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1232) );
INV_X1 U980 ( .A(n1068), .ZN(n1069) );
NOR2_X1 U981 ( .A1(n1067), .A2(n1066), .ZN(n1068) );
INV_X1 U982 ( .A(n1222), .ZN(n1066) );
NAND2_X1 U983 ( .A1(G214), .A2(n1161), .ZN(n1222) );
XOR2_X1 U984 ( .A(n1079), .B(n1081), .Z(n1067) );
AND2_X1 U985 ( .A1(G210), .A2(n1270), .ZN(n1081) );
XNOR2_X1 U986 ( .A(KEYINPUT31), .B(n1161), .ZN(n1270) );
NAND2_X1 U987 ( .A1(n1271), .A2(n1268), .ZN(n1161) );
NAND2_X1 U988 ( .A1(n1272), .A2(n1245), .ZN(n1079) );
XOR2_X1 U989 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U990 ( .A(n1254), .B(n1159), .ZN(n1274) );
XOR2_X1 U991 ( .A(n1275), .B(n1276), .Z(n1159) );
NOR2_X1 U992 ( .A1(G953), .A2(n1110), .ZN(n1276) );
INV_X1 U993 ( .A(G224), .ZN(n1110) );
XOR2_X1 U994 ( .A(n1264), .B(G125), .Z(n1275) );
NAND3_X1 U995 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1264) );
NAND2_X1 U996 ( .A1(G146), .A2(n1280), .ZN(n1279) );
NAND2_X1 U997 ( .A1(KEYINPUT19), .A2(n1281), .ZN(n1278) );
NAND2_X1 U998 ( .A1(n1282), .A2(n1205), .ZN(n1281) );
XNOR2_X1 U999 ( .A(KEYINPUT57), .B(n1280), .ZN(n1282) );
NAND2_X1 U1000 ( .A1(n1283), .A2(n1284), .ZN(n1277) );
INV_X1 U1001 ( .A(KEYINPUT19), .ZN(n1284) );
NAND2_X1 U1002 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U1003 ( .A1(KEYINPUT57), .A2(n1280), .ZN(n1286) );
OR3_X1 U1004 ( .A1(G146), .A2(KEYINPUT57), .A3(n1280), .ZN(n1285) );
XNOR2_X1 U1005 ( .A(G110), .B(n1224), .ZN(n1254) );
XOR2_X1 U1006 ( .A(G122), .B(n1203), .Z(n1273) );
NOR2_X1 U1007 ( .A1(KEYINPUT4), .A2(n1119), .ZN(n1203) );
XOR2_X1 U1008 ( .A(n1287), .B(n1288), .Z(n1119) );
XNOR2_X1 U1009 ( .A(n1289), .B(n1290), .ZN(n1288) );
NOR2_X1 U1010 ( .A1(KEYINPUT39), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U1011 ( .A(G116), .B(G119), .ZN(n1291) );
INV_X1 U1012 ( .A(G113), .ZN(n1289) );
NAND2_X1 U1013 ( .A1(n1292), .A2(n1293), .ZN(n1287) );
NAND2_X1 U1014 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
INV_X1 U1015 ( .A(KEYINPUT10), .ZN(n1295) );
NAND2_X1 U1016 ( .A1(KEYINPUT10), .A2(n1296), .ZN(n1292) );
XNOR2_X1 U1017 ( .A(G101), .B(n1297), .ZN(n1296) );
NOR2_X1 U1018 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U1019 ( .A(n1178), .ZN(n1041) );
NAND2_X1 U1020 ( .A1(n1043), .A2(n1042), .ZN(n1178) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1244), .ZN(n1042) );
NAND2_X1 U1022 ( .A1(n1271), .A2(G234), .ZN(n1244) );
XNOR2_X1 U1023 ( .A(KEYINPUT59), .B(G902), .ZN(n1271) );
XOR2_X1 U1024 ( .A(n1090), .B(n1300), .Z(n1043) );
NOR2_X1 U1025 ( .A1(G469), .A2(KEYINPUT23), .ZN(n1300) );
NAND2_X1 U1026 ( .A1(n1301), .A2(n1245), .ZN(n1090) );
XOR2_X1 U1027 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1028 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U1029 ( .A1(G110), .A2(KEYINPUT33), .ZN(n1305) );
NAND3_X1 U1030 ( .A1(n1306), .A2(n1307), .A3(KEYINPUT49), .ZN(n1304) );
NAND2_X1 U1031 ( .A1(KEYINPUT28), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1032 ( .A(n1309), .B(n1310), .ZN(n1308) );
NOR2_X1 U1033 ( .A1(KEYINPUT17), .A2(n1311), .ZN(n1310) );
NAND3_X1 U1034 ( .A1(n1309), .A2(n1311), .A3(n1312), .ZN(n1306) );
INV_X1 U1035 ( .A(KEYINPUT28), .ZN(n1312) );
XNOR2_X1 U1036 ( .A(n1148), .B(n1224), .ZN(n1311) );
INV_X1 U1037 ( .A(G128), .ZN(n1224) );
XNOR2_X1 U1038 ( .A(n1294), .B(n1100), .ZN(n1148) );
NAND3_X1 U1039 ( .A1(n1313), .A2(n1314), .A3(KEYINPUT0), .ZN(n1100) );
NAND2_X1 U1040 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U1041 ( .A(KEYINPUT16), .B(n1280), .ZN(n1316) );
XNOR2_X1 U1042 ( .A(KEYINPUT36), .B(G146), .ZN(n1315) );
NAND2_X1 U1043 ( .A1(n1317), .A2(n1318), .ZN(n1313) );
XNOR2_X1 U1044 ( .A(KEYINPUT26), .B(n1280), .ZN(n1318) );
INV_X1 U1045 ( .A(G143), .ZN(n1280) );
XNOR2_X1 U1046 ( .A(KEYINPUT36), .B(n1205), .ZN(n1317) );
XOR2_X1 U1047 ( .A(n1319), .B(n1299), .Z(n1294) );
XOR2_X1 U1048 ( .A(G104), .B(KEYINPUT7), .Z(n1299) );
XNOR2_X1 U1049 ( .A(G101), .B(n1298), .ZN(n1319) );
XNOR2_X1 U1050 ( .A(G134), .B(n1150), .ZN(n1309) );
XNOR2_X1 U1051 ( .A(n1214), .B(n1320), .ZN(n1150) );
INV_X1 U1052 ( .A(G137), .ZN(n1214) );
XNOR2_X1 U1053 ( .A(G227), .B(n1149), .ZN(n1302) );
INV_X1 U1054 ( .A(G140), .ZN(n1149) );
NOR2_X1 U1055 ( .A1(n1207), .A2(n1208), .ZN(n1062) );
XNOR2_X1 U1056 ( .A(n1321), .B(G475), .ZN(n1208) );
NAND2_X1 U1057 ( .A1(n1135), .A2(n1245), .ZN(n1321) );
XOR2_X1 U1058 ( .A(n1322), .B(n1323), .Z(n1135) );
XOR2_X1 U1059 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1060 ( .A(G104), .B(n1326), .ZN(n1325) );
NAND2_X1 U1061 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1062 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1063 ( .A1(KEYINPUT25), .A2(n1331), .ZN(n1330) );
NAND2_X1 U1064 ( .A1(G131), .A2(n1332), .ZN(n1331) );
NAND2_X1 U1065 ( .A1(n1333), .A2(n1320), .ZN(n1327) );
INV_X1 U1066 ( .A(G131), .ZN(n1320) );
NAND2_X1 U1067 ( .A1(n1332), .A2(n1334), .ZN(n1333) );
NAND2_X1 U1068 ( .A1(n1335), .A2(KEYINPUT25), .ZN(n1334) );
INV_X1 U1069 ( .A(n1329), .ZN(n1335) );
XNOR2_X1 U1070 ( .A(n1336), .B(n1337), .ZN(n1329) );
AND3_X1 U1071 ( .A1(G214), .A2(n1045), .A3(n1268), .ZN(n1337) );
INV_X1 U1072 ( .A(G237), .ZN(n1268) );
NAND2_X1 U1073 ( .A1(KEYINPUT1), .A2(G143), .ZN(n1336) );
INV_X1 U1074 ( .A(KEYINPUT21), .ZN(n1332) );
NOR2_X1 U1075 ( .A1(G140), .A2(KEYINPUT14), .ZN(n1324) );
XOR2_X1 U1076 ( .A(n1338), .B(n1339), .Z(n1322) );
XNOR2_X1 U1077 ( .A(n1205), .B(G125), .ZN(n1339) );
INV_X1 U1078 ( .A(G146), .ZN(n1205) );
XNOR2_X1 U1079 ( .A(G113), .B(G122), .ZN(n1338) );
XNOR2_X1 U1080 ( .A(n1340), .B(G478), .ZN(n1207) );
NAND2_X1 U1081 ( .A1(n1245), .A2(n1130), .ZN(n1340) );
NAND2_X1 U1082 ( .A1(n1341), .A2(n1342), .ZN(n1130) );
NAND4_X1 U1083 ( .A1(G217), .A2(G234), .A3(n1343), .A4(n1045), .ZN(n1342) );
NAND2_X1 U1084 ( .A1(n1344), .A2(n1345), .ZN(n1341) );
NAND3_X1 U1085 ( .A1(G234), .A2(n1045), .A3(G217), .ZN(n1345) );
INV_X1 U1086 ( .A(G953), .ZN(n1045) );
XOR2_X1 U1087 ( .A(KEYINPUT20), .B(n1343), .Z(n1344) );
XNOR2_X1 U1088 ( .A(n1346), .B(n1347), .ZN(n1343) );
XNOR2_X1 U1089 ( .A(G143), .B(n1348), .ZN(n1347) );
XNOR2_X1 U1090 ( .A(KEYINPUT8), .B(KEYINPUT51), .ZN(n1348) );
XOR2_X1 U1091 ( .A(n1349), .B(n1298), .Z(n1346) );
XOR2_X1 U1092 ( .A(G107), .B(KEYINPUT44), .Z(n1298) );
XOR2_X1 U1093 ( .A(n1266), .B(G122), .Z(n1349) );
XNOR2_X1 U1094 ( .A(G116), .B(n1151), .ZN(n1266) );
XNOR2_X1 U1095 ( .A(n1215), .B(G128), .ZN(n1151) );
INV_X1 U1096 ( .A(G134), .ZN(n1215) );
INV_X1 U1097 ( .A(G902), .ZN(n1245) );
endmodule


