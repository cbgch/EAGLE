//Key = 0100000010010101111100000010100010000001000101100001100011000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;

XOR2_X1 U702 ( .A(G107), .B(n962), .Z(G9) );
NOR2_X1 U703 ( .A1(n963), .A2(n964), .ZN(G75) );
NOR4_X1 U704 ( .A1(G953), .A2(n965), .A3(n966), .A4(n967), .ZN(n964) );
XOR2_X1 U705 ( .A(n968), .B(KEYINPUT20), .Z(n966) );
NAND3_X1 U706 ( .A1(n969), .A2(n970), .A3(n971), .ZN(n968) );
NAND2_X1 U707 ( .A1(n972), .A2(n973), .ZN(n970) );
NAND2_X1 U708 ( .A1(n974), .A2(n975), .ZN(n973) );
NAND3_X1 U709 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n975) );
NAND2_X1 U710 ( .A1(n979), .A2(n980), .ZN(n977) );
NAND3_X1 U711 ( .A1(n981), .A2(n982), .A3(KEYINPUT3), .ZN(n979) );
NAND3_X1 U712 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n976) );
NAND2_X1 U713 ( .A1(n986), .A2(n987), .ZN(n984) );
OR2_X1 U714 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND2_X1 U715 ( .A1(n981), .A2(n990), .ZN(n983) );
NAND2_X1 U716 ( .A1(n991), .A2(n992), .ZN(n990) );
OR2_X1 U717 ( .A1(n993), .A2(KEYINPUT3), .ZN(n992) );
NAND2_X1 U718 ( .A1(n994), .A2(n995), .ZN(n991) );
NAND3_X1 U719 ( .A1(n986), .A2(n996), .A3(n981), .ZN(n974) );
NAND3_X1 U720 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NAND2_X1 U721 ( .A1(n1000), .A2(n985), .ZN(n999) );
NAND3_X1 U722 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n998) );
XOR2_X1 U723 ( .A(KEYINPUT12), .B(n985), .Z(n1001) );
NAND2_X1 U724 ( .A1(n978), .A2(n1004), .ZN(n997) );
NAND2_X1 U725 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U726 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
INV_X1 U727 ( .A(n1009), .ZN(n972) );
NOR3_X1 U728 ( .A1(n1010), .A2(G953), .A3(n965), .ZN(n963) );
AND4_X1 U729 ( .A1(n986), .A2(n985), .A3(n1011), .A4(n1012), .ZN(n965) );
NOR4_X1 U730 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
XOR2_X1 U731 ( .A(n1017), .B(KEYINPUT25), .Z(n1016) );
NAND2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
XNOR2_X1 U733 ( .A(n1020), .B(KEYINPUT13), .ZN(n1015) );
NOR2_X1 U734 ( .A1(n1021), .A2(n1022), .ZN(n1014) );
NOR2_X1 U735 ( .A1(G902), .A2(n1023), .ZN(n1021) );
XOR2_X1 U736 ( .A(n1024), .B(KEYINPUT11), .Z(n1011) );
NAND3_X1 U737 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
OR3_X1 U738 ( .A1(n1028), .A2(n1029), .A3(KEYINPUT23), .ZN(n1026) );
NAND2_X1 U739 ( .A1(KEYINPUT23), .A2(n1029), .ZN(n1025) );
XOR2_X1 U740 ( .A(KEYINPUT59), .B(G952), .Z(n1010) );
XOR2_X1 U741 ( .A(n1030), .B(n1031), .Z(G72) );
XOR2_X1 U742 ( .A(n1032), .B(n1033), .Z(n1031) );
NOR3_X1 U743 ( .A1(n969), .A2(KEYINPUT30), .A3(G953), .ZN(n1033) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
XOR2_X1 U745 ( .A(n1036), .B(n1037), .Z(n1035) );
XNOR2_X1 U746 ( .A(n1038), .B(n1039), .ZN(n1037) );
NOR2_X1 U747 ( .A1(KEYINPUT0), .A2(n1040), .ZN(n1039) );
XOR2_X1 U748 ( .A(n1041), .B(n1042), .Z(n1036) );
XOR2_X1 U749 ( .A(KEYINPUT6), .B(G125), .Z(n1042) );
NAND2_X1 U750 ( .A1(KEYINPUT15), .A2(n1043), .ZN(n1041) );
NOR2_X1 U751 ( .A1(G900), .A2(n1044), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1044), .ZN(n1030) );
AND2_X1 U753 ( .A1(G227), .A2(G900), .ZN(n1045) );
XOR2_X1 U754 ( .A(n1046), .B(n1047), .Z(G69) );
NOR2_X1 U755 ( .A1(n1048), .A2(n1044), .ZN(n1047) );
AND2_X1 U756 ( .A1(G224), .A2(G898), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
NAND3_X1 U758 ( .A1(n1051), .A2(n1052), .A3(n971), .ZN(n1050) );
XOR2_X1 U759 ( .A(n1053), .B(n1054), .Z(n1052) );
NAND2_X1 U760 ( .A1(G953), .A2(n1055), .ZN(n1051) );
XOR2_X1 U761 ( .A(n1056), .B(KEYINPUT9), .Z(n1049) );
NAND3_X1 U762 ( .A1(n1057), .A2(n1044), .A3(n1058), .ZN(n1056) );
XOR2_X1 U763 ( .A(n1054), .B(n1059), .Z(n1058) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(G66) );
XOR2_X1 U765 ( .A(n1062), .B(n1063), .Z(n1061) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U767 ( .A1(n1060), .A2(n1066), .ZN(G63) );
XOR2_X1 U768 ( .A(n1067), .B(n1023), .Z(n1066) );
NOR3_X1 U769 ( .A1(n1022), .A2(n1068), .A3(n1069), .ZN(n1067) );
XOR2_X1 U770 ( .A(n1070), .B(KEYINPUT56), .Z(n1069) );
INV_X1 U771 ( .A(n1071), .ZN(n1068) );
INV_X1 U772 ( .A(G478), .ZN(n1022) );
NOR2_X1 U773 ( .A1(n1060), .A2(n1072), .ZN(G60) );
XOR2_X1 U774 ( .A(n1073), .B(n1074), .Z(n1072) );
NAND2_X1 U775 ( .A1(n1064), .A2(G475), .ZN(n1073) );
XOR2_X1 U776 ( .A(n1075), .B(n1076), .Z(G6) );
NOR2_X1 U777 ( .A1(n1060), .A2(n1077), .ZN(G57) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U779 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
AND2_X1 U781 ( .A1(KEYINPUT40), .A2(n1084), .ZN(n1083) );
NOR2_X1 U782 ( .A1(KEYINPUT44), .A2(n1084), .ZN(n1082) );
XOR2_X1 U783 ( .A(n1085), .B(n1086), .Z(n1078) );
XOR2_X1 U784 ( .A(n1087), .B(G101), .Z(n1086) );
NAND2_X1 U785 ( .A1(n1064), .A2(G472), .ZN(n1087) );
NAND3_X1 U786 ( .A1(n1088), .A2(G210), .A3(KEYINPUT52), .ZN(n1085) );
NOR2_X1 U787 ( .A1(n1060), .A2(n1089), .ZN(G54) );
XOR2_X1 U788 ( .A(n1090), .B(n1091), .Z(n1089) );
AND2_X1 U789 ( .A1(G469), .A2(n1064), .ZN(n1091) );
NAND2_X1 U790 ( .A1(KEYINPUT51), .A2(n1092), .ZN(n1090) );
XOR2_X1 U791 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U792 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U793 ( .A1(KEYINPUT34), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U794 ( .A(n1098), .B(n1099), .ZN(n1093) );
XOR2_X1 U795 ( .A(KEYINPUT16), .B(G140), .Z(n1099) );
NOR2_X1 U796 ( .A1(n1060), .A2(n1100), .ZN(G51) );
XOR2_X1 U797 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U798 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U799 ( .A1(n1064), .A2(n1105), .ZN(n1103) );
AND2_X1 U800 ( .A1(n1070), .A2(n1071), .ZN(n1064) );
NAND2_X1 U801 ( .A1(n971), .A2(n1106), .ZN(n1071) );
XOR2_X1 U802 ( .A(KEYINPUT47), .B(n969), .Z(n1106) );
AND4_X1 U803 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n969) );
NOR4_X1 U804 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NOR2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1109) );
NOR3_X1 U806 ( .A1(n1117), .A2(n1118), .A3(n1005), .ZN(n1116) );
XNOR2_X1 U807 ( .A(n986), .B(KEYINPUT21), .ZN(n1118) );
INV_X1 U808 ( .A(n1057), .ZN(n971) );
NAND4_X1 U809 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1057) );
AND4_X1 U810 ( .A1(n1123), .A2(n1124), .A3(n1076), .A4(n1125), .ZN(n1122) );
NAND3_X1 U811 ( .A1(n981), .A2(n1126), .A3(n1000), .ZN(n1125) );
NAND3_X1 U812 ( .A1(n1126), .A2(n978), .A3(n988), .ZN(n1076) );
NOR2_X1 U813 ( .A1(n1127), .A2(n962), .ZN(n1121) );
AND3_X1 U814 ( .A1(n989), .A2(n978), .A3(n1126), .ZN(n962) );
XOR2_X1 U815 ( .A(n1128), .B(KEYINPUT18), .Z(n1070) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(n1101) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U818 ( .A1(KEYINPUT41), .A2(n1133), .ZN(n1132) );
XOR2_X1 U819 ( .A(n1134), .B(KEYINPUT38), .Z(n1133) );
AND2_X1 U820 ( .A1(n1135), .A2(n967), .ZN(n1060) );
INV_X1 U821 ( .A(G952), .ZN(n967) );
XOR2_X1 U822 ( .A(KEYINPUT50), .B(G953), .Z(n1135) );
XOR2_X1 U823 ( .A(n1136), .B(n1115), .Z(G48) );
AND3_X1 U824 ( .A1(n988), .A2(n1137), .A3(n1138), .ZN(n1115) );
XOR2_X1 U825 ( .A(n1139), .B(KEYINPUT32), .Z(n1136) );
XNOR2_X1 U826 ( .A(G143), .B(n1107), .ZN(G45) );
NAND4_X1 U827 ( .A1(n982), .A2(n1137), .A3(n1000), .A4(n1140), .ZN(n1107) );
AND3_X1 U828 ( .A1(n1020), .A2(n1141), .A3(n1142), .ZN(n1140) );
XOR2_X1 U829 ( .A(n1143), .B(n1114), .Z(G42) );
NOR3_X1 U830 ( .A1(n980), .A2(n993), .A3(n1117), .ZN(n1114) );
XOR2_X1 U831 ( .A(n1043), .B(KEYINPUT19), .Z(n1143) );
NAND2_X1 U832 ( .A1(n1144), .A2(n1145), .ZN(G39) );
NAND2_X1 U833 ( .A1(G137), .A2(n1108), .ZN(n1145) );
XOR2_X1 U834 ( .A(KEYINPUT1), .B(n1146), .Z(n1144) );
NOR2_X1 U835 ( .A1(G137), .A2(n1108), .ZN(n1146) );
NAND3_X1 U836 ( .A1(n981), .A2(n985), .A3(n1138), .ZN(n1108) );
XOR2_X1 U837 ( .A(G134), .B(n1113), .Z(G36) );
AND2_X1 U838 ( .A1(n1147), .A2(n989), .ZN(n1113) );
XOR2_X1 U839 ( .A(G131), .B(n1112), .Z(G33) );
AND2_X1 U840 ( .A1(n1147), .A2(n988), .ZN(n1112) );
AND4_X1 U841 ( .A1(n1000), .A2(n985), .A3(n982), .A4(n1142), .ZN(n1147) );
INV_X1 U842 ( .A(n980), .ZN(n985) );
NAND2_X1 U843 ( .A1(n1008), .A2(n1148), .ZN(n980) );
XOR2_X1 U844 ( .A(G128), .B(n1111), .Z(G30) );
AND3_X1 U845 ( .A1(n989), .A2(n1137), .A3(n1138), .ZN(n1111) );
AND4_X1 U846 ( .A1(n982), .A2(n1149), .A3(n1142), .A4(n1002), .ZN(n1138) );
XOR2_X1 U847 ( .A(n1150), .B(n1151), .Z(G3) );
NAND4_X1 U848 ( .A1(n1152), .A2(n1153), .A3(n982), .A4(n1154), .ZN(n1151) );
AND2_X1 U849 ( .A1(n1000), .A2(n981), .ZN(n1154) );
XNOR2_X1 U850 ( .A(KEYINPUT48), .B(n1155), .ZN(n1152) );
XOR2_X1 U851 ( .A(G125), .B(n1156), .Z(G27) );
NOR2_X1 U852 ( .A1(n1157), .A2(n1117), .ZN(n1156) );
NAND4_X1 U853 ( .A1(n988), .A2(n1003), .A3(n1142), .A4(n1002), .ZN(n1117) );
NAND2_X1 U854 ( .A1(n1009), .A2(n1158), .ZN(n1142) );
NAND4_X1 U855 ( .A1(n1159), .A2(G953), .A3(G902), .A4(n1160), .ZN(n1158) );
XNOR2_X1 U856 ( .A(G900), .B(KEYINPUT5), .ZN(n1159) );
XNOR2_X1 U857 ( .A(G122), .B(n1124), .ZN(G24) );
NAND4_X1 U858 ( .A1(n1161), .A2(n978), .A3(n1020), .A4(n1141), .ZN(n1124) );
NOR2_X1 U859 ( .A1(n1162), .A2(n1002), .ZN(n978) );
XOR2_X1 U860 ( .A(n1163), .B(n1123), .Z(G21) );
NAND4_X1 U861 ( .A1(n1161), .A2(n981), .A3(n1149), .A4(n1002), .ZN(n1123) );
XOR2_X1 U862 ( .A(n1119), .B(n1164), .Z(G18) );
XNOR2_X1 U863 ( .A(G116), .B(KEYINPUT42), .ZN(n1164) );
NAND3_X1 U864 ( .A1(n1000), .A2(n989), .A3(n1161), .ZN(n1119) );
NOR2_X1 U865 ( .A1(n1157), .A2(n1165), .ZN(n1161) );
NAND2_X1 U866 ( .A1(n986), .A2(n1137), .ZN(n1157) );
NOR2_X1 U867 ( .A1(n1020), .A2(n1166), .ZN(n989) );
XOR2_X1 U868 ( .A(n1167), .B(G113), .Z(G15) );
NAND2_X1 U869 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U870 ( .A1(n1127), .A2(n1170), .ZN(n1169) );
INV_X1 U871 ( .A(KEYINPUT10), .ZN(n1170) );
NOR2_X1 U872 ( .A1(n1171), .A2(n1155), .ZN(n1127) );
NAND3_X1 U873 ( .A1(n1172), .A2(n1155), .A3(KEYINPUT10), .ZN(n1168) );
INV_X1 U874 ( .A(n1171), .ZN(n1172) );
NAND4_X1 U875 ( .A1(n1000), .A2(n988), .A3(n986), .A4(n1153), .ZN(n1171) );
NOR2_X1 U876 ( .A1(n1173), .A2(n994), .ZN(n986) );
INV_X1 U877 ( .A(n995), .ZN(n1173) );
AND2_X1 U878 ( .A1(n1166), .A2(n1020), .ZN(n988) );
INV_X1 U879 ( .A(n1141), .ZN(n1166) );
NOR2_X1 U880 ( .A1(n1002), .A2(n1174), .ZN(n1000) );
INV_X1 U881 ( .A(n1149), .ZN(n1174) );
XOR2_X1 U882 ( .A(n1003), .B(KEYINPUT62), .Z(n1149) );
XNOR2_X1 U883 ( .A(G110), .B(n1175), .ZN(G12) );
NAND2_X1 U884 ( .A1(KEYINPUT8), .A2(n1176), .ZN(n1175) );
INV_X1 U885 ( .A(n1120), .ZN(n1176) );
NAND4_X1 U886 ( .A1(n981), .A2(n1126), .A3(n1003), .A4(n1002), .ZN(n1120) );
NAND2_X1 U887 ( .A1(n1027), .A2(n1177), .ZN(n1002) );
NAND2_X1 U888 ( .A1(n1065), .A2(n1178), .ZN(n1177) );
INV_X1 U889 ( .A(n1028), .ZN(n1065) );
NAND2_X1 U890 ( .A1(n1029), .A2(n1028), .ZN(n1027) );
NAND2_X1 U891 ( .A1(G217), .A2(n1179), .ZN(n1028) );
INV_X1 U892 ( .A(n1178), .ZN(n1029) );
NAND2_X1 U893 ( .A1(n1063), .A2(n1128), .ZN(n1178) );
XOR2_X1 U894 ( .A(n1180), .B(n1181), .Z(n1063) );
XOR2_X1 U895 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U896 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U897 ( .A1(KEYINPUT27), .A2(n1186), .ZN(n1185) );
XOR2_X1 U898 ( .A(n1139), .B(n1187), .Z(n1186) );
NAND2_X1 U899 ( .A1(n1188), .A2(G221), .ZN(n1184) );
NAND3_X1 U900 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1182) );
NAND2_X1 U901 ( .A1(KEYINPUT54), .A2(G128), .ZN(n1191) );
NAND3_X1 U902 ( .A1(n1192), .A2(n1193), .A3(G119), .ZN(n1190) );
NAND2_X1 U903 ( .A1(n1194), .A2(n1163), .ZN(n1189) );
NAND2_X1 U904 ( .A1(n1195), .A2(n1193), .ZN(n1194) );
INV_X1 U905 ( .A(KEYINPUT54), .ZN(n1193) );
XOR2_X1 U906 ( .A(n1192), .B(KEYINPUT37), .Z(n1195) );
INV_X1 U907 ( .A(G128), .ZN(n1192) );
XOR2_X1 U908 ( .A(n1097), .B(n1196), .Z(n1180) );
NOR2_X1 U909 ( .A1(G137), .A2(KEYINPUT55), .ZN(n1196) );
INV_X1 U910 ( .A(n1162), .ZN(n1003) );
NAND2_X1 U911 ( .A1(n1197), .A2(n1019), .ZN(n1162) );
NAND3_X1 U912 ( .A1(n1198), .A2(n1128), .A3(n1199), .ZN(n1019) );
INV_X1 U913 ( .A(G472), .ZN(n1198) );
XOR2_X1 U914 ( .A(n1018), .B(KEYINPUT31), .Z(n1197) );
NAND2_X1 U915 ( .A1(G472), .A2(n1200), .ZN(n1018) );
NAND2_X1 U916 ( .A1(n1199), .A2(n1128), .ZN(n1200) );
XOR2_X1 U917 ( .A(n1201), .B(n1202), .Z(n1199) );
XOR2_X1 U918 ( .A(G101), .B(n1203), .Z(n1202) );
NOR2_X1 U919 ( .A1(KEYINPUT60), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U920 ( .A(n1084), .B(n1080), .ZN(n1204) );
XNOR2_X1 U921 ( .A(n1205), .B(n1206), .ZN(n1080) );
XOR2_X1 U922 ( .A(G113), .B(n1207), .Z(n1206) );
NOR2_X1 U923 ( .A1(KEYINPUT35), .A2(n1163), .ZN(n1207) );
XNOR2_X1 U924 ( .A(G116), .B(KEYINPUT58), .ZN(n1205) );
NAND3_X1 U925 ( .A1(n1088), .A2(G210), .A3(KEYINPUT43), .ZN(n1201) );
NOR3_X1 U926 ( .A1(n1155), .A2(n1165), .A3(n993), .ZN(n1126) );
INV_X1 U927 ( .A(n982), .ZN(n993) );
NOR2_X1 U928 ( .A1(n995), .A2(n994), .ZN(n982) );
AND2_X1 U929 ( .A1(G221), .A2(n1179), .ZN(n994) );
NAND2_X1 U930 ( .A1(G234), .A2(n1128), .ZN(n1179) );
XOR2_X1 U931 ( .A(n1208), .B(G469), .Z(n995) );
NAND2_X1 U932 ( .A1(n1209), .A2(n1128), .ZN(n1208) );
XOR2_X1 U933 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U934 ( .A(n1095), .B(n1097), .ZN(n1211) );
XOR2_X1 U935 ( .A(n1212), .B(n1213), .Z(n1095) );
XOR2_X1 U936 ( .A(n1084), .B(G101), .Z(n1212) );
XNOR2_X1 U937 ( .A(n1040), .B(n1038), .ZN(n1084) );
XNOR2_X1 U938 ( .A(n1104), .B(G131), .ZN(n1038) );
XOR2_X1 U939 ( .A(G134), .B(G137), .Z(n1040) );
XOR2_X1 U940 ( .A(n1214), .B(n1215), .Z(n1210) );
NOR2_X1 U941 ( .A1(KEYINPUT33), .A2(G140), .ZN(n1215) );
NAND2_X1 U942 ( .A1(KEYINPUT45), .A2(n1098), .ZN(n1214) );
AND2_X1 U943 ( .A1(G227), .A2(n1044), .ZN(n1098) );
INV_X1 U944 ( .A(n1153), .ZN(n1165) );
NAND2_X1 U945 ( .A1(n1009), .A2(n1216), .ZN(n1153) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1160), .A4(n1055), .ZN(n1216) );
INV_X1 U947 ( .A(G898), .ZN(n1055) );
NAND3_X1 U948 ( .A1(n1160), .A2(n1044), .A3(G952), .ZN(n1009) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1160) );
XOR2_X1 U950 ( .A(n1005), .B(KEYINPUT49), .Z(n1155) );
INV_X1 U951 ( .A(n1137), .ZN(n1005) );
NOR2_X1 U952 ( .A1(n1008), .A2(n1007), .ZN(n1137) );
INV_X1 U953 ( .A(n1148), .ZN(n1007) );
NAND2_X1 U954 ( .A1(n1217), .A2(n1218), .ZN(n1148) );
XOR2_X1 U955 ( .A(KEYINPUT7), .B(G214), .Z(n1217) );
XOR2_X1 U956 ( .A(n1219), .B(n1105), .Z(n1008) );
AND2_X1 U957 ( .A1(G210), .A2(n1218), .ZN(n1105) );
NAND2_X1 U958 ( .A1(n1220), .A2(n1128), .ZN(n1218) );
NAND2_X1 U959 ( .A1(n1221), .A2(n1128), .ZN(n1219) );
XOR2_X1 U960 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U961 ( .A(n1224), .B(n1104), .Z(n1223) );
XOR2_X1 U962 ( .A(G146), .B(n1225), .Z(n1104) );
NAND2_X1 U963 ( .A1(KEYINPUT26), .A2(n1131), .ZN(n1224) );
XOR2_X1 U964 ( .A(n1129), .B(n1134), .Z(n1222) );
NAND2_X1 U965 ( .A1(G224), .A2(n1044), .ZN(n1134) );
NAND2_X1 U966 ( .A1(n1226), .A2(n1227), .ZN(n1129) );
NAND2_X1 U967 ( .A1(n1228), .A2(n1059), .ZN(n1227) );
XOR2_X1 U968 ( .A(KEYINPUT57), .B(n1229), .Z(n1226) );
NOR2_X1 U969 ( .A1(n1059), .A2(n1228), .ZN(n1229) );
XNOR2_X1 U970 ( .A(KEYINPUT53), .B(n1054), .ZN(n1228) );
XOR2_X1 U971 ( .A(n1230), .B(n1231), .Z(n1054) );
XOR2_X1 U972 ( .A(G113), .B(n1232), .Z(n1231) );
NOR2_X1 U973 ( .A1(KEYINPUT2), .A2(n1233), .ZN(n1232) );
XOR2_X1 U974 ( .A(G116), .B(n1163), .Z(n1233) );
INV_X1 U975 ( .A(G119), .ZN(n1163) );
XOR2_X1 U976 ( .A(n1234), .B(n1213), .Z(n1230) );
XOR2_X1 U977 ( .A(G104), .B(G107), .Z(n1213) );
NAND2_X1 U978 ( .A1(KEYINPUT46), .A2(n1150), .ZN(n1234) );
INV_X1 U979 ( .A(G101), .ZN(n1150) );
INV_X1 U980 ( .A(n1053), .ZN(n1059) );
XNOR2_X1 U981 ( .A(n1235), .B(n1097), .ZN(n1053) );
XNOR2_X1 U982 ( .A(G110), .B(KEYINPUT39), .ZN(n1097) );
NOR2_X1 U983 ( .A1(n1141), .A2(n1020), .ZN(n981) );
XNOR2_X1 U984 ( .A(n1236), .B(G475), .ZN(n1020) );
NAND2_X1 U985 ( .A1(n1074), .A2(n1128), .ZN(n1236) );
INV_X1 U986 ( .A(G902), .ZN(n1128) );
XNOR2_X1 U987 ( .A(n1237), .B(n1238), .ZN(n1074) );
XOR2_X1 U988 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U989 ( .A(n1241), .B(n1242), .Z(n1240) );
AND2_X1 U990 ( .A1(G214), .A2(n1088), .ZN(n1242) );
AND2_X1 U991 ( .A1(n1243), .A2(n1044), .ZN(n1088) );
XOR2_X1 U992 ( .A(n1220), .B(KEYINPUT4), .Z(n1243) );
INV_X1 U993 ( .A(G237), .ZN(n1220) );
NAND2_X1 U994 ( .A1(n1244), .A2(n1245), .ZN(n1241) );
NAND4_X1 U995 ( .A1(KEYINPUT28), .A2(n1187), .A3(n1139), .A4(n1246), .ZN(n1245) );
NAND2_X1 U996 ( .A1(n1247), .A2(n1248), .ZN(n1244) );
NAND2_X1 U997 ( .A1(n1249), .A2(n1139), .ZN(n1248) );
INV_X1 U998 ( .A(G146), .ZN(n1139) );
OR2_X1 U999 ( .A1(n1187), .A2(KEYINPUT28), .ZN(n1249) );
NAND2_X1 U1000 ( .A1(n1187), .A2(n1246), .ZN(n1247) );
INV_X1 U1001 ( .A(KEYINPUT22), .ZN(n1246) );
XOR2_X1 U1002 ( .A(n1131), .B(n1043), .Z(n1187) );
INV_X1 U1003 ( .A(G140), .ZN(n1043) );
INV_X1 U1004 ( .A(G125), .ZN(n1131) );
NAND3_X1 U1005 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1239) );
NAND2_X1 U1006 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U1007 ( .A1(KEYINPUT29), .A2(n1255), .ZN(n1251) );
NAND2_X1 U1008 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U1009 ( .A(KEYINPUT24), .B(G113), .Z(n1257) );
NAND2_X1 U1010 ( .A1(n1258), .A2(n1259), .ZN(n1250) );
INV_X1 U1011 ( .A(KEYINPUT29), .ZN(n1259) );
NAND2_X1 U1012 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NAND2_X1 U1013 ( .A1(KEYINPUT24), .A2(n1254), .ZN(n1261) );
OR3_X1 U1014 ( .A1(n1253), .A2(KEYINPUT24), .A3(n1254), .ZN(n1260) );
INV_X1 U1015 ( .A(G113), .ZN(n1254) );
INV_X1 U1016 ( .A(n1256), .ZN(n1253) );
XOR2_X1 U1017 ( .A(n1235), .B(KEYINPUT17), .Z(n1256) );
XOR2_X1 U1018 ( .A(n1075), .B(n1262), .Z(n1237) );
XOR2_X1 U1019 ( .A(G143), .B(G131), .Z(n1262) );
INV_X1 U1020 ( .A(G104), .ZN(n1075) );
NAND2_X1 U1021 ( .A1(n1263), .A2(n1264), .ZN(n1141) );
NAND2_X1 U1022 ( .A1(G478), .A2(n1265), .ZN(n1264) );
OR3_X1 U1023 ( .A1(G902), .A2(KEYINPUT63), .A3(n1023), .ZN(n1265) );
NAND2_X1 U1024 ( .A1(n1013), .A2(n1266), .ZN(n1263) );
INV_X1 U1025 ( .A(KEYINPUT63), .ZN(n1266) );
NOR3_X1 U1026 ( .A1(G478), .A2(G902), .A3(n1023), .ZN(n1013) );
XNOR2_X1 U1027 ( .A(n1267), .B(n1268), .ZN(n1023) );
XOR2_X1 U1028 ( .A(n1269), .B(n1235), .Z(n1268) );
XNOR2_X1 U1029 ( .A(G122), .B(KEYINPUT61), .ZN(n1235) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1188), .ZN(n1269) );
AND2_X1 U1031 ( .A1(G234), .A2(n1044), .ZN(n1188) );
INV_X1 U1032 ( .A(G953), .ZN(n1044) );
XOR2_X1 U1033 ( .A(n1270), .B(n1271), .Z(n1267) );
NOR2_X1 U1034 ( .A1(KEYINPUT36), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U1035 ( .A(G134), .B(n1273), .ZN(n1272) );
NOR2_X1 U1036 ( .A1(KEYINPUT14), .A2(n1225), .ZN(n1273) );
XNOR2_X1 U1037 ( .A(G143), .B(G128), .ZN(n1225) );
XNOR2_X1 U1038 ( .A(G107), .B(G116), .ZN(n1270) );
endmodule


