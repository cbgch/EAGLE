//Key = 1100101111001001000111101100010101000011011111011110110101111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308;

XOR2_X1 U722 ( .A(n985), .B(n986), .Z(G9) );
NOR2_X1 U723 ( .A1(n987), .A2(n988), .ZN(n985) );
XOR2_X1 U724 ( .A(KEYINPUT44), .B(KEYINPUT38), .Z(n988) );
NOR2_X1 U725 ( .A1(n989), .A2(n990), .ZN(G75) );
NOR4_X1 U726 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
XOR2_X1 U727 ( .A(KEYINPUT37), .B(n995), .Z(n992) );
NOR3_X1 U728 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NAND3_X1 U729 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n996) );
NAND3_X1 U730 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n991) );
NAND2_X1 U731 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U732 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND3_X1 U733 ( .A1(n1000), .A2(n1009), .A3(n1010), .ZN(n1008) );
NAND2_X1 U734 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND3_X1 U735 ( .A1(n1013), .A2(n1001), .A3(KEYINPUT42), .ZN(n1012) );
NAND2_X1 U736 ( .A1(n1014), .A2(n1015), .ZN(n1011) );
NAND2_X1 U737 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U738 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U739 ( .A1(n1001), .A2(n1020), .ZN(n1007) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
OR4_X1 U741 ( .A1(n1023), .A2(n997), .A3(n1000), .A4(KEYINPUT42), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1014), .A2(n1024), .ZN(n1021) );
NAND2_X1 U743 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U744 ( .A1(n1010), .A2(n1027), .ZN(n1026) );
NAND2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1000), .A2(n1032), .ZN(n1025) );
NAND2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
INV_X1 U750 ( .A(n1037), .ZN(n1001) );
INV_X1 U751 ( .A(n998), .ZN(n1005) );
AND3_X1 U752 ( .A1(n1002), .A2(n1003), .A3(n1038), .ZN(n989) );
NAND4_X1 U753 ( .A1(n1039), .A2(n1010), .A3(n1040), .A4(n1041), .ZN(n1002) );
NOR3_X1 U754 ( .A1(n1037), .A2(n1042), .A3(n1043), .ZN(n1041) );
XOR2_X1 U755 ( .A(n1044), .B(KEYINPUT33), .Z(n1040) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XOR2_X1 U758 ( .A(KEYINPUT53), .B(n1049), .Z(n1045) );
NOR2_X1 U759 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
XNOR2_X1 U760 ( .A(KEYINPUT54), .B(G472), .ZN(n1047) );
INV_X1 U761 ( .A(n997), .ZN(n1010) );
XNOR2_X1 U762 ( .A(n1050), .B(KEYINPUT32), .ZN(n1039) );
XOR2_X1 U763 ( .A(n1051), .B(n1052), .Z(G72) );
XOR2_X1 U764 ( .A(n1053), .B(n1054), .Z(n1052) );
NAND2_X1 U765 ( .A1(G953), .A2(n1055), .ZN(n1054) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1055) );
NAND2_X1 U767 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND2_X1 U768 ( .A1(G953), .A2(n1058), .ZN(n1057) );
XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n1059), .ZN(n1058) );
XOR2_X1 U770 ( .A(n1060), .B(n1061), .Z(n1056) );
NOR2_X1 U771 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XOR2_X1 U772 ( .A(n1064), .B(KEYINPUT49), .Z(n1063) );
NAND2_X1 U773 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U774 ( .A1(n1066), .A2(n1065), .ZN(n1062) );
XNOR2_X1 U775 ( .A(n1067), .B(n1068), .ZN(n1065) );
XNOR2_X1 U776 ( .A(G131), .B(KEYINPUT5), .ZN(n1067) );
NAND2_X1 U777 ( .A1(KEYINPUT12), .A2(n1069), .ZN(n1060) );
XOR2_X1 U778 ( .A(G140), .B(G125), .Z(n1069) );
NOR2_X1 U779 ( .A1(n1070), .A2(G953), .ZN(n1051) );
XOR2_X1 U780 ( .A(n1071), .B(n1072), .Z(G69) );
NOR2_X1 U781 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U782 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NAND2_X1 U783 ( .A1(n1077), .A2(n1003), .ZN(n1076) );
NAND2_X1 U784 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
OR2_X1 U785 ( .A1(n1080), .A2(n1033), .ZN(n1079) );
NAND2_X1 U786 ( .A1(n1081), .A2(G953), .ZN(n1075) );
XOR2_X1 U787 ( .A(KEYINPUT22), .B(n1082), .Z(n1081) );
AND2_X1 U788 ( .A1(G224), .A2(G898), .ZN(n1082) );
NOR2_X1 U789 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U790 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND3_X1 U791 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
OR2_X1 U792 ( .A1(n1090), .A2(KEYINPUT30), .ZN(n1088) );
NAND2_X1 U793 ( .A1(KEYINPUT30), .A2(n1091), .ZN(n1087) );
NAND2_X1 U794 ( .A1(n1092), .A2(G902), .ZN(n1091) );
NOR2_X1 U795 ( .A1(n1083), .A2(n1093), .ZN(G63) );
XOR2_X1 U796 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U797 ( .A1(n1090), .A2(G478), .ZN(n1094) );
NOR2_X1 U798 ( .A1(n1083), .A2(n1096), .ZN(G60) );
XNOR2_X1 U799 ( .A(n1097), .B(n1098), .ZN(n1096) );
NOR3_X1 U800 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
NOR2_X1 U801 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U802 ( .A(KEYINPUT10), .ZN(n1103) );
NOR2_X1 U803 ( .A1(G902), .A2(n1092), .ZN(n1102) );
NOR2_X1 U804 ( .A1(KEYINPUT10), .A2(n1090), .ZN(n1100) );
XNOR2_X1 U805 ( .A(n1104), .B(n1105), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1106), .A2(n1023), .ZN(n1105) );
NOR3_X1 U807 ( .A1(n1083), .A2(n1107), .A3(n1108), .ZN(G57) );
NOR2_X1 U808 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U809 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
AND2_X1 U810 ( .A1(n1113), .A2(KEYINPUT35), .ZN(n1112) );
NOR3_X1 U811 ( .A1(KEYINPUT35), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR2_X1 U812 ( .A1(n1115), .A2(n1116), .ZN(n1107) );
INV_X1 U813 ( .A(n1109), .ZN(n1116) );
XNOR2_X1 U814 ( .A(n1117), .B(n1118), .ZN(n1109) );
NOR3_X1 U815 ( .A1(n1119), .A2(KEYINPUT3), .A3(n1120), .ZN(n1118) );
INV_X1 U816 ( .A(n1090), .ZN(n1119) );
NAND2_X1 U817 ( .A1(n1121), .A2(n1122), .ZN(n1117) );
NAND2_X1 U818 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U819 ( .A(n1125), .B(KEYINPUT51), .Z(n1121) );
OR2_X1 U820 ( .A1(n1124), .A2(n1123), .ZN(n1125) );
XNOR2_X1 U821 ( .A(n1126), .B(n1127), .ZN(n1124) );
NAND2_X1 U822 ( .A1(KEYINPUT52), .A2(n1128), .ZN(n1126) );
NOR2_X1 U823 ( .A1(n1113), .A2(n1114), .ZN(n1115) );
INV_X1 U824 ( .A(KEYINPUT45), .ZN(n1114) );
XNOR2_X1 U825 ( .A(n1129), .B(KEYINPUT15), .ZN(n1113) );
NOR2_X1 U826 ( .A1(n1083), .A2(n1130), .ZN(G54) );
XOR2_X1 U827 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U828 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U829 ( .A1(n1090), .A2(G469), .ZN(n1134) );
NAND2_X1 U830 ( .A1(n1135), .A2(KEYINPUT20), .ZN(n1133) );
XNOR2_X1 U831 ( .A(n1136), .B(KEYINPUT62), .ZN(n1135) );
XOR2_X1 U832 ( .A(KEYINPUT39), .B(n1137), .Z(n1131) );
NOR2_X1 U833 ( .A1(n1083), .A2(n1138), .ZN(G51) );
NOR2_X1 U834 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U835 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U836 ( .A1(KEYINPUT6), .A2(n1143), .ZN(n1142) );
NAND2_X1 U837 ( .A1(n1090), .A2(n1144), .ZN(n1141) );
NOR2_X1 U838 ( .A1(n1145), .A2(n1092), .ZN(n1090) );
AND2_X1 U839 ( .A1(n1070), .A2(n1146), .ZN(n1092) );
XNOR2_X1 U840 ( .A(KEYINPUT11), .B(n993), .ZN(n1146) );
NAND2_X1 U841 ( .A1(n1078), .A2(n1147), .ZN(n993) );
XOR2_X1 U842 ( .A(KEYINPUT4), .B(n1148), .Z(n1147) );
NOR2_X1 U843 ( .A1(n1033), .A2(n1080), .ZN(n1148) );
AND4_X1 U844 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1078) );
NOR4_X1 U845 ( .A1(n986), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1152) );
INV_X1 U846 ( .A(n1156), .ZN(n1154) );
NOR2_X1 U847 ( .A1(n1157), .A2(n1106), .ZN(n986) );
NAND3_X1 U848 ( .A1(n1000), .A2(n1158), .A3(n1159), .ZN(n1106) );
INV_X1 U849 ( .A(n999), .ZN(n1157) );
NAND4_X1 U850 ( .A1(n1013), .A2(n1159), .A3(n1000), .A4(n1160), .ZN(n1151) );
XNOR2_X1 U851 ( .A(KEYINPUT41), .B(n1158), .ZN(n1160) );
NAND3_X1 U852 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1149) );
XNOR2_X1 U853 ( .A(KEYINPUT43), .B(n1158), .ZN(n1162) );
INV_X1 U854 ( .A(n994), .ZN(n1070) );
NAND4_X1 U855 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n994) );
AND4_X1 U856 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR3_X1 U857 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1166) );
NOR2_X1 U858 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
INV_X1 U859 ( .A(KEYINPUT58), .ZN(n1175) );
NOR2_X1 U860 ( .A1(KEYINPUT58), .A2(n1177), .ZN(n1173) );
NAND4_X1 U861 ( .A1(n1178), .A2(n1179), .A3(n1013), .A4(n1180), .ZN(n1177) );
NOR3_X1 U862 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NOR2_X1 U863 ( .A1(KEYINPUT6), .A2(n1143), .ZN(n1139) );
XNOR2_X1 U864 ( .A(n1184), .B(n1185), .ZN(n1143) );
AND2_X1 U865 ( .A1(n1186), .A2(n1038), .ZN(n1083) );
INV_X1 U866 ( .A(G952), .ZN(n1038) );
XNOR2_X1 U867 ( .A(G953), .B(KEYINPUT55), .ZN(n1186) );
XNOR2_X1 U868 ( .A(G146), .B(n1176), .ZN(G48) );
NAND2_X1 U869 ( .A1(n1187), .A2(n1013), .ZN(n1176) );
NAND2_X1 U870 ( .A1(n1188), .A2(n1189), .ZN(G45) );
NAND2_X1 U871 ( .A1(G143), .A2(n1190), .ZN(n1189) );
XOR2_X1 U872 ( .A(n1191), .B(KEYINPUT40), .Z(n1188) );
NAND2_X1 U873 ( .A1(n1172), .A2(n1192), .ZN(n1191) );
INV_X1 U874 ( .A(n1190), .ZN(n1172) );
NAND3_X1 U875 ( .A1(n1193), .A2(n1159), .A3(n1194), .ZN(n1190) );
NOR3_X1 U876 ( .A1(n1195), .A2(n1183), .A3(n1196), .ZN(n1194) );
XNOR2_X1 U877 ( .A(G140), .B(n1164), .ZN(G42) );
NAND2_X1 U878 ( .A1(n1197), .A2(n1198), .ZN(n1164) );
XNOR2_X1 U879 ( .A(G137), .B(n1165), .ZN(G39) );
NAND3_X1 U880 ( .A1(n1197), .A2(n1179), .A3(n1199), .ZN(n1165) );
XNOR2_X1 U881 ( .A(G134), .B(n1171), .ZN(G36) );
NAND3_X1 U882 ( .A1(n1193), .A2(n999), .A3(n1197), .ZN(n1171) );
XNOR2_X1 U883 ( .A(G131), .B(n1170), .ZN(G33) );
NAND2_X1 U884 ( .A1(n1197), .A2(n1163), .ZN(n1170) );
NOR3_X1 U885 ( .A1(n1016), .A2(n1183), .A3(n997), .ZN(n1197) );
NAND2_X1 U886 ( .A1(n1036), .A2(n1200), .ZN(n997) );
INV_X1 U887 ( .A(n1201), .ZN(n1183) );
XNOR2_X1 U888 ( .A(G128), .B(n1169), .ZN(G30) );
NAND2_X1 U889 ( .A1(n1187), .A2(n999), .ZN(n1169) );
AND4_X1 U890 ( .A1(n1030), .A2(n1159), .A3(n1179), .A4(n1201), .ZN(n1187) );
XOR2_X1 U891 ( .A(G101), .B(n1202), .Z(G3) );
NOR3_X1 U892 ( .A1(n1203), .A2(KEYINPUT2), .A3(n1033), .ZN(n1202) );
XNOR2_X1 U893 ( .A(KEYINPUT8), .B(n1080), .ZN(n1203) );
NAND4_X1 U894 ( .A1(n1014), .A2(n1193), .A3(n1182), .A4(n1158), .ZN(n1080) );
XNOR2_X1 U895 ( .A(G125), .B(n1168), .ZN(G27) );
NAND3_X1 U896 ( .A1(n1161), .A2(n1201), .A3(n1198), .ZN(n1168) );
NOR3_X1 U897 ( .A1(n1179), .A2(n1181), .A3(n1023), .ZN(n1198) );
NAND2_X1 U898 ( .A1(n998), .A2(n1204), .ZN(n1201) );
NAND4_X1 U899 ( .A1(G902), .A2(G953), .A3(n1205), .A4(n1059), .ZN(n1204) );
INV_X1 U900 ( .A(G900), .ZN(n1059) );
XNOR2_X1 U901 ( .A(G122), .B(n1150), .ZN(G24) );
NAND4_X1 U902 ( .A1(n1206), .A2(n1000), .A3(n1050), .A4(n1043), .ZN(n1150) );
AND2_X1 U903 ( .A1(n1207), .A2(n1181), .ZN(n1000) );
XNOR2_X1 U904 ( .A(KEYINPUT1), .B(n1031), .ZN(n1207) );
XOR2_X1 U905 ( .A(G119), .B(n1155), .Z(G21) );
AND3_X1 U906 ( .A1(n1199), .A2(n1179), .A3(n1206), .ZN(n1155) );
XNOR2_X1 U907 ( .A(G116), .B(n1156), .ZN(G18) );
NAND3_X1 U908 ( .A1(n1193), .A2(n999), .A3(n1206), .ZN(n1156) );
NOR2_X1 U909 ( .A1(n1043), .A2(n1195), .ZN(n999) );
INV_X1 U910 ( .A(n1050), .ZN(n1195) );
INV_X1 U911 ( .A(n1028), .ZN(n1193) );
XOR2_X1 U912 ( .A(n1208), .B(n1209), .Z(G15) );
NOR2_X1 U913 ( .A1(G113), .A2(KEYINPUT14), .ZN(n1209) );
NAND2_X1 U914 ( .A1(n1206), .A2(n1163), .ZN(n1208) );
NOR2_X1 U915 ( .A1(n1028), .A2(n1023), .ZN(n1163) );
INV_X1 U916 ( .A(n1013), .ZN(n1023) );
NOR2_X1 U917 ( .A1(n1050), .A2(n1196), .ZN(n1013) );
INV_X1 U918 ( .A(n1043), .ZN(n1196) );
NAND2_X1 U919 ( .A1(n1210), .A2(n1179), .ZN(n1028) );
INV_X1 U920 ( .A(n1031), .ZN(n1179) );
XNOR2_X1 U921 ( .A(KEYINPUT56), .B(n1030), .ZN(n1210) );
AND2_X1 U922 ( .A1(n1161), .A2(n1158), .ZN(n1206) );
NOR2_X1 U923 ( .A1(n1037), .A2(n1033), .ZN(n1161) );
NAND2_X1 U924 ( .A1(n1019), .A2(n1211), .ZN(n1037) );
XNOR2_X1 U925 ( .A(n1153), .B(n1212), .ZN(G12) );
XNOR2_X1 U926 ( .A(KEYINPUT47), .B(n1213), .ZN(n1212) );
AND4_X1 U927 ( .A1(n1199), .A2(n1159), .A3(n1031), .A4(n1158), .ZN(n1153) );
NAND2_X1 U928 ( .A1(n998), .A2(n1214), .ZN(n1158) );
NAND3_X1 U929 ( .A1(n1073), .A2(n1205), .A3(G902), .ZN(n1214) );
NOR2_X1 U930 ( .A1(n1003), .A2(G898), .ZN(n1073) );
NAND3_X1 U931 ( .A1(n1205), .A2(n1003), .A3(G952), .ZN(n998) );
NAND2_X1 U932 ( .A1(G237), .A2(G234), .ZN(n1205) );
XOR2_X1 U933 ( .A(n1048), .B(n1120), .Z(n1031) );
INV_X1 U934 ( .A(G472), .ZN(n1120) );
AND2_X1 U935 ( .A1(n1215), .A2(n1145), .ZN(n1048) );
XOR2_X1 U936 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U937 ( .A(n1123), .B(n1127), .Z(n1217) );
XOR2_X1 U938 ( .A(G146), .B(n1218), .Z(n1127) );
XOR2_X1 U939 ( .A(n1219), .B(n1220), .Z(n1123) );
NAND2_X1 U940 ( .A1(KEYINPUT48), .A2(n1221), .ZN(n1219) );
XNOR2_X1 U941 ( .A(n1128), .B(n1222), .ZN(n1216) );
NOR2_X1 U942 ( .A1(KEYINPUT46), .A2(n1129), .ZN(n1222) );
XNOR2_X1 U943 ( .A(n1223), .B(G101), .ZN(n1129) );
NAND2_X1 U944 ( .A1(G210), .A2(n1224), .ZN(n1223) );
NOR2_X1 U945 ( .A1(n1033), .A2(n1016), .ZN(n1159) );
INV_X1 U946 ( .A(n1182), .ZN(n1016) );
NOR2_X1 U947 ( .A1(n1019), .A2(n1018), .ZN(n1182) );
INV_X1 U948 ( .A(n1211), .ZN(n1018) );
NAND2_X1 U949 ( .A1(G221), .A2(n1225), .ZN(n1211) );
XOR2_X1 U950 ( .A(n1226), .B(G469), .Z(n1019) );
NAND2_X1 U951 ( .A1(n1227), .A2(n1145), .ZN(n1226) );
XOR2_X1 U952 ( .A(n1228), .B(n1137), .Z(n1227) );
AND2_X1 U953 ( .A1(n1229), .A2(n1230), .ZN(n1137) );
NAND3_X1 U954 ( .A1(n1231), .A2(G227), .A3(n1232), .ZN(n1230) );
XNOR2_X1 U955 ( .A(G110), .B(G140), .ZN(n1232) );
NAND2_X1 U956 ( .A1(n1233), .A2(n1234), .ZN(n1229) );
NAND2_X1 U957 ( .A1(n1231), .A2(G227), .ZN(n1234) );
XNOR2_X1 U958 ( .A(KEYINPUT34), .B(G953), .ZN(n1231) );
XNOR2_X1 U959 ( .A(G140), .B(n1213), .ZN(n1233) );
INV_X1 U960 ( .A(G110), .ZN(n1213) );
NAND2_X1 U961 ( .A1(KEYINPUT0), .A2(n1136), .ZN(n1228) );
XNOR2_X1 U962 ( .A(n1235), .B(n1236), .ZN(n1136) );
XNOR2_X1 U963 ( .A(n1237), .B(n1128), .ZN(n1236) );
XOR2_X1 U964 ( .A(n1068), .B(n1238), .Z(n1128) );
XNOR2_X1 U965 ( .A(n1239), .B(KEYINPUT60), .ZN(n1238) );
NAND2_X1 U966 ( .A1(KEYINPUT25), .A2(n1240), .ZN(n1239) );
INV_X1 U967 ( .A(G131), .ZN(n1240) );
XOR2_X1 U968 ( .A(G134), .B(G137), .Z(n1068) );
NAND2_X1 U969 ( .A1(KEYINPUT50), .A2(n1241), .ZN(n1237) );
XNOR2_X1 U970 ( .A(n1104), .B(n1242), .ZN(n1241) );
XNOR2_X1 U971 ( .A(KEYINPUT9), .B(n987), .ZN(n1242) );
XNOR2_X1 U972 ( .A(n1066), .B(n1243), .ZN(n1235) );
XNOR2_X1 U973 ( .A(n1244), .B(n1245), .ZN(n1066) );
XOR2_X1 U974 ( .A(KEYINPUT24), .B(G146), .Z(n1245) );
XOR2_X1 U975 ( .A(n1246), .B(G128), .Z(n1244) );
NAND2_X1 U976 ( .A1(KEYINPUT31), .A2(n1192), .ZN(n1246) );
INV_X1 U977 ( .A(n1178), .ZN(n1033) );
NOR2_X1 U978 ( .A1(n1036), .A2(n1035), .ZN(n1178) );
INV_X1 U979 ( .A(n1200), .ZN(n1035) );
NAND2_X1 U980 ( .A1(n1247), .A2(n1248), .ZN(n1200) );
XOR2_X1 U981 ( .A(KEYINPUT16), .B(G214), .Z(n1247) );
XOR2_X1 U982 ( .A(n1249), .B(n1144), .Z(n1036) );
AND2_X1 U983 ( .A1(G210), .A2(n1248), .ZN(n1144) );
OR2_X1 U984 ( .A1(G902), .A2(G237), .ZN(n1248) );
NAND2_X1 U985 ( .A1(n1250), .A2(n1145), .ZN(n1249) );
XNOR2_X1 U986 ( .A(n1251), .B(n1252), .ZN(n1250) );
INV_X1 U987 ( .A(n1184), .ZN(n1252) );
XNOR2_X1 U988 ( .A(n1074), .B(n1253), .ZN(n1184) );
XOR2_X1 U989 ( .A(n1254), .B(n1218), .Z(n1253) );
XOR2_X1 U990 ( .A(n1255), .B(n1256), .Z(n1074) );
XOR2_X1 U991 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U992 ( .A(n1221), .B(G110), .ZN(n1258) );
INV_X1 U993 ( .A(G116), .ZN(n1221) );
XNOR2_X1 U994 ( .A(KEYINPUT13), .B(n1259), .ZN(n1257) );
XOR2_X1 U995 ( .A(n1260), .B(n1261), .Z(n1255) );
XOR2_X1 U996 ( .A(n1220), .B(n1243), .Z(n1261) );
XOR2_X1 U997 ( .A(G101), .B(KEYINPUT59), .Z(n1243) );
XOR2_X1 U998 ( .A(G113), .B(G119), .Z(n1220) );
XNOR2_X1 U999 ( .A(G107), .B(n1262), .ZN(n1260) );
NOR2_X1 U1000 ( .A1(KEYINPUT28), .A2(n1104), .ZN(n1262) );
NAND2_X1 U1001 ( .A1(KEYINPUT19), .A2(n1185), .ZN(n1251) );
AND2_X1 U1002 ( .A1(G224), .A2(n1003), .ZN(n1185) );
AND2_X1 U1003 ( .A1(n1014), .A2(n1030), .ZN(n1199) );
INV_X1 U1004 ( .A(n1181), .ZN(n1030) );
XOR2_X1 U1005 ( .A(n1042), .B(KEYINPUT57), .Z(n1181) );
XOR2_X1 U1006 ( .A(n1089), .B(n1263), .Z(n1042) );
AND2_X1 U1007 ( .A1(n1145), .A2(n1086), .ZN(n1263) );
XNOR2_X1 U1008 ( .A(n1264), .B(n1265), .ZN(n1086) );
NOR2_X1 U1009 ( .A1(KEYINPUT26), .A2(n1266), .ZN(n1265) );
XOR2_X1 U1010 ( .A(n1267), .B(G137), .Z(n1266) );
NAND2_X1 U1011 ( .A1(G221), .A2(n1268), .ZN(n1267) );
NAND3_X1 U1012 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1264) );
NAND2_X1 U1013 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
OR3_X1 U1014 ( .A1(n1273), .A2(n1272), .A3(KEYINPUT18), .ZN(n1270) );
XNOR2_X1 U1015 ( .A(n1274), .B(KEYINPUT29), .ZN(n1272) );
OR2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1275), .ZN(n1273) );
NAND2_X1 U1017 ( .A1(KEYINPUT18), .A2(n1275), .ZN(n1269) );
XNOR2_X1 U1018 ( .A(G110), .B(n1276), .ZN(n1275) );
XOR2_X1 U1019 ( .A(G128), .B(G119), .Z(n1276) );
AND2_X1 U1020 ( .A1(G217), .A2(n1225), .ZN(n1089) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1145), .ZN(n1225) );
NOR2_X1 U1022 ( .A1(n1050), .A2(n1043), .ZN(n1014) );
XOR2_X1 U1023 ( .A(n1277), .B(n1099), .Z(n1043) );
INV_X1 U1024 ( .A(G475), .ZN(n1099) );
NAND2_X1 U1025 ( .A1(n1145), .A2(n1098), .ZN(n1277) );
NAND3_X1 U1026 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1098) );
OR2_X1 U1027 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U1028 ( .A1(n1283), .A2(n1284), .ZN(n1279) );
INV_X1 U1029 ( .A(KEYINPUT63), .ZN(n1284) );
NAND2_X1 U1030 ( .A1(n1285), .A2(n1281), .ZN(n1283) );
XNOR2_X1 U1031 ( .A(KEYINPUT36), .B(n1286), .ZN(n1285) );
NAND2_X1 U1032 ( .A1(KEYINPUT63), .A2(n1287), .ZN(n1278) );
NAND2_X1 U1033 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND3_X1 U1034 ( .A1(n1282), .A2(n1281), .A3(n1290), .ZN(n1289) );
INV_X1 U1035 ( .A(KEYINPUT36), .ZN(n1290) );
XNOR2_X1 U1036 ( .A(n1291), .B(n1292), .ZN(n1281) );
XNOR2_X1 U1037 ( .A(G113), .B(n1104), .ZN(n1292) );
INV_X1 U1038 ( .A(G104), .ZN(n1104) );
NAND2_X1 U1039 ( .A1(KEYINPUT7), .A2(n1259), .ZN(n1291) );
NAND2_X1 U1040 ( .A1(KEYINPUT36), .A2(n1286), .ZN(n1288) );
INV_X1 U1041 ( .A(n1282), .ZN(n1286) );
XNOR2_X1 U1042 ( .A(n1293), .B(n1294), .ZN(n1282) );
XNOR2_X1 U1043 ( .A(n1192), .B(G131), .ZN(n1294) );
XOR2_X1 U1044 ( .A(n1274), .B(n1295), .Z(n1293) );
AND2_X1 U1045 ( .A1(n1224), .A2(G214), .ZN(n1295) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1224) );
XNOR2_X1 U1047 ( .A(G140), .B(n1254), .ZN(n1274) );
XOR2_X1 U1048 ( .A(G125), .B(G146), .Z(n1254) );
XNOR2_X1 U1049 ( .A(n1296), .B(G478), .ZN(n1050) );
NAND2_X1 U1050 ( .A1(n1095), .A2(n1145), .ZN(n1296) );
INV_X1 U1051 ( .A(G902), .ZN(n1145) );
XNOR2_X1 U1052 ( .A(n1297), .B(n1298), .ZN(n1095) );
XNOR2_X1 U1053 ( .A(n1299), .B(n1218), .ZN(n1298) );
XNOR2_X1 U1054 ( .A(G128), .B(n1192), .ZN(n1218) );
INV_X1 U1055 ( .A(G143), .ZN(n1192) );
NAND2_X1 U1056 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U1057 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U1058 ( .A(KEYINPUT23), .B(n987), .ZN(n1303) );
INV_X1 U1059 ( .A(G107), .ZN(n987) );
XNOR2_X1 U1060 ( .A(G122), .B(n1304), .ZN(n1302) );
XOR2_X1 U1061 ( .A(n1305), .B(KEYINPUT61), .Z(n1300) );
NAND2_X1 U1062 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U1063 ( .A(n1259), .B(n1304), .ZN(n1307) );
NOR2_X1 U1064 ( .A1(G116), .A2(KEYINPUT17), .ZN(n1304) );
INV_X1 U1065 ( .A(G122), .ZN(n1259) );
XNOR2_X1 U1066 ( .A(KEYINPUT23), .B(G107), .ZN(n1306) );
XOR2_X1 U1067 ( .A(n1308), .B(G134), .Z(n1297) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1268), .ZN(n1308) );
AND2_X1 U1069 ( .A1(G234), .A2(n1003), .ZN(n1268) );
INV_X1 U1070 ( .A(G953), .ZN(n1003) );
endmodule


