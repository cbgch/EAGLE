//Key = 0010100001101001101111011000011101000011000100000111000100011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215;

NAND2_X1 U683 ( .A1(n925), .A2(n926), .ZN(G9) );
NAND2_X1 U684 ( .A1(G107), .A2(n927), .ZN(n926) );
XOR2_X1 U685 ( .A(n928), .B(KEYINPUT54), .Z(n925) );
NAND2_X1 U686 ( .A1(n929), .A2(n930), .ZN(n928) );
NOR2_X1 U687 ( .A1(n931), .A2(n932), .ZN(G75) );
NOR4_X1 U688 ( .A1(G953), .A2(n933), .A3(n934), .A4(n935), .ZN(n932) );
NOR2_X1 U689 ( .A1(n936), .A2(n937), .ZN(n934) );
NOR2_X1 U690 ( .A1(n938), .A2(n939), .ZN(n937) );
NOR3_X1 U691 ( .A1(n940), .A2(n941), .A3(n942), .ZN(n939) );
NOR2_X1 U692 ( .A1(n943), .A2(n944), .ZN(n941) );
AND2_X1 U693 ( .A1(n945), .A2(n946), .ZN(n944) );
NOR3_X1 U694 ( .A1(n947), .A2(n948), .A3(n949), .ZN(n943) );
NOR3_X1 U695 ( .A1(n950), .A2(n951), .A3(n952), .ZN(n949) );
NOR2_X1 U696 ( .A1(n946), .A2(n953), .ZN(n948) );
NOR4_X1 U697 ( .A1(n950), .A2(n954), .A3(n955), .A4(n947), .ZN(n938) );
INV_X1 U698 ( .A(n956), .ZN(n947) );
INV_X1 U699 ( .A(n946), .ZN(n955) );
NOR2_X1 U700 ( .A1(n957), .A2(n958), .ZN(n954) );
NOR2_X1 U701 ( .A1(n959), .A2(n940), .ZN(n958) );
INV_X1 U702 ( .A(n960), .ZN(n940) );
NOR2_X1 U703 ( .A1(n961), .A2(n962), .ZN(n959) );
NOR2_X1 U704 ( .A1(n963), .A2(n942), .ZN(n957) );
NOR2_X1 U705 ( .A1(n964), .A2(n965), .ZN(n963) );
AND3_X1 U706 ( .A1(n966), .A2(n967), .A3(G221), .ZN(n964) );
NOR3_X1 U707 ( .A1(n933), .A2(G953), .A3(G952), .ZN(n931) );
AND4_X1 U708 ( .A1(n956), .A2(n953), .A3(n960), .A4(n968), .ZN(n933) );
NOR4_X1 U709 ( .A1(n969), .A2(n970), .A3(n971), .A4(n972), .ZN(n968) );
XOR2_X1 U710 ( .A(KEYINPUT5), .B(n973), .Z(n972) );
XOR2_X1 U711 ( .A(n974), .B(KEYINPUT0), .Z(n971) );
NAND2_X1 U712 ( .A1(n975), .A2(n976), .ZN(n974) );
NAND2_X1 U713 ( .A1(n977), .A2(n978), .ZN(n976) );
XOR2_X1 U714 ( .A(KEYINPUT13), .B(n979), .Z(n977) );
NAND2_X1 U715 ( .A1(n980), .A2(G475), .ZN(n975) );
XOR2_X1 U716 ( .A(KEYINPUT4), .B(n979), .Z(n980) );
AND2_X1 U717 ( .A1(n981), .A2(KEYINPUT48), .ZN(n970) );
NOR2_X1 U718 ( .A1(KEYINPUT48), .A2(n982), .ZN(n969) );
XOR2_X1 U719 ( .A(n983), .B(n984), .Z(G72) );
NOR2_X1 U720 ( .A1(n985), .A2(n986), .ZN(n984) );
NOR3_X1 U721 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
XOR2_X1 U722 ( .A(n990), .B(KEYINPUT38), .Z(n989) );
NOR2_X1 U723 ( .A1(n991), .A2(n992), .ZN(n988) );
XOR2_X1 U724 ( .A(n993), .B(KEYINPUT15), .Z(n991) );
NOR2_X1 U725 ( .A1(n994), .A2(n990), .ZN(n985) );
NAND2_X1 U726 ( .A1(n995), .A2(n992), .ZN(n990) );
NAND2_X1 U727 ( .A1(n996), .A2(n997), .ZN(n995) );
INV_X1 U728 ( .A(n987), .ZN(n994) );
XOR2_X1 U729 ( .A(n998), .B(n999), .Z(n987) );
XOR2_X1 U730 ( .A(n1000), .B(n1001), .Z(n999) );
XOR2_X1 U731 ( .A(n1002), .B(n1003), .Z(n998) );
XOR2_X1 U732 ( .A(G137), .B(G134), .Z(n1003) );
NAND2_X1 U733 ( .A1(G953), .A2(n1004), .ZN(n983) );
NAND2_X1 U734 ( .A1(G900), .A2(G227), .ZN(n1004) );
NAND3_X1 U735 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(G69) );
XOR2_X1 U736 ( .A(n1008), .B(KEYINPUT32), .Z(n1007) );
OR2_X1 U737 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U738 ( .A1(n1010), .A2(n1009), .ZN(n1006) );
NAND2_X1 U739 ( .A1(G953), .A2(n1011), .ZN(n1009) );
NAND2_X1 U740 ( .A1(G898), .A2(G224), .ZN(n1011) );
NOR2_X1 U741 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
XOR2_X1 U742 ( .A(n1014), .B(KEYINPUT53), .Z(n1012) );
NAND2_X1 U743 ( .A1(n1014), .A2(n1013), .ZN(n1005) );
NAND2_X1 U744 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
XOR2_X1 U745 ( .A(KEYINPUT33), .B(n1017), .Z(n1016) );
NOR2_X1 U746 ( .A1(G898), .A2(n992), .ZN(n1017) );
XOR2_X1 U747 ( .A(KEYINPUT10), .B(n1018), .Z(n1015) );
INV_X1 U748 ( .A(n1019), .ZN(n1018) );
NOR2_X1 U749 ( .A1(G953), .A2(n1020), .ZN(n1014) );
NOR2_X1 U750 ( .A1(n1021), .A2(n1022), .ZN(G66) );
XOR2_X1 U751 ( .A(n1023), .B(n1024), .Z(n1022) );
NOR2_X1 U752 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U753 ( .A1(n1021), .A2(n1027), .ZN(G63) );
XOR2_X1 U754 ( .A(n1028), .B(n1029), .Z(n1027) );
AND2_X1 U755 ( .A1(G478), .A2(n1030), .ZN(n1028) );
NOR2_X1 U756 ( .A1(n1021), .A2(n1031), .ZN(G60) );
XOR2_X1 U757 ( .A(n1032), .B(n1033), .Z(n1031) );
NAND2_X1 U758 ( .A1(KEYINPUT50), .A2(n1034), .ZN(n1032) );
NAND2_X1 U759 ( .A1(n1030), .A2(G475), .ZN(n1034) );
XOR2_X1 U760 ( .A(n1035), .B(n1036), .Z(G6) );
NOR2_X1 U761 ( .A1(n1021), .A2(n1037), .ZN(G57) );
XOR2_X1 U762 ( .A(n1038), .B(n1039), .Z(n1037) );
XOR2_X1 U763 ( .A(n1040), .B(n1041), .Z(n1039) );
NAND4_X1 U764 ( .A1(KEYINPUT20), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1041) );
OR3_X1 U765 ( .A1(n1045), .A2(KEYINPUT17), .A3(G101), .ZN(n1044) );
NAND2_X1 U766 ( .A1(G101), .A2(n1045), .ZN(n1043) );
NAND2_X1 U767 ( .A1(KEYINPUT63), .A2(n1046), .ZN(n1045) );
NAND2_X1 U768 ( .A1(KEYINPUT17), .A2(n1047), .ZN(n1042) );
INV_X1 U769 ( .A(n1046), .ZN(n1047) );
XNOR2_X1 U770 ( .A(n1048), .B(KEYINPUT1), .ZN(n1046) );
NAND2_X1 U771 ( .A1(n1049), .A2(n1050), .ZN(n1040) );
NAND2_X1 U772 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U773 ( .A(n1053), .B(KEYINPUT27), .Z(n1049) );
OR2_X1 U774 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
AND2_X1 U775 ( .A1(G472), .A2(n1030), .ZN(n1038) );
NOR2_X1 U776 ( .A1(n1021), .A2(n1054), .ZN(G54) );
XOR2_X1 U777 ( .A(n1055), .B(n1056), .Z(n1054) );
XNOR2_X1 U778 ( .A(n1057), .B(KEYINPUT23), .ZN(n1056) );
NAND3_X1 U779 ( .A1(n1030), .A2(G469), .A3(KEYINPUT31), .ZN(n1057) );
INV_X1 U780 ( .A(n1026), .ZN(n1030) );
NOR2_X1 U781 ( .A1(n1021), .A2(n1058), .ZN(G51) );
XOR2_X1 U782 ( .A(n1019), .B(n1059), .Z(n1058) );
XOR2_X1 U783 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR3_X1 U784 ( .A1(n1026), .A2(n1062), .A3(n1063), .ZN(n1061) );
NAND2_X1 U785 ( .A1(G902), .A2(n935), .ZN(n1026) );
NAND3_X1 U786 ( .A1(n996), .A2(n1064), .A3(n1020), .ZN(n935) );
AND4_X1 U787 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1020) );
AND4_X1 U788 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1036), .ZN(n1068) );
NAND3_X1 U789 ( .A1(n1072), .A2(n982), .A3(n951), .ZN(n1036) );
NOR2_X1 U790 ( .A1(n1073), .A2(n929), .ZN(n1067) );
INV_X1 U791 ( .A(n927), .ZN(n929) );
NAND3_X1 U792 ( .A1(n952), .A2(n982), .A3(n1072), .ZN(n927) );
XOR2_X1 U793 ( .A(KEYINPUT34), .B(n997), .Z(n1064) );
AND4_X1 U794 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n997) );
AND4_X1 U795 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n996) );
NAND2_X1 U796 ( .A1(KEYINPUT21), .A2(n1082), .ZN(n1060) );
INV_X1 U797 ( .A(n1083), .ZN(n1082) );
NOR2_X1 U798 ( .A1(n992), .A2(G952), .ZN(n1021) );
XNOR2_X1 U799 ( .A(G146), .B(n1078), .ZN(G48) );
NAND4_X1 U800 ( .A1(n965), .A2(n1084), .A3(n951), .A4(n1085), .ZN(n1078) );
XOR2_X1 U801 ( .A(n1086), .B(G143), .Z(G45) );
NAND2_X1 U802 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U803 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
OR2_X1 U804 ( .A1(n1079), .A2(n1091), .ZN(n1087) );
INV_X1 U805 ( .A(KEYINPUT18), .ZN(n1091) );
NAND2_X1 U806 ( .A1(n1089), .A2(n1092), .ZN(n1079) );
AND4_X1 U807 ( .A1(n965), .A2(n961), .A3(n945), .A4(n1085), .ZN(n1089) );
XNOR2_X1 U808 ( .A(G140), .B(n1080), .ZN(G42) );
NAND3_X1 U809 ( .A1(n951), .A2(n962), .A3(n1093), .ZN(n1080) );
XOR2_X1 U810 ( .A(n1081), .B(n1094), .Z(G39) );
NOR2_X1 U811 ( .A1(G137), .A2(KEYINPUT6), .ZN(n1094) );
NAND4_X1 U812 ( .A1(n1095), .A2(n1093), .A3(n946), .A4(n1096), .ZN(n1081) );
XOR2_X1 U813 ( .A(n1097), .B(n1074), .Z(G36) );
NAND3_X1 U814 ( .A1(n961), .A2(n952), .A3(n1093), .ZN(n1074) );
XNOR2_X1 U815 ( .A(G131), .B(n1075), .ZN(G33) );
NAND3_X1 U816 ( .A1(n961), .A2(n951), .A3(n1093), .ZN(n1075) );
AND4_X1 U817 ( .A1(n965), .A2(n956), .A3(n1085), .A4(n953), .ZN(n1093) );
XNOR2_X1 U818 ( .A(n1098), .B(KEYINPUT29), .ZN(n965) );
XOR2_X1 U819 ( .A(n1099), .B(n1076), .Z(G30) );
NAND4_X1 U820 ( .A1(n1084), .A2(n952), .A3(n1098), .A4(n1085), .ZN(n1076) );
XNOR2_X1 U821 ( .A(G101), .B(n1071), .ZN(G3) );
NAND3_X1 U822 ( .A1(n946), .A2(n1072), .A3(n961), .ZN(n1071) );
XOR2_X1 U823 ( .A(n1002), .B(n1077), .Z(G27) );
NAND4_X1 U824 ( .A1(n945), .A2(n1085), .A3(n960), .A4(n1100), .ZN(n1077) );
NOR2_X1 U825 ( .A1(n981), .A2(n1101), .ZN(n1100) );
NAND2_X1 U826 ( .A1(n1102), .A2(n1103), .ZN(n1085) );
NAND2_X1 U827 ( .A1(n1104), .A2(n993), .ZN(n1103) );
INV_X1 U828 ( .A(G900), .ZN(n993) );
XOR2_X1 U829 ( .A(G122), .B(n1105), .Z(G24) );
NOR2_X1 U830 ( .A1(KEYINPUT62), .A2(n1070), .ZN(n1105) );
NAND4_X1 U831 ( .A1(n1092), .A2(n1106), .A3(n982), .A4(n945), .ZN(n1070) );
INV_X1 U832 ( .A(n942), .ZN(n982) );
NAND2_X1 U833 ( .A1(n1107), .A2(n1108), .ZN(n942) );
INV_X1 U834 ( .A(n1090), .ZN(n1092) );
NAND2_X1 U835 ( .A1(n1109), .A2(n973), .ZN(n1090) );
XOR2_X1 U836 ( .A(G119), .B(n1110), .Z(G21) );
NOR2_X1 U837 ( .A1(KEYINPUT61), .A2(n1069), .ZN(n1110) );
NAND3_X1 U838 ( .A1(n1106), .A2(n946), .A3(n1084), .ZN(n1069) );
AND3_X1 U839 ( .A1(n945), .A2(n1096), .A3(n1095), .ZN(n1084) );
XOR2_X1 U840 ( .A(n1111), .B(n1065), .Z(G18) );
NAND4_X1 U841 ( .A1(n961), .A2(n1106), .A3(n952), .A4(n945), .ZN(n1065) );
XOR2_X1 U842 ( .A(n1112), .B(KEYINPUT28), .Z(n945) );
NOR2_X1 U843 ( .A1(n1109), .A2(n1113), .ZN(n952) );
XNOR2_X1 U844 ( .A(G113), .B(n1066), .ZN(G15) );
NAND4_X1 U845 ( .A1(n961), .A2(n951), .A3(n1106), .A4(n1112), .ZN(n1066) );
AND2_X1 U846 ( .A1(n960), .A2(n1114), .ZN(n1106) );
NOR2_X1 U847 ( .A1(n1115), .A2(n1116), .ZN(n960) );
AND2_X1 U848 ( .A1(G221), .A2(n967), .ZN(n1116) );
INV_X1 U849 ( .A(n1101), .ZN(n951) );
NAND2_X1 U850 ( .A1(n1113), .A2(n1109), .ZN(n1101) );
AND2_X1 U851 ( .A1(n1095), .A2(n1107), .ZN(n961) );
XOR2_X1 U852 ( .A(n1108), .B(KEYINPUT60), .Z(n1095) );
XOR2_X1 U853 ( .A(G110), .B(n1073), .Z(G12) );
AND3_X1 U854 ( .A1(n946), .A2(n1072), .A3(n962), .ZN(n1073) );
INV_X1 U855 ( .A(n981), .ZN(n962) );
NAND2_X1 U856 ( .A1(n1108), .A2(n1096), .ZN(n981) );
INV_X1 U857 ( .A(n1107), .ZN(n1096) );
XNOR2_X1 U858 ( .A(n1117), .B(n1025), .ZN(n1107) );
NAND2_X1 U859 ( .A1(G217), .A2(n967), .ZN(n1025) );
OR2_X1 U860 ( .A1(n1024), .A2(n1118), .ZN(n1117) );
XNOR2_X1 U861 ( .A(n1119), .B(n1120), .ZN(n1024) );
XOR2_X1 U862 ( .A(KEYINPUT47), .B(KEYINPUT24), .Z(n1120) );
XOR2_X1 U863 ( .A(n1121), .B(n1122), .Z(n1119) );
XOR2_X1 U864 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U865 ( .A(G119), .B(G110), .Z(n1124) );
XOR2_X1 U866 ( .A(G146), .B(G137), .Z(n1123) );
XOR2_X1 U867 ( .A(n1125), .B(n1126), .Z(n1121) );
XNOR2_X1 U868 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U869 ( .A1(G128), .A2(KEYINPUT56), .ZN(n1128) );
NAND2_X1 U870 ( .A1(KEYINPUT12), .A2(n1002), .ZN(n1127) );
INV_X1 U871 ( .A(G125), .ZN(n1002) );
XOR2_X1 U872 ( .A(n1129), .B(n1130), .Z(n1125) );
NAND2_X1 U873 ( .A1(n1131), .A2(G221), .ZN(n1129) );
XOR2_X1 U874 ( .A(n1132), .B(G472), .Z(n1108) );
NAND3_X1 U875 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U876 ( .A1(KEYINPUT49), .A2(n1136), .ZN(n1134) );
NAND3_X1 U877 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NAND2_X1 U878 ( .A1(n1140), .A2(KEYINPUT8), .ZN(n1139) );
NAND3_X1 U879 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1138) );
INV_X1 U880 ( .A(KEYINPUT8), .ZN(n1142) );
OR2_X1 U881 ( .A1(n1143), .A2(n1141), .ZN(n1137) );
NOR2_X1 U882 ( .A1(n1140), .A2(KEYINPUT22), .ZN(n1141) );
NAND4_X1 U883 ( .A1(n1144), .A2(n1145), .A3(n1143), .A4(n1146), .ZN(n1133) );
INV_X1 U884 ( .A(KEYINPUT49), .ZN(n1146) );
XNOR2_X1 U885 ( .A(n1147), .B(n1051), .ZN(n1143) );
XOR2_X1 U886 ( .A(G113), .B(n1148), .Z(n1051) );
XOR2_X1 U887 ( .A(G119), .B(G116), .Z(n1148) );
XNOR2_X1 U888 ( .A(n1052), .B(KEYINPUT7), .ZN(n1147) );
XNOR2_X1 U889 ( .A(n1149), .B(n1150), .ZN(n1052) );
NAND2_X1 U890 ( .A1(KEYINPUT8), .A2(n1151), .ZN(n1145) );
OR2_X1 U891 ( .A1(n1140), .A2(KEYINPUT22), .ZN(n1151) );
OR2_X1 U892 ( .A1(n1140), .A2(KEYINPUT8), .ZN(n1144) );
XOR2_X1 U893 ( .A(n1048), .B(G101), .Z(n1140) );
NAND2_X1 U894 ( .A1(n1152), .A2(G210), .ZN(n1048) );
AND3_X1 U895 ( .A1(n1112), .A2(n1114), .A3(n1098), .ZN(n1072) );
AND2_X1 U896 ( .A1(n1115), .A2(n1153), .ZN(n1098) );
NAND2_X1 U897 ( .A1(G221), .A2(n967), .ZN(n1153) );
NAND2_X1 U898 ( .A1(G234), .A2(n1154), .ZN(n967) );
INV_X1 U899 ( .A(n966), .ZN(n1115) );
XOR2_X1 U900 ( .A(n1155), .B(G469), .Z(n966) );
NAND2_X1 U901 ( .A1(n1156), .A2(n1135), .ZN(n1155) );
XOR2_X1 U902 ( .A(KEYINPUT37), .B(n1055), .Z(n1156) );
XNOR2_X1 U903 ( .A(n1157), .B(n1158), .ZN(n1055) );
XOR2_X1 U904 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U905 ( .A(KEYINPUT14), .B(G104), .Z(n1160) );
XOR2_X1 U906 ( .A(KEYINPUT44), .B(KEYINPUT35), .Z(n1159) );
XOR2_X1 U907 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U908 ( .A(n1163), .B(n1001), .Z(n1162) );
XOR2_X1 U909 ( .A(G140), .B(n1164), .Z(n1001) );
NOR2_X1 U910 ( .A1(KEYINPUT3), .A2(n1165), .ZN(n1164) );
XOR2_X1 U911 ( .A(n1149), .B(n1166), .Z(n1161) );
AND2_X1 U912 ( .A1(n992), .A2(G227), .ZN(n1166) );
XOR2_X1 U913 ( .A(n1167), .B(n1000), .Z(n1149) );
XNOR2_X1 U914 ( .A(n1168), .B(n1169), .ZN(n1000) );
XNOR2_X1 U915 ( .A(G131), .B(KEYINPUT26), .ZN(n1168) );
NAND2_X1 U916 ( .A1(KEYINPUT43), .A2(n1170), .ZN(n1167) );
XNOR2_X1 U917 ( .A(G137), .B(n1171), .ZN(n1170) );
NAND2_X1 U918 ( .A1(KEYINPUT30), .A2(n1097), .ZN(n1171) );
INV_X1 U919 ( .A(G134), .ZN(n1097) );
NAND2_X1 U920 ( .A1(n1102), .A2(n1172), .ZN(n1114) );
NAND2_X1 U921 ( .A1(n1104), .A2(n1173), .ZN(n1172) );
INV_X1 U922 ( .A(G898), .ZN(n1173) );
NOR3_X1 U923 ( .A1(n1174), .A2(n936), .A3(n992), .ZN(n1104) );
INV_X1 U924 ( .A(n1175), .ZN(n936) );
NAND3_X1 U925 ( .A1(n1175), .A2(n992), .A3(n1176), .ZN(n1102) );
XNOR2_X1 U926 ( .A(G952), .B(KEYINPUT19), .ZN(n1176) );
NAND2_X1 U927 ( .A1(G234), .A2(n1177), .ZN(n1175) );
XOR2_X1 U928 ( .A(KEYINPUT41), .B(G237), .Z(n1177) );
NOR2_X1 U929 ( .A1(n956), .A2(n950), .ZN(n1112) );
INV_X1 U930 ( .A(n953), .ZN(n950) );
NAND2_X1 U931 ( .A1(G214), .A2(n1178), .ZN(n953) );
INV_X1 U932 ( .A(n1062), .ZN(n1178) );
XOR2_X1 U933 ( .A(n1179), .B(n1180), .Z(n956) );
NOR2_X1 U934 ( .A1(n1062), .A2(n1063), .ZN(n1180) );
INV_X1 U935 ( .A(G210), .ZN(n1063) );
NOR2_X1 U936 ( .A1(n1181), .A2(G237), .ZN(n1062) );
INV_X1 U937 ( .A(n1154), .ZN(n1181) );
XOR2_X1 U938 ( .A(n1174), .B(KEYINPUT52), .Z(n1154) );
INV_X1 U939 ( .A(G902), .ZN(n1174) );
NAND2_X1 U940 ( .A1(n1182), .A2(n1135), .ZN(n1179) );
XOR2_X1 U941 ( .A(n1019), .B(n1183), .Z(n1182) );
NOR2_X1 U942 ( .A1(KEYINPUT45), .A2(n1083), .ZN(n1183) );
XOR2_X1 U943 ( .A(n1184), .B(n1185), .Z(n1083) );
XOR2_X1 U944 ( .A(G125), .B(n1150), .Z(n1185) );
NOR2_X1 U945 ( .A1(KEYINPUT25), .A2(n1165), .ZN(n1150) );
XOR2_X1 U946 ( .A(G143), .B(KEYINPUT40), .Z(n1165) );
XOR2_X1 U947 ( .A(n1186), .B(n1169), .Z(n1184) );
XOR2_X1 U948 ( .A(G128), .B(G146), .Z(n1169) );
NAND2_X1 U949 ( .A1(G224), .A2(n992), .ZN(n1186) );
XNOR2_X1 U950 ( .A(n1163), .B(n1187), .ZN(n1019) );
XOR2_X1 U951 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U952 ( .A1(KEYINPUT55), .A2(n1190), .ZN(n1188) );
XOR2_X1 U953 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U954 ( .A(KEYINPUT39), .B(G116), .Z(n1192) );
NOR2_X1 U955 ( .A1(G119), .A2(KEYINPUT11), .ZN(n1191) );
XOR2_X1 U956 ( .A(G101), .B(n1193), .Z(n1163) );
XOR2_X1 U957 ( .A(G110), .B(G107), .Z(n1193) );
NOR2_X1 U958 ( .A1(n973), .A2(n1109), .ZN(n946) );
XOR2_X1 U959 ( .A(n979), .B(n1194), .Z(n1109) );
NOR2_X1 U960 ( .A1(KEYINPUT58), .A2(n978), .ZN(n1194) );
INV_X1 U961 ( .A(G475), .ZN(n978) );
NOR2_X1 U962 ( .A1(n1033), .A2(n1118), .ZN(n979) );
XNOR2_X1 U963 ( .A(n1195), .B(n1196), .ZN(n1033) );
XOR2_X1 U964 ( .A(n1189), .B(n1197), .Z(n1196) );
XOR2_X1 U965 ( .A(n1198), .B(n1130), .Z(n1197) );
XOR2_X1 U966 ( .A(G140), .B(KEYINPUT36), .Z(n1130) );
NAND2_X1 U967 ( .A1(n1199), .A2(KEYINPUT2), .ZN(n1198) );
XOR2_X1 U968 ( .A(n1200), .B(G143), .Z(n1199) );
NAND2_X1 U969 ( .A1(n1152), .A2(G214), .ZN(n1200) );
NOR2_X1 U970 ( .A1(G953), .A2(G237), .ZN(n1152) );
XOR2_X1 U971 ( .A(n1035), .B(n1201), .Z(n1189) );
XOR2_X1 U972 ( .A(G122), .B(G113), .Z(n1201) );
INV_X1 U973 ( .A(G104), .ZN(n1035) );
XOR2_X1 U974 ( .A(n1202), .B(n1203), .Z(n1195) );
XOR2_X1 U975 ( .A(G125), .B(n1204), .Z(n1203) );
NOR2_X1 U976 ( .A1(G146), .A2(KEYINPUT46), .ZN(n1204) );
XNOR2_X1 U977 ( .A(G131), .B(KEYINPUT9), .ZN(n1202) );
INV_X1 U978 ( .A(n1113), .ZN(n973) );
XOR2_X1 U979 ( .A(n1205), .B(G478), .Z(n1113) );
OR2_X1 U980 ( .A1(n1029), .A2(n1118), .ZN(n1205) );
INV_X1 U981 ( .A(n1135), .ZN(n1118) );
XOR2_X1 U982 ( .A(G902), .B(KEYINPUT59), .Z(n1135) );
XNOR2_X1 U983 ( .A(n1206), .B(n1207), .ZN(n1029) );
XOR2_X1 U984 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U985 ( .A(n1210), .B(n1211), .ZN(n1209) );
NAND2_X1 U986 ( .A1(KEYINPUT16), .A2(G122), .ZN(n1211) );
NAND2_X1 U987 ( .A1(KEYINPUT51), .A2(n930), .ZN(n1210) );
INV_X1 U988 ( .A(G107), .ZN(n930) );
NAND2_X1 U989 ( .A1(G217), .A2(n1131), .ZN(n1208) );
AND2_X1 U990 ( .A1(G234), .A2(n992), .ZN(n1131) );
INV_X1 U991 ( .A(G953), .ZN(n992) );
XOR2_X1 U992 ( .A(n1212), .B(n1213), .Z(n1206) );
NOR2_X1 U993 ( .A1(KEYINPUT42), .A2(n1214), .ZN(n1213) );
XOR2_X1 U994 ( .A(n1099), .B(n1215), .Z(n1214) );
XOR2_X1 U995 ( .A(G143), .B(G134), .Z(n1215) );
INV_X1 U996 ( .A(G128), .ZN(n1099) );
XOR2_X1 U997 ( .A(n1111), .B(KEYINPUT57), .Z(n1212) );
INV_X1 U998 ( .A(G116), .ZN(n1111) );
endmodule


