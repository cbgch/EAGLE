//Key = 1010100111010011010101010101100010011100010110101000111000110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313;

XOR2_X1 U720 ( .A(G107), .B(n1003), .Z(G9) );
NOR2_X1 U721 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR4_X1 U722 ( .A1(G953), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1005) );
NOR2_X1 U723 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U724 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U725 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U728 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR3_X1 U729 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR2_X1 U730 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XNOR2_X1 U731 ( .A(n1026), .B(KEYINPUT4), .ZN(n1025) );
NOR3_X1 U732 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1022) );
NOR4_X1 U733 ( .A1(n1030), .A2(n1027), .A3(n1031), .A4(n1032), .ZN(n1019) );
INV_X1 U734 ( .A(n1033), .ZN(n1031) );
NOR3_X1 U735 ( .A1(n1034), .A2(n1030), .A3(n1027), .ZN(n1015) );
AND4_X1 U736 ( .A1(n1026), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1030) );
NAND2_X1 U737 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U738 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
OR2_X1 U739 ( .A1(n1042), .A2(KEYINPUT38), .ZN(n1041) );
NAND2_X1 U740 ( .A1(n1033), .A2(n1032), .ZN(n1040) );
INV_X1 U741 ( .A(KEYINPUT63), .ZN(n1032) );
INV_X1 U742 ( .A(n1018), .ZN(n1038) );
NAND3_X1 U743 ( .A1(KEYINPUT38), .A2(n1043), .A3(n1018), .ZN(n1036) );
NAND2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR4_X1 U747 ( .A1(n1021), .A2(n1050), .A3(n1034), .A4(n1018), .ZN(n1011) );
INV_X1 U748 ( .A(n1026), .ZN(n1034) );
INV_X1 U749 ( .A(n1044), .ZN(n1021) );
NOR3_X1 U750 ( .A1(n1006), .A2(G953), .A3(G952), .ZN(n1004) );
AND4_X1 U751 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1006) );
NOR4_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
XNOR2_X1 U753 ( .A(n1059), .B(n1060), .ZN(n1058) );
XNOR2_X1 U754 ( .A(n1061), .B(KEYINPUT15), .ZN(n1055) );
NOR3_X1 U755 ( .A1(n1062), .A2(n1027), .A3(n1048), .ZN(n1053) );
INV_X1 U756 ( .A(n1063), .ZN(n1048) );
AND2_X1 U757 ( .A1(n1064), .A2(G472), .ZN(n1062) );
XOR2_X1 U758 ( .A(KEYINPUT14), .B(n1065), .Z(n1052) );
NOR2_X1 U759 ( .A1(G472), .A2(n1064), .ZN(n1065) );
XOR2_X1 U760 ( .A(KEYINPUT33), .B(n1066), .Z(n1051) );
NOR2_X1 U761 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(G72) );
NAND2_X1 U764 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U765 ( .A(n1075), .B(n1076), .Z(n1073) );
NAND2_X1 U766 ( .A1(KEYINPUT2), .A2(n1077), .ZN(n1076) );
NAND2_X1 U767 ( .A1(n1078), .A2(G953), .ZN(n1071) );
XOR2_X1 U768 ( .A(n1075), .B(n1079), .Z(n1078) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U770 ( .A1(n1082), .A2(n1083), .ZN(n1075) );
NAND2_X1 U771 ( .A1(G953), .A2(n1081), .ZN(n1083) );
XOR2_X1 U772 ( .A(n1084), .B(n1085), .Z(n1082) );
XNOR2_X1 U773 ( .A(n1086), .B(n1087), .ZN(n1085) );
XNOR2_X1 U774 ( .A(n1088), .B(n1089), .ZN(n1087) );
NOR2_X1 U775 ( .A1(G134), .A2(KEYINPUT61), .ZN(n1089) );
NAND2_X1 U776 ( .A1(KEYINPUT23), .A2(G125), .ZN(n1088) );
XNOR2_X1 U777 ( .A(n1090), .B(n1091), .ZN(n1084) );
XNOR2_X1 U778 ( .A(n1092), .B(G137), .ZN(n1091) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(G69) );
XOR2_X1 U780 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U782 ( .A(n1099), .B(n1100), .ZN(n1098) );
NOR2_X1 U783 ( .A1(G898), .A2(n1074), .ZN(n1097) );
NOR2_X1 U784 ( .A1(n1101), .A2(G953), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U786 ( .A1(n1104), .A2(n1074), .ZN(n1093) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U790 ( .A1(n1111), .A2(n1070), .ZN(n1109) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1112), .ZN(G63) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U793 ( .A1(n1111), .A2(G478), .ZN(n1113) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1115), .ZN(G60) );
XOR2_X1 U795 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U796 ( .A1(n1111), .A2(G475), .ZN(n1116) );
XOR2_X1 U797 ( .A(G104), .B(n1102), .Z(G6) );
NOR2_X1 U798 ( .A1(n1107), .A2(n1118), .ZN(G57) );
XOR2_X1 U799 ( .A(n1119), .B(n1120), .Z(n1118) );
XNOR2_X1 U800 ( .A(n1121), .B(n1122), .ZN(n1120) );
NAND3_X1 U801 ( .A1(n1111), .A2(G472), .A3(KEYINPUT52), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1119) );
XOR2_X1 U803 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U804 ( .A1(KEYINPUT49), .A2(n1127), .ZN(n1126) );
NAND2_X1 U805 ( .A1(KEYINPUT7), .A2(n1086), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(G54) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1132) );
NOR2_X1 U810 ( .A1(KEYINPUT29), .A2(n1086), .ZN(n1135) );
NAND2_X1 U811 ( .A1(n1111), .A2(G469), .ZN(n1134) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1130) );
XNOR2_X1 U813 ( .A(KEYINPUT31), .B(n1092), .ZN(n1137) );
XNOR2_X1 U814 ( .A(n1138), .B(n1139), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1140), .A2(KEYINPUT55), .ZN(n1139) );
NOR2_X1 U816 ( .A1(KEYINPUT39), .A2(n1141), .ZN(n1138) );
XNOR2_X1 U817 ( .A(n1107), .B(KEYINPUT59), .ZN(n1128) );
NOR2_X1 U818 ( .A1(n1107), .A2(n1142), .ZN(G51) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U820 ( .A(n1145), .B(n1146), .ZN(n1144) );
XOR2_X1 U821 ( .A(n1147), .B(n1148), .Z(n1143) );
NOR2_X1 U822 ( .A1(KEYINPUT62), .A2(n1149), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1147) );
NAND3_X1 U824 ( .A1(n1111), .A2(n1152), .A3(n1153), .ZN(n1150) );
XNOR2_X1 U825 ( .A(G210), .B(KEYINPUT35), .ZN(n1153) );
AND2_X1 U826 ( .A1(G902), .A2(n1008), .ZN(n1111) );
OR3_X1 U827 ( .A1(n1077), .A2(n1103), .A3(n1154), .ZN(n1008) );
XOR2_X1 U828 ( .A(n1102), .B(KEYINPUT20), .Z(n1154) );
AND3_X1 U829 ( .A1(n1155), .A2(n1026), .A3(n1043), .ZN(n1102) );
NAND4_X1 U830 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1103) );
NOR4_X1 U831 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1003), .ZN(n1159) );
AND3_X1 U832 ( .A1(n1033), .A2(n1026), .A3(n1155), .ZN(n1003) );
INV_X1 U833 ( .A(n1163), .ZN(n1160) );
NAND4_X1 U834 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1077) );
NOR4_X1 U835 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
INV_X1 U836 ( .A(n1172), .ZN(n1168) );
NOR2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1050), .A2(n1175), .ZN(n1174) );
NOR3_X1 U839 ( .A1(n1176), .A2(n1177), .A3(n1042), .ZN(n1173) );
XOR2_X1 U840 ( .A(KEYINPUT53), .B(n1028), .Z(n1176) );
NOR2_X1 U841 ( .A1(n1074), .A2(G952), .ZN(n1107) );
XNOR2_X1 U842 ( .A(G146), .B(n1164), .ZN(G48) );
NAND3_X1 U843 ( .A1(n1178), .A2(n1179), .A3(n1043), .ZN(n1164) );
XNOR2_X1 U844 ( .A(G143), .B(n1165), .ZN(G45) );
NAND4_X1 U845 ( .A1(n1029), .A2(n1178), .A3(n1061), .A4(n1056), .ZN(n1165) );
XNOR2_X1 U846 ( .A(n1092), .B(n1180), .ZN(G42) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1181), .ZN(n1180) );
INV_X1 U848 ( .A(n1182), .ZN(n1177) );
XNOR2_X1 U849 ( .A(n1171), .B(n1183), .ZN(G39) );
NAND2_X1 U850 ( .A1(KEYINPUT8), .A2(G137), .ZN(n1183) );
AND3_X1 U851 ( .A1(n1179), .A2(n1044), .A3(n1182), .ZN(n1171) );
XNOR2_X1 U852 ( .A(n1184), .B(n1170), .ZN(G36) );
AND3_X1 U853 ( .A1(n1182), .A2(n1033), .A3(n1029), .ZN(n1170) );
XNOR2_X1 U854 ( .A(n1090), .B(n1169), .ZN(G33) );
AND3_X1 U855 ( .A1(n1043), .A2(n1182), .A3(n1029), .ZN(n1169) );
NOR4_X1 U856 ( .A1(n1185), .A2(n1046), .A3(n1014), .A4(n1027), .ZN(n1182) );
INV_X1 U857 ( .A(n1024), .ZN(n1027) );
XNOR2_X1 U858 ( .A(G128), .B(n1172), .ZN(G30) );
NAND3_X1 U859 ( .A1(n1179), .A2(n1033), .A3(n1178), .ZN(n1172) );
NOR3_X1 U860 ( .A1(n1046), .A2(n1050), .A3(n1185), .ZN(n1178) );
XOR2_X1 U861 ( .A(G101), .B(n1162), .Z(G3) );
AND3_X1 U862 ( .A1(n1155), .A2(n1044), .A3(n1029), .ZN(n1162) );
XOR2_X1 U863 ( .A(n1186), .B(n1187), .Z(G27) );
XNOR2_X1 U864 ( .A(KEYINPUT3), .B(n1149), .ZN(n1187) );
NOR2_X1 U865 ( .A1(n1188), .A2(n1050), .ZN(n1186) );
XOR2_X1 U866 ( .A(n1175), .B(KEYINPUT6), .Z(n1188) );
OR3_X1 U867 ( .A1(n1181), .A2(n1185), .A3(n1018), .ZN(n1175) );
NAND2_X1 U868 ( .A1(n1189), .A2(n1190), .ZN(n1185) );
NAND2_X1 U869 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND3_X1 U870 ( .A1(G902), .A2(n1081), .A3(G953), .ZN(n1191) );
INV_X1 U871 ( .A(G900), .ZN(n1081) );
NAND2_X1 U872 ( .A1(n1028), .A2(n1043), .ZN(n1181) );
XNOR2_X1 U873 ( .A(G122), .B(n1158), .ZN(G24) );
NAND4_X1 U874 ( .A1(n1193), .A2(n1026), .A3(n1061), .A4(n1056), .ZN(n1158) );
NOR2_X1 U875 ( .A1(n1194), .A2(n1195), .ZN(n1026) );
XNOR2_X1 U876 ( .A(G119), .B(n1156), .ZN(G21) );
NAND3_X1 U877 ( .A1(n1179), .A2(n1044), .A3(n1193), .ZN(n1156) );
NOR2_X1 U878 ( .A1(n1196), .A2(n1197), .ZN(n1179) );
XOR2_X1 U879 ( .A(G116), .B(n1161), .Z(G18) );
AND3_X1 U880 ( .A1(n1029), .A2(n1033), .A3(n1193), .ZN(n1161) );
XNOR2_X1 U881 ( .A(G113), .B(n1157), .ZN(G15) );
NAND3_X1 U882 ( .A1(n1029), .A2(n1043), .A3(n1193), .ZN(n1157) );
NOR2_X1 U883 ( .A1(n1018), .A2(n1198), .ZN(n1193) );
NAND2_X1 U884 ( .A1(n1049), .A2(n1199), .ZN(n1018) );
XNOR2_X1 U885 ( .A(KEYINPUT17), .B(n1063), .ZN(n1199) );
INV_X1 U886 ( .A(n1057), .ZN(n1049) );
INV_X1 U887 ( .A(n1042), .ZN(n1043) );
NAND2_X1 U888 ( .A1(n1200), .A2(n1056), .ZN(n1042) );
XNOR2_X1 U889 ( .A(n1061), .B(KEYINPUT5), .ZN(n1200) );
NOR2_X1 U890 ( .A1(n1196), .A2(n1194), .ZN(n1029) );
XNOR2_X1 U891 ( .A(G110), .B(n1163), .ZN(G12) );
NAND3_X1 U892 ( .A1(n1155), .A2(n1044), .A3(n1028), .ZN(n1163) );
NOR2_X1 U893 ( .A1(n1195), .A2(n1197), .ZN(n1028) );
INV_X1 U894 ( .A(n1194), .ZN(n1197) );
NAND3_X1 U895 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1194) );
INV_X1 U896 ( .A(n1068), .ZN(n1203) );
NOR2_X1 U897 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
OR2_X1 U898 ( .A1(n1070), .A2(KEYINPUT0), .ZN(n1202) );
NAND3_X1 U899 ( .A1(n1070), .A2(n1069), .A3(KEYINPUT0), .ZN(n1201) );
NAND2_X1 U900 ( .A1(n1110), .A2(n1204), .ZN(n1069) );
XNOR2_X1 U901 ( .A(n1205), .B(n1206), .ZN(n1110) );
XOR2_X1 U902 ( .A(G137), .B(n1207), .Z(n1206) );
AND3_X1 U903 ( .A1(G221), .A2(n1074), .A3(G234), .ZN(n1207) );
NAND4_X1 U904 ( .A1(KEYINPUT44), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1205) );
NAND3_X1 U905 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
INV_X1 U906 ( .A(KEYINPUT22), .ZN(n1212) );
OR2_X1 U907 ( .A1(n1213), .A2(n1211), .ZN(n1209) );
NOR2_X1 U908 ( .A1(KEYINPUT57), .A2(n1214), .ZN(n1211) );
XOR2_X1 U909 ( .A(n1215), .B(n1216), .Z(n1213) );
XNOR2_X1 U910 ( .A(KEYINPUT27), .B(n1217), .ZN(n1216) );
INV_X1 U911 ( .A(G146), .ZN(n1217) );
XNOR2_X1 U912 ( .A(n1218), .B(n1149), .ZN(n1215) );
NAND2_X1 U913 ( .A1(KEYINPUT9), .A2(G140), .ZN(n1218) );
NAND2_X1 U914 ( .A1(KEYINPUT22), .A2(n1214), .ZN(n1208) );
XNOR2_X1 U915 ( .A(n1141), .B(n1219), .ZN(n1214) );
NOR2_X1 U916 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XOR2_X1 U917 ( .A(n1222), .B(KEYINPUT58), .Z(n1221) );
NAND2_X1 U918 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U919 ( .A(KEYINPUT30), .B(G119), .Z(n1223) );
NOR2_X1 U920 ( .A1(G119), .A2(n1224), .ZN(n1220) );
INV_X1 U921 ( .A(G128), .ZN(n1224) );
AND2_X1 U922 ( .A1(G217), .A2(n1225), .ZN(n1070) );
INV_X1 U923 ( .A(n1196), .ZN(n1195) );
XNOR2_X1 U924 ( .A(n1064), .B(n1226), .ZN(n1196) );
XOR2_X1 U925 ( .A(KEYINPUT54), .B(G472), .Z(n1226) );
NAND2_X1 U926 ( .A1(n1227), .A2(n1204), .ZN(n1064) );
XNOR2_X1 U927 ( .A(n1228), .B(n1127), .ZN(n1227) );
NAND2_X1 U928 ( .A1(n1229), .A2(G210), .ZN(n1127) );
XOR2_X1 U929 ( .A(n1230), .B(G101), .Z(n1228) );
NAND2_X1 U930 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U931 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U932 ( .A1(KEYINPUT48), .A2(n1235), .ZN(n1234) );
OR2_X1 U933 ( .A1(n1125), .A2(KEYINPUT13), .ZN(n1235) );
NAND2_X1 U934 ( .A1(n1236), .A2(n1125), .ZN(n1231) );
NAND2_X1 U935 ( .A1(n1237), .A2(n1238), .ZN(n1125) );
NAND2_X1 U936 ( .A1(G113), .A2(n1239), .ZN(n1238) );
XOR2_X1 U937 ( .A(KEYINPUT11), .B(n1240), .Z(n1237) );
NOR2_X1 U938 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U939 ( .A(KEYINPUT42), .B(n1239), .Z(n1242) );
XNOR2_X1 U940 ( .A(G113), .B(KEYINPUT36), .ZN(n1241) );
NAND2_X1 U941 ( .A1(n1243), .A2(n1244), .ZN(n1236) );
NAND2_X1 U942 ( .A1(KEYINPUT48), .A2(n1245), .ZN(n1244) );
INV_X1 U943 ( .A(n1233), .ZN(n1245) );
XOR2_X1 U944 ( .A(n1246), .B(n1086), .Z(n1233) );
INV_X1 U945 ( .A(KEYINPUT13), .ZN(n1243) );
NAND2_X1 U946 ( .A1(n1247), .A2(n1248), .ZN(n1044) );
OR3_X1 U947 ( .A1(n1056), .A2(n1061), .A3(KEYINPUT5), .ZN(n1248) );
NAND2_X1 U948 ( .A1(KEYINPUT5), .A2(n1033), .ZN(n1247) );
NOR2_X1 U949 ( .A1(n1056), .A2(n1249), .ZN(n1033) );
INV_X1 U950 ( .A(n1061), .ZN(n1249) );
XNOR2_X1 U951 ( .A(n1250), .B(G478), .ZN(n1061) );
NAND2_X1 U952 ( .A1(n1114), .A2(n1204), .ZN(n1250) );
XNOR2_X1 U953 ( .A(n1251), .B(n1252), .ZN(n1114) );
NOR2_X1 U954 ( .A1(KEYINPUT40), .A2(n1253), .ZN(n1252) );
XOR2_X1 U955 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U956 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U957 ( .A1(KEYINPUT43), .A2(n1258), .ZN(n1256) );
XOR2_X1 U958 ( .A(G122), .B(G116), .Z(n1258) );
XNOR2_X1 U959 ( .A(G107), .B(n1259), .ZN(n1254) );
XNOR2_X1 U960 ( .A(n1184), .B(G128), .ZN(n1259) );
INV_X1 U961 ( .A(G134), .ZN(n1184) );
NAND3_X1 U962 ( .A1(G234), .A2(n1074), .A3(G217), .ZN(n1251) );
XNOR2_X1 U963 ( .A(n1260), .B(G475), .ZN(n1056) );
NAND2_X1 U964 ( .A1(n1117), .A2(n1204), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1261), .B(n1262), .ZN(n1117) );
XNOR2_X1 U966 ( .A(n1263), .B(G104), .ZN(n1262) );
XOR2_X1 U967 ( .A(n1264), .B(n1265), .Z(n1261) );
XOR2_X1 U968 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U969 ( .A(n1090), .B(G125), .ZN(n1267) );
INV_X1 U970 ( .A(G131), .ZN(n1090) );
XOR2_X1 U971 ( .A(KEYINPUT47), .B(KEYINPUT28), .Z(n1266) );
XOR2_X1 U972 ( .A(n1268), .B(n1269), .Z(n1264) );
XOR2_X1 U973 ( .A(G122), .B(n1270), .Z(n1269) );
NOR2_X1 U974 ( .A1(G140), .A2(KEYINPUT50), .ZN(n1270) );
XNOR2_X1 U975 ( .A(n1271), .B(n1272), .ZN(n1268) );
AND2_X1 U976 ( .A1(G214), .A2(n1229), .ZN(n1272) );
NOR2_X1 U977 ( .A1(G953), .A2(G237), .ZN(n1229) );
NOR2_X1 U978 ( .A1(n1198), .A2(n1046), .ZN(n1155) );
NAND2_X1 U979 ( .A1(n1057), .A2(n1063), .ZN(n1046) );
NAND2_X1 U980 ( .A1(G221), .A2(n1225), .ZN(n1063) );
NAND2_X1 U981 ( .A1(n1273), .A2(G234), .ZN(n1225) );
XNOR2_X1 U982 ( .A(n1274), .B(G469), .ZN(n1057) );
NAND2_X1 U983 ( .A1(n1275), .A2(n1204), .ZN(n1274) );
XOR2_X1 U984 ( .A(n1276), .B(n1133), .Z(n1275) );
XNOR2_X1 U985 ( .A(n1277), .B(n1122), .ZN(n1133) );
XOR2_X1 U986 ( .A(G101), .B(n1246), .Z(n1122) );
XOR2_X1 U987 ( .A(G131), .B(n1278), .Z(n1246) );
NOR2_X1 U988 ( .A1(KEYINPUT10), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U989 ( .A(G134), .B(G137), .ZN(n1279) );
NAND2_X1 U990 ( .A1(KEYINPUT21), .A2(n1280), .ZN(n1277) );
XNOR2_X1 U991 ( .A(n1281), .B(n1086), .ZN(n1276) );
INV_X1 U992 ( .A(n1145), .ZN(n1086) );
NAND2_X1 U993 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND3_X1 U994 ( .A1(n1092), .A2(n1284), .A3(n1285), .ZN(n1283) );
XOR2_X1 U995 ( .A(n1140), .B(n1286), .Z(n1285) );
NOR2_X1 U996 ( .A1(n1141), .A2(n1287), .ZN(n1286) );
INV_X1 U997 ( .A(G110), .ZN(n1141) );
NAND2_X1 U998 ( .A1(n1288), .A2(n1289), .ZN(n1282) );
NAND2_X1 U999 ( .A1(n1092), .A2(n1284), .ZN(n1289) );
INV_X1 U1000 ( .A(KEYINPUT26), .ZN(n1284) );
INV_X1 U1001 ( .A(G140), .ZN(n1092) );
XOR2_X1 U1002 ( .A(n1140), .B(n1290), .Z(n1288) );
NOR2_X1 U1003 ( .A1(G110), .A2(n1287), .ZN(n1290) );
INV_X1 U1004 ( .A(KEYINPUT41), .ZN(n1287) );
NOR2_X1 U1005 ( .A1(n1080), .A2(G953), .ZN(n1140) );
INV_X1 U1006 ( .A(G227), .ZN(n1080) );
OR3_X1 U1007 ( .A1(n1291), .A2(n1009), .A3(n1050), .ZN(n1198) );
NAND2_X1 U1008 ( .A1(n1014), .A2(n1024), .ZN(n1050) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1152), .ZN(n1024) );
INV_X1 U1010 ( .A(n1292), .ZN(n1152) );
XOR2_X1 U1011 ( .A(n1059), .B(n1293), .Z(n1014) );
NOR2_X1 U1012 ( .A1(n1060), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U1013 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n1294) );
NOR2_X1 U1014 ( .A1(n1292), .A2(n1295), .ZN(n1060) );
INV_X1 U1015 ( .A(G210), .ZN(n1295) );
NOR2_X1 U1016 ( .A1(n1296), .A2(G237), .ZN(n1292) );
INV_X1 U1017 ( .A(n1273), .ZN(n1296) );
XNOR2_X1 U1018 ( .A(G902), .B(KEYINPUT34), .ZN(n1273) );
NAND2_X1 U1019 ( .A1(n1297), .A2(n1204), .ZN(n1059) );
INV_X1 U1020 ( .A(G902), .ZN(n1204) );
XOR2_X1 U1021 ( .A(n1298), .B(n1146), .Z(n1297) );
XNOR2_X1 U1022 ( .A(n1299), .B(n1100), .ZN(n1146) );
XNOR2_X1 U1023 ( .A(n1300), .B(n1301), .ZN(n1100) );
XNOR2_X1 U1024 ( .A(n1302), .B(n1303), .ZN(n1301) );
NOR2_X1 U1025 ( .A1(G122), .A2(KEYINPUT56), .ZN(n1303) );
NAND2_X1 U1026 ( .A1(KEYINPUT32), .A2(n1239), .ZN(n1302) );
XOR2_X1 U1027 ( .A(G116), .B(G119), .Z(n1239) );
XNOR2_X1 U1028 ( .A(G110), .B(n1304), .ZN(n1300) );
XNOR2_X1 U1029 ( .A(KEYINPUT25), .B(n1263), .ZN(n1304) );
INV_X1 U1030 ( .A(G113), .ZN(n1263) );
NAND2_X1 U1031 ( .A1(KEYINPUT46), .A2(n1099), .ZN(n1299) );
XNOR2_X1 U1032 ( .A(n1305), .B(n1306), .ZN(n1099) );
XOR2_X1 U1033 ( .A(n1307), .B(n1280), .Z(n1306) );
XOR2_X1 U1034 ( .A(G104), .B(G107), .Z(n1280) );
NOR2_X1 U1035 ( .A1(G101), .A2(KEYINPUT45), .ZN(n1307) );
XNOR2_X1 U1036 ( .A(KEYINPUT24), .B(KEYINPUT16), .ZN(n1305) );
NOR2_X1 U1037 ( .A1(KEYINPUT60), .A2(n1308), .ZN(n1298) );
XOR2_X1 U1038 ( .A(n1309), .B(n1310), .Z(n1308) );
XNOR2_X1 U1039 ( .A(n1149), .B(n1151), .ZN(n1310) );
NOR2_X1 U1040 ( .A1(n1105), .A2(G953), .ZN(n1151) );
INV_X1 U1041 ( .A(G224), .ZN(n1105) );
INV_X1 U1042 ( .A(G125), .ZN(n1149) );
NAND2_X1 U1043 ( .A1(n1311), .A2(KEYINPUT37), .ZN(n1309) );
XNOR2_X1 U1044 ( .A(n1145), .B(KEYINPUT1), .ZN(n1311) );
XOR2_X1 U1045 ( .A(G128), .B(n1271), .Z(n1145) );
XNOR2_X1 U1046 ( .A(G146), .B(n1257), .ZN(n1271) );
XNOR2_X1 U1047 ( .A(G143), .B(KEYINPUT51), .ZN(n1257) );
INV_X1 U1048 ( .A(n1189), .ZN(n1009) );
NAND2_X1 U1049 ( .A1(G237), .A2(G234), .ZN(n1189) );
AND2_X1 U1050 ( .A1(n1192), .A2(n1312), .ZN(n1291) );
NAND3_X1 U1051 ( .A1(G902), .A2(n1106), .A3(G953), .ZN(n1312) );
INV_X1 U1052 ( .A(G898), .ZN(n1106) );
NAND2_X1 U1053 ( .A1(n1313), .A2(n1074), .ZN(n1192) );
INV_X1 U1054 ( .A(G953), .ZN(n1074) );
XOR2_X1 U1055 ( .A(KEYINPUT12), .B(G952), .Z(n1313) );
endmodule


