//Key = 0000011000110000011010100000000110110101000001111101001111110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429;

XNOR2_X1 U781 ( .A(n1083), .B(n1084), .ZN(G9) );
NAND2_X1 U782 ( .A1(KEYINPUT11), .A2(n1085), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(G75) );
NOR4_X1 U784 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1087) );
NOR4_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1090) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
NOR2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR3_X1 U788 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
NOR3_X1 U789 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1100) );
XNOR2_X1 U791 ( .A(n1108), .B(n1109), .ZN(n1106) );
NOR3_X1 U792 ( .A1(n1107), .A2(n1110), .A3(n1104), .ZN(n1096) );
NOR2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U794 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1088) );
NAND4_X1 U795 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1104), .ZN(n1118) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U798 ( .A(n1123), .B(KEYINPUT6), .ZN(n1122) );
INV_X1 U799 ( .A(n1095), .ZN(n1116) );
NOR3_X1 U800 ( .A1(n1124), .A2(G953), .A3(n1125), .ZN(n1086) );
INV_X1 U801 ( .A(n1113), .ZN(n1125) );
NAND4_X1 U802 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1113) );
NOR4_X1 U803 ( .A1(n1130), .A2(n1131), .A3(n1104), .A4(n1132), .ZN(n1129) );
INV_X1 U804 ( .A(n1133), .ZN(n1104) );
XOR2_X1 U805 ( .A(KEYINPUT30), .B(n1134), .Z(n1131) );
NOR2_X1 U806 ( .A1(G472), .A2(n1135), .ZN(n1134) );
NAND3_X1 U807 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1130) );
XOR2_X1 U808 ( .A(n1139), .B(KEYINPUT36), .Z(n1138) );
NAND2_X1 U809 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
XNOR2_X1 U810 ( .A(KEYINPUT3), .B(n1142), .ZN(n1140) );
NAND2_X1 U811 ( .A1(n1143), .A2(G478), .ZN(n1136) );
XNOR2_X1 U812 ( .A(n1144), .B(KEYINPUT60), .ZN(n1143) );
AND3_X1 U813 ( .A1(n1145), .A2(n1146), .A3(n1103), .ZN(n1128) );
NAND2_X1 U814 ( .A1(n1147), .A2(n1148), .ZN(n1127) );
NAND2_X1 U815 ( .A1(G472), .A2(n1135), .ZN(n1126) );
XNOR2_X1 U816 ( .A(KEYINPUT28), .B(n1091), .ZN(n1124) );
INV_X1 U817 ( .A(G952), .ZN(n1091) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(G72) );
NOR2_X1 U819 ( .A1(n1151), .A2(n1114), .ZN(n1150) );
AND2_X1 U820 ( .A1(G227), .A2(G900), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NAND2_X1 U822 ( .A1(n1154), .A2(n1114), .ZN(n1153) );
XNOR2_X1 U823 ( .A(n1155), .B(n1156), .ZN(n1154) );
NAND3_X1 U824 ( .A1(G900), .A2(n1155), .A3(G953), .ZN(n1152) );
XNOR2_X1 U825 ( .A(n1157), .B(n1158), .ZN(n1155) );
XOR2_X1 U826 ( .A(KEYINPUT5), .B(n1159), .Z(n1158) );
XOR2_X1 U827 ( .A(n1160), .B(n1161), .Z(n1157) );
NAND4_X1 U828 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1160) );
NAND3_X1 U829 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
NAND3_X1 U830 ( .A1(G131), .A2(n1167), .A3(G137), .ZN(n1164) );
XOR2_X1 U831 ( .A(n1169), .B(n1170), .Z(G69) );
XOR2_X1 U832 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U833 ( .A1(G953), .A2(n1173), .ZN(n1172) );
NAND2_X1 U834 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
NAND2_X1 U835 ( .A1(G224), .A2(G898), .ZN(n1175) );
XNOR2_X1 U836 ( .A(G953), .B(KEYINPUT59), .ZN(n1174) );
NAND2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(n1169) );
OR2_X1 U838 ( .A1(n1114), .A2(G898), .ZN(n1177) );
XOR2_X1 U839 ( .A(n1178), .B(n1179), .Z(n1176) );
NOR2_X1 U840 ( .A1(n1180), .A2(n1181), .ZN(G66) );
XNOR2_X1 U841 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U843 ( .A1(n1180), .A2(n1186), .ZN(G63) );
NOR3_X1 U844 ( .A1(n1144), .A2(n1187), .A3(n1188), .ZN(n1186) );
AND4_X1 U845 ( .A1(n1189), .A2(KEYINPUT22), .A3(G478), .A4(n1190), .ZN(n1188) );
NOR2_X1 U846 ( .A1(n1191), .A2(n1189), .ZN(n1187) );
AND3_X1 U847 ( .A1(KEYINPUT22), .A2(n1089), .A3(G478), .ZN(n1191) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1192), .ZN(G60) );
XOR2_X1 U849 ( .A(n1193), .B(n1194), .Z(n1192) );
AND2_X1 U850 ( .A1(G475), .A2(n1190), .ZN(n1193) );
XNOR2_X1 U851 ( .A(G104), .B(n1195), .ZN(G6) );
NAND2_X1 U852 ( .A1(n1112), .A2(n1196), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1180), .A2(n1197), .ZN(G57) );
XNOR2_X1 U854 ( .A(n1198), .B(n1199), .ZN(n1197) );
XOR2_X1 U855 ( .A(n1200), .B(n1201), .Z(n1198) );
NOR2_X1 U856 ( .A1(KEYINPUT63), .A2(G101), .ZN(n1201) );
NAND2_X1 U857 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
NAND2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND2_X1 U859 ( .A1(KEYINPUT45), .A2(n1206), .ZN(n1204) );
NAND2_X1 U860 ( .A1(KEYINPUT17), .A2(n1207), .ZN(n1206) );
NAND2_X1 U861 ( .A1(n1208), .A2(n1209), .ZN(n1202) );
NAND2_X1 U862 ( .A1(KEYINPUT17), .A2(n1210), .ZN(n1209) );
NAND2_X1 U863 ( .A1(n1211), .A2(KEYINPUT45), .ZN(n1210) );
INV_X1 U864 ( .A(n1205), .ZN(n1211) );
NAND2_X1 U865 ( .A1(n1190), .A2(G472), .ZN(n1205) );
INV_X1 U866 ( .A(n1207), .ZN(n1208) );
XNOR2_X1 U867 ( .A(n1212), .B(n1213), .ZN(n1207) );
NOR3_X1 U868 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NOR2_X1 U869 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XNOR2_X1 U870 ( .A(KEYINPUT19), .B(n1219), .ZN(n1217) );
AND3_X1 U871 ( .A1(n1218), .A2(n1220), .A3(n1221), .ZN(n1215) );
INV_X1 U872 ( .A(KEYINPUT52), .ZN(n1218) );
NOR2_X1 U873 ( .A1(n1221), .A2(n1220), .ZN(n1214) );
NOR2_X1 U874 ( .A1(KEYINPUT38), .A2(n1222), .ZN(n1221) );
XNOR2_X1 U875 ( .A(KEYINPUT19), .B(n1223), .ZN(n1222) );
NAND2_X1 U876 ( .A1(KEYINPUT32), .A2(n1224), .ZN(n1212) );
NOR2_X1 U877 ( .A1(n1180), .A2(n1225), .ZN(G54) );
XOR2_X1 U878 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U879 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U880 ( .A(n1230), .B(n1231), .Z(n1226) );
AND2_X1 U881 ( .A1(G469), .A2(n1190), .ZN(n1231) );
INV_X1 U882 ( .A(n1185), .ZN(n1190) );
XNOR2_X1 U883 ( .A(G110), .B(KEYINPUT33), .ZN(n1230) );
NOR2_X1 U884 ( .A1(n1180), .A2(n1232), .ZN(G51) );
NOR3_X1 U885 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
NOR3_X1 U886 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
NOR3_X1 U887 ( .A1(n1185), .A2(KEYINPUT40), .A3(n1239), .ZN(n1237) );
NOR2_X1 U888 ( .A1(KEYINPUT10), .A2(n1240), .ZN(n1234) );
NOR3_X1 U889 ( .A1(n1185), .A2(n1241), .A3(n1239), .ZN(n1233) );
NOR2_X1 U890 ( .A1(n1242), .A2(n1236), .ZN(n1241) );
INV_X1 U891 ( .A(KEYINPUT10), .ZN(n1236) );
NOR2_X1 U892 ( .A1(KEYINPUT40), .A2(n1240), .ZN(n1242) );
INV_X1 U893 ( .A(n1238), .ZN(n1240) );
XNOR2_X1 U894 ( .A(n1243), .B(n1244), .ZN(n1238) );
NAND2_X1 U895 ( .A1(KEYINPUT34), .A2(n1245), .ZN(n1243) );
NAND2_X1 U896 ( .A1(G902), .A2(n1089), .ZN(n1185) );
NAND2_X1 U897 ( .A1(n1156), .A2(n1173), .ZN(n1089) );
AND4_X1 U898 ( .A1(n1246), .A2(n1084), .A3(n1247), .A4(n1248), .ZN(n1173) );
NOR4_X1 U899 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1248) );
NOR2_X1 U900 ( .A1(n1253), .A2(n1254), .ZN(n1247) );
NOR2_X1 U901 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U902 ( .A(KEYINPUT48), .B(n1257), .ZN(n1256) );
INV_X1 U903 ( .A(n1196), .ZN(n1255) );
NOR3_X1 U904 ( .A1(n1099), .A2(n1258), .A3(n1259), .ZN(n1253) );
NAND2_X1 U905 ( .A1(n1111), .A2(n1196), .ZN(n1084) );
NOR3_X1 U906 ( .A1(n1093), .A2(n1094), .A3(n1258), .ZN(n1196) );
AND4_X1 U907 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1156) );
AND4_X1 U908 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1263) );
OR2_X1 U909 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U910 ( .A(n1270), .B(KEYINPUT2), .ZN(n1268) );
AND2_X1 U911 ( .A1(n1271), .A2(n1272), .ZN(n1262) );
NAND2_X1 U912 ( .A1(n1273), .A2(n1274), .ZN(n1260) );
XNOR2_X1 U913 ( .A(KEYINPUT9), .B(n1107), .ZN(n1274) );
NOR2_X1 U914 ( .A1(n1114), .A2(G952), .ZN(n1180) );
NAND2_X1 U915 ( .A1(n1275), .A2(n1276), .ZN(G48) );
NAND2_X1 U916 ( .A1(KEYINPUT62), .A2(n1277), .ZN(n1276) );
XOR2_X1 U917 ( .A(n1278), .B(n1279), .Z(n1275) );
NOR2_X1 U918 ( .A1(n1280), .A2(n1269), .ZN(n1279) );
NAND3_X1 U919 ( .A1(n1112), .A2(n1281), .A3(n1282), .ZN(n1269) );
OR2_X1 U920 ( .A1(n1277), .A2(KEYINPUT62), .ZN(n1278) );
XNOR2_X1 U921 ( .A(n1283), .B(n1284), .ZN(G45) );
NOR2_X1 U922 ( .A1(KEYINPUT14), .A2(n1266), .ZN(n1284) );
NAND3_X1 U923 ( .A1(n1121), .A2(n1282), .A3(n1285), .ZN(n1266) );
XNOR2_X1 U924 ( .A(G140), .B(n1265), .ZN(G42) );
NAND4_X1 U925 ( .A1(n1282), .A2(n1119), .A3(n1123), .A4(n1112), .ZN(n1265) );
XNOR2_X1 U926 ( .A(n1261), .B(n1286), .ZN(G39) );
NOR2_X1 U927 ( .A1(KEYINPUT4), .A2(n1168), .ZN(n1286) );
NAND4_X1 U928 ( .A1(n1117), .A2(n1270), .A3(n1282), .A4(n1119), .ZN(n1261) );
XNOR2_X1 U929 ( .A(n1167), .B(n1287), .ZN(G36) );
NOR2_X1 U930 ( .A1(n1288), .A2(n1107), .ZN(n1287) );
INV_X1 U931 ( .A(n1119), .ZN(n1107) );
XNOR2_X1 U932 ( .A(n1273), .B(KEYINPUT15), .ZN(n1288) );
AND3_X1 U933 ( .A1(n1282), .A2(n1111), .A3(n1121), .ZN(n1273) );
XNOR2_X1 U934 ( .A(G131), .B(n1272), .ZN(G33) );
NAND4_X1 U935 ( .A1(n1121), .A2(n1282), .A3(n1119), .A4(n1112), .ZN(n1272) );
NOR2_X1 U936 ( .A1(n1105), .A2(n1289), .ZN(n1119) );
INV_X1 U937 ( .A(n1103), .ZN(n1289) );
XNOR2_X1 U938 ( .A(G128), .B(n1264), .ZN(G30) );
NAND4_X1 U939 ( .A1(n1270), .A2(n1282), .A3(n1111), .A4(n1281), .ZN(n1264) );
AND3_X1 U940 ( .A1(n1290), .A2(n1291), .A3(n1109), .ZN(n1282) );
XNOR2_X1 U941 ( .A(n1252), .B(n1292), .ZN(G3) );
NAND2_X1 U942 ( .A1(KEYINPUT47), .A2(G101), .ZN(n1292) );
NOR3_X1 U943 ( .A1(n1293), .A2(n1258), .A3(n1099), .ZN(n1252) );
XOR2_X1 U944 ( .A(n1271), .B(n1294), .Z(G27) );
NAND2_X1 U945 ( .A1(KEYINPUT51), .A2(G125), .ZN(n1294) );
NAND4_X1 U946 ( .A1(n1123), .A2(n1101), .A3(n1112), .A4(n1290), .ZN(n1271) );
NAND2_X1 U947 ( .A1(n1095), .A2(n1295), .ZN(n1290) );
NAND2_X1 U948 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
INV_X1 U949 ( .A(G900), .ZN(n1297) );
INV_X1 U950 ( .A(n1257), .ZN(n1112) );
INV_X1 U951 ( .A(n1259), .ZN(n1123) );
NAND2_X1 U952 ( .A1(n1298), .A2(n1299), .ZN(G24) );
NAND2_X1 U953 ( .A1(G122), .A2(n1246), .ZN(n1299) );
XOR2_X1 U954 ( .A(n1300), .B(KEYINPUT0), .Z(n1298) );
OR2_X1 U955 ( .A1(n1246), .A2(G122), .ZN(n1300) );
NAND3_X1 U956 ( .A1(n1285), .A2(n1133), .A3(n1301), .ZN(n1246) );
NOR3_X1 U957 ( .A1(n1094), .A2(n1302), .A3(n1093), .ZN(n1301) );
INV_X1 U958 ( .A(n1303), .ZN(n1302) );
AND3_X1 U959 ( .A1(n1304), .A2(n1132), .A3(n1281), .ZN(n1285) );
XNOR2_X1 U960 ( .A(n1251), .B(n1305), .ZN(G21) );
XNOR2_X1 U961 ( .A(G119), .B(KEYINPUT1), .ZN(n1305) );
AND4_X1 U962 ( .A1(n1117), .A2(n1270), .A3(n1101), .A4(n1303), .ZN(n1251) );
INV_X1 U963 ( .A(n1280), .ZN(n1270) );
NAND2_X1 U964 ( .A1(n1093), .A2(n1094), .ZN(n1280) );
XNOR2_X1 U965 ( .A(G116), .B(n1306), .ZN(G18) );
NOR2_X1 U966 ( .A1(n1250), .A2(KEYINPUT27), .ZN(n1306) );
AND4_X1 U967 ( .A1(n1121), .A2(n1101), .A3(n1111), .A4(n1303), .ZN(n1250) );
NOR2_X1 U968 ( .A1(n1132), .A2(n1307), .ZN(n1111) );
AND2_X1 U969 ( .A1(n1133), .A2(n1281), .ZN(n1101) );
NAND2_X1 U970 ( .A1(n1308), .A2(n1309), .ZN(G15) );
NAND2_X1 U971 ( .A1(n1249), .A2(n1310), .ZN(n1309) );
XOR2_X1 U972 ( .A(KEYINPUT20), .B(n1311), .Z(n1308) );
NOR2_X1 U973 ( .A1(n1249), .A2(n1310), .ZN(n1311) );
INV_X1 U974 ( .A(G113), .ZN(n1310) );
AND4_X1 U975 ( .A1(n1312), .A2(n1303), .A3(n1133), .A4(n1313), .ZN(n1249) );
NOR2_X1 U976 ( .A1(n1257), .A2(n1293), .ZN(n1313) );
INV_X1 U977 ( .A(n1121), .ZN(n1293) );
NOR2_X1 U978 ( .A1(n1094), .A2(n1314), .ZN(n1121) );
NAND2_X1 U979 ( .A1(n1307), .A2(n1132), .ZN(n1257) );
NOR2_X1 U980 ( .A1(n1109), .A2(n1108), .ZN(n1133) );
INV_X1 U981 ( .A(n1291), .ZN(n1108) );
XNOR2_X1 U982 ( .A(n1315), .B(n1316), .ZN(G12) );
NOR3_X1 U983 ( .A1(n1317), .A2(n1258), .A3(n1259), .ZN(n1316) );
NAND2_X1 U984 ( .A1(n1314), .A2(n1094), .ZN(n1259) );
NAND2_X1 U985 ( .A1(n1139), .A2(n1145), .ZN(n1094) );
NAND3_X1 U986 ( .A1(n1318), .A2(n1319), .A3(n1182), .ZN(n1145) );
NAND2_X1 U987 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
NAND2_X1 U988 ( .A1(n1320), .A2(n1322), .ZN(n1139) );
NAND2_X1 U989 ( .A1(n1323), .A2(n1319), .ZN(n1322) );
NAND2_X1 U990 ( .A1(n1324), .A2(n1321), .ZN(n1323) );
INV_X1 U991 ( .A(n1182), .ZN(n1324) );
XNOR2_X1 U992 ( .A(n1325), .B(n1326), .ZN(n1182) );
XNOR2_X1 U993 ( .A(n1315), .B(n1327), .ZN(n1326) );
XNOR2_X1 U994 ( .A(n1277), .B(G137), .ZN(n1327) );
INV_X1 U995 ( .A(G146), .ZN(n1277) );
XNOR2_X1 U996 ( .A(n1161), .B(n1328), .ZN(n1325) );
XNOR2_X1 U997 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U998 ( .A1(G119), .A2(KEYINPUT7), .ZN(n1330) );
NAND2_X1 U999 ( .A1(KEYINPUT49), .A2(n1331), .ZN(n1329) );
NAND3_X1 U1000 ( .A1(G234), .A2(n1114), .A3(G221), .ZN(n1331) );
XOR2_X1 U1001 ( .A(G125), .B(n1228), .Z(n1161) );
XNOR2_X1 U1002 ( .A(n1332), .B(G140), .ZN(n1228) );
XNOR2_X1 U1003 ( .A(KEYINPUT29), .B(n1184), .ZN(n1320) );
INV_X1 U1004 ( .A(n1093), .ZN(n1314) );
XNOR2_X1 U1005 ( .A(n1135), .B(G472), .ZN(n1093) );
NAND2_X1 U1006 ( .A1(n1333), .A2(n1319), .ZN(n1135) );
XOR2_X1 U1007 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1008 ( .A(n1336), .B(n1224), .Z(n1335) );
XNOR2_X1 U1009 ( .A(G113), .B(n1337), .ZN(n1224) );
NAND2_X1 U1010 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
NAND2_X1 U1011 ( .A1(n1220), .A2(n1340), .ZN(n1339) );
NAND2_X1 U1012 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1013 ( .A1(KEYINPUT56), .A2(n1223), .ZN(n1342) );
NAND2_X1 U1014 ( .A1(n1219), .A2(n1343), .ZN(n1338) );
NAND2_X1 U1015 ( .A1(KEYINPUT56), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1016 ( .A1(n1345), .A2(n1341), .ZN(n1344) );
INV_X1 U1017 ( .A(KEYINPUT53), .ZN(n1341) );
INV_X1 U1018 ( .A(n1223), .ZN(n1219) );
XOR2_X1 U1019 ( .A(n1199), .B(G101), .Z(n1334) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1346), .ZN(n1199) );
NAND4_X1 U1021 ( .A1(n1312), .A2(n1109), .A3(n1303), .A4(n1291), .ZN(n1258) );
NAND2_X1 U1022 ( .A1(G221), .A2(n1347), .ZN(n1291) );
NAND2_X1 U1023 ( .A1(G234), .A2(n1319), .ZN(n1347) );
NAND2_X1 U1024 ( .A1(n1095), .A2(n1348), .ZN(n1303) );
NAND2_X1 U1025 ( .A1(n1296), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1026 ( .A(KEYINPUT35), .B(G898), .Z(n1349) );
AND3_X1 U1027 ( .A1(n1350), .A2(n1351), .A3(G953), .ZN(n1296) );
XNOR2_X1 U1028 ( .A(KEYINPUT42), .B(n1319), .ZN(n1350) );
NAND3_X1 U1029 ( .A1(n1351), .A2(n1114), .A3(G952), .ZN(n1095) );
NAND2_X1 U1030 ( .A1(G237), .A2(G234), .ZN(n1351) );
XNOR2_X1 U1031 ( .A(n1352), .B(G469), .ZN(n1109) );
NAND2_X1 U1032 ( .A1(n1353), .A2(n1319), .ZN(n1352) );
XOR2_X1 U1033 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1034 ( .A(n1229), .B(G128), .ZN(n1355) );
XNOR2_X1 U1035 ( .A(n1356), .B(n1357), .ZN(n1229) );
XNOR2_X1 U1036 ( .A(n1220), .B(n1358), .ZN(n1357) );
NAND2_X1 U1037 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
OR2_X1 U1038 ( .A1(n1361), .A2(G101), .ZN(n1360) );
XOR2_X1 U1039 ( .A(n1362), .B(KEYINPUT21), .Z(n1359) );
NAND2_X1 U1040 ( .A1(G101), .A2(n1361), .ZN(n1362) );
XOR2_X1 U1041 ( .A(n1363), .B(n1085), .Z(n1361) );
NAND2_X1 U1042 ( .A1(KEYINPUT54), .A2(G104), .ZN(n1363) );
INV_X1 U1043 ( .A(n1345), .ZN(n1220) );
NAND2_X1 U1044 ( .A1(n1364), .A2(n1365), .ZN(n1345) );
NAND2_X1 U1045 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NAND2_X1 U1046 ( .A1(G134), .A2(n1368), .ZN(n1367) );
XNOR2_X1 U1047 ( .A(G131), .B(G137), .ZN(n1366) );
NAND2_X1 U1048 ( .A1(n1369), .A2(n1368), .ZN(n1364) );
INV_X1 U1049 ( .A(KEYINPUT50), .ZN(n1368) );
NAND2_X1 U1050 ( .A1(n1163), .A2(n1162), .ZN(n1369) );
NAND3_X1 U1051 ( .A1(G131), .A2(n1168), .A3(G134), .ZN(n1162) );
INV_X1 U1052 ( .A(G137), .ZN(n1168) );
NAND3_X1 U1053 ( .A1(G134), .A2(n1166), .A3(G137), .ZN(n1163) );
INV_X1 U1054 ( .A(G131), .ZN(n1166) );
XOR2_X1 U1055 ( .A(n1370), .B(n1159), .Z(n1356) );
NOR2_X1 U1056 ( .A1(KEYINPUT24), .A2(n1371), .ZN(n1159) );
XNOR2_X1 U1057 ( .A(G143), .B(G146), .ZN(n1371) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1114), .ZN(n1370) );
NAND2_X1 U1059 ( .A1(n1372), .A2(n1373), .ZN(n1354) );
NAND2_X1 U1060 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
INV_X1 U1061 ( .A(KEYINPUT13), .ZN(n1375) );
XNOR2_X1 U1062 ( .A(G110), .B(G140), .ZN(n1374) );
NAND3_X1 U1063 ( .A1(G140), .A2(n1315), .A3(KEYINPUT13), .ZN(n1372) );
XNOR2_X1 U1064 ( .A(n1281), .B(KEYINPUT31), .ZN(n1312) );
AND2_X1 U1065 ( .A1(n1103), .A2(n1105), .ZN(n1281) );
NAND3_X1 U1066 ( .A1(n1376), .A2(n1377), .A3(n1146), .ZN(n1105) );
OR2_X1 U1067 ( .A1(n1148), .A2(n1147), .ZN(n1146) );
OR2_X1 U1068 ( .A1(n1147), .A2(KEYINPUT46), .ZN(n1377) );
NAND3_X1 U1069 ( .A1(n1147), .A2(n1148), .A3(KEYINPUT46), .ZN(n1376) );
NAND2_X1 U1070 ( .A1(n1378), .A2(n1319), .ZN(n1148) );
XOR2_X1 U1071 ( .A(n1379), .B(n1244), .Z(n1378) );
XNOR2_X1 U1072 ( .A(n1380), .B(n1223), .ZN(n1244) );
XNOR2_X1 U1073 ( .A(n1381), .B(n1382), .ZN(n1223) );
NOR2_X1 U1074 ( .A1(G146), .A2(KEYINPUT44), .ZN(n1382) );
XNOR2_X1 U1075 ( .A(G143), .B(n1383), .ZN(n1381) );
NOR2_X1 U1076 ( .A1(KEYINPUT61), .A2(n1332), .ZN(n1383) );
INV_X1 U1077 ( .A(G128), .ZN(n1332) );
XNOR2_X1 U1078 ( .A(G125), .B(n1384), .ZN(n1380) );
AND2_X1 U1079 ( .A1(n1114), .A2(G224), .ZN(n1384) );
INV_X1 U1080 ( .A(G953), .ZN(n1114) );
XOR2_X1 U1081 ( .A(n1245), .B(KEYINPUT55), .Z(n1379) );
XOR2_X1 U1082 ( .A(n1178), .B(n1385), .Z(n1245) );
NOR2_X1 U1083 ( .A1(KEYINPUT43), .A2(n1179), .ZN(n1385) );
XNOR2_X1 U1084 ( .A(n1315), .B(n1386), .ZN(n1179) );
NOR2_X1 U1085 ( .A1(G122), .A2(KEYINPUT41), .ZN(n1386) );
XOR2_X1 U1086 ( .A(n1387), .B(n1388), .Z(n1178) );
XNOR2_X1 U1087 ( .A(n1085), .B(G101), .ZN(n1388) );
INV_X1 U1088 ( .A(G107), .ZN(n1085) );
XOR2_X1 U1089 ( .A(n1389), .B(n1390), .Z(n1387) );
NOR2_X1 U1090 ( .A1(G104), .A2(KEYINPUT23), .ZN(n1390) );
NAND2_X1 U1091 ( .A1(n1391), .A2(n1392), .ZN(n1389) );
NAND2_X1 U1092 ( .A1(G113), .A2(n1337), .ZN(n1392) );
XOR2_X1 U1093 ( .A(KEYINPUT37), .B(n1393), .Z(n1391) );
NOR2_X1 U1094 ( .A1(G113), .A2(n1337), .ZN(n1393) );
XNOR2_X1 U1095 ( .A(n1394), .B(G119), .ZN(n1337) );
INV_X1 U1096 ( .A(n1239), .ZN(n1147) );
NAND2_X1 U1097 ( .A1(G210), .A2(n1395), .ZN(n1239) );
NAND2_X1 U1098 ( .A1(G214), .A2(n1395), .ZN(n1103) );
NAND2_X1 U1099 ( .A1(n1396), .A2(n1319), .ZN(n1395) );
INV_X1 U1100 ( .A(G902), .ZN(n1319) );
INV_X1 U1101 ( .A(G237), .ZN(n1396) );
XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1099), .ZN(n1317) );
INV_X1 U1103 ( .A(n1117), .ZN(n1099) );
NOR2_X1 U1104 ( .A1(n1132), .A2(n1304), .ZN(n1117) );
INV_X1 U1105 ( .A(n1307), .ZN(n1304) );
XOR2_X1 U1106 ( .A(n1397), .B(n1142), .Z(n1307) );
INV_X1 U1107 ( .A(n1144), .ZN(n1142) );
NOR2_X1 U1108 ( .A1(n1189), .A2(G902), .ZN(n1144) );
XOR2_X1 U1109 ( .A(n1398), .B(n1399), .Z(n1189) );
XOR2_X1 U1110 ( .A(n1400), .B(n1401), .Z(n1399) );
XNOR2_X1 U1111 ( .A(n1402), .B(n1403), .ZN(n1401) );
NOR2_X1 U1112 ( .A1(KEYINPUT26), .A2(n1404), .ZN(n1403) );
XNOR2_X1 U1113 ( .A(n1283), .B(G128), .ZN(n1404) );
NAND2_X1 U1114 ( .A1(KEYINPUT18), .A2(n1394), .ZN(n1402) );
INV_X1 U1115 ( .A(G116), .ZN(n1394) );
NOR4_X1 U1116 ( .A1(KEYINPUT12), .A2(G953), .A3(n1184), .A4(n1321), .ZN(n1400) );
INV_X1 U1117 ( .A(G234), .ZN(n1321) );
INV_X1 U1118 ( .A(G217), .ZN(n1184) );
XNOR2_X1 U1119 ( .A(G107), .B(n1405), .ZN(n1398) );
XNOR2_X1 U1120 ( .A(n1167), .B(G122), .ZN(n1405) );
INV_X1 U1121 ( .A(G134), .ZN(n1167) );
NAND2_X1 U1122 ( .A1(KEYINPUT57), .A2(n1141), .ZN(n1397) );
INV_X1 U1123 ( .A(G478), .ZN(n1141) );
XNOR2_X1 U1124 ( .A(n1406), .B(G475), .ZN(n1132) );
OR2_X1 U1125 ( .A1(n1194), .A2(G902), .ZN(n1406) );
XNOR2_X1 U1126 ( .A(n1407), .B(n1408), .ZN(n1194) );
XOR2_X1 U1127 ( .A(n1409), .B(n1410), .Z(n1408) );
XOR2_X1 U1128 ( .A(n1411), .B(n1412), .Z(n1410) );
NOR2_X1 U1129 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
XOR2_X1 U1130 ( .A(n1415), .B(KEYINPUT39), .Z(n1414) );
NAND2_X1 U1131 ( .A1(G146), .A2(n1416), .ZN(n1415) );
NOR2_X1 U1132 ( .A1(G146), .A2(n1416), .ZN(n1413) );
NAND3_X1 U1133 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1416) );
NAND2_X1 U1134 ( .A1(G140), .A2(n1420), .ZN(n1419) );
NAND2_X1 U1135 ( .A1(KEYINPUT16), .A2(n1421), .ZN(n1418) );
NAND2_X1 U1136 ( .A1(n1422), .A2(n1423), .ZN(n1421) );
INV_X1 U1137 ( .A(G140), .ZN(n1423) );
XNOR2_X1 U1138 ( .A(KEYINPUT25), .B(n1420), .ZN(n1422) );
NAND2_X1 U1139 ( .A1(n1424), .A2(n1425), .ZN(n1417) );
INV_X1 U1140 ( .A(KEYINPUT16), .ZN(n1425) );
NAND2_X1 U1141 ( .A1(n1426), .A2(n1427), .ZN(n1424) );
OR3_X1 U1142 ( .A1(n1420), .A2(G140), .A3(KEYINPUT25), .ZN(n1427) );
NAND2_X1 U1143 ( .A1(KEYINPUT25), .A2(n1420), .ZN(n1426) );
INV_X1 U1144 ( .A(G125), .ZN(n1420) );
NOR2_X1 U1145 ( .A1(KEYINPUT8), .A2(G122), .ZN(n1411) );
AND2_X1 U1146 ( .A1(n1346), .A2(G214), .ZN(n1409) );
NOR2_X1 U1147 ( .A1(G953), .A2(G237), .ZN(n1346) );
XOR2_X1 U1148 ( .A(n1428), .B(n1429), .Z(n1407) );
XNOR2_X1 U1149 ( .A(n1283), .B(G131), .ZN(n1429) );
INV_X1 U1150 ( .A(G143), .ZN(n1283) );
XNOR2_X1 U1151 ( .A(G104), .B(G113), .ZN(n1428) );
INV_X1 U1152 ( .A(G110), .ZN(n1315) );
endmodule


