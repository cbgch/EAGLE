//Key = 1100001010100000111100110000001111100111000100001111111100010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;

XNOR2_X1 U751 ( .A(G107), .B(n1031), .ZN(G9) );
NOR2_X1 U752 ( .A1(n1032), .A2(n1033), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1034), .A2(n1035), .A3(G953), .A4(n1036), .ZN(n1033) );
NAND3_X1 U754 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1034) );
XOR2_X1 U755 ( .A(n1040), .B(KEYINPUT31), .Z(n1039) );
NAND2_X1 U756 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND4_X1 U757 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NAND3_X1 U758 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND3_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1048) );
XOR2_X1 U761 ( .A(KEYINPUT56), .B(n1050), .Z(n1053) );
NAND2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1047) );
NAND2_X1 U763 ( .A1(n1055), .A2(n1057), .ZN(n1041) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND4_X1 U765 ( .A1(n1044), .A2(n1060), .A3(n1045), .A4(n1061), .ZN(n1059) );
XNOR2_X1 U766 ( .A(KEYINPUT13), .B(n1062), .ZN(n1061) );
NAND4_X1 U767 ( .A1(n1043), .A2(n1050), .A3(n1063), .A4(n1064), .ZN(n1058) );
NAND2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1045), .A2(n1067), .ZN(n1065) );
NAND2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
OR3_X1 U771 ( .A1(n1070), .A2(n1071), .A3(n1066), .ZN(n1063) );
INV_X1 U772 ( .A(n1044), .ZN(n1066) );
INV_X1 U773 ( .A(n1062), .ZN(n1043) );
NOR3_X1 U774 ( .A1(n1036), .A2(G953), .A3(G952), .ZN(n1032) );
AND4_X1 U775 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1036) );
NOR4_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
INV_X1 U778 ( .A(KEYINPUT42), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
INV_X1 U780 ( .A(n1084), .ZN(n1082) );
NOR3_X1 U781 ( .A1(KEYINPUT42), .A2(n1085), .A3(n1083), .ZN(n1078) );
XNOR2_X1 U782 ( .A(n1086), .B(n1087), .ZN(n1077) );
NAND3_X1 U783 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1076) );
XOR2_X1 U784 ( .A(G469), .B(n1091), .Z(n1089) );
NOR2_X1 U785 ( .A1(n1092), .A2(KEYINPUT41), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1085), .A2(n1083), .ZN(n1088) );
XNOR2_X1 U787 ( .A(n1093), .B(KEYINPUT25), .ZN(n1083) );
NOR2_X1 U788 ( .A1(n1084), .A2(KEYINPUT40), .ZN(n1085) );
NOR3_X1 U789 ( .A1(n1054), .A2(n1094), .A3(n1095), .ZN(n1074) );
XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(n1072) );
NAND2_X1 U791 ( .A1(KEYINPUT6), .A2(n1098), .ZN(n1097) );
XOR2_X1 U792 ( .A(n1099), .B(n1100), .Z(G72) );
NAND2_X1 U793 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND4_X1 U794 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
NAND2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
NAND3_X1 U796 ( .A1(n1109), .A2(n1108), .A3(n1107), .ZN(n1101) );
NAND2_X1 U797 ( .A1(n1037), .A2(n1110), .ZN(n1107) );
NAND2_X1 U798 ( .A1(n1103), .A2(n1105), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1105) );
XNOR2_X1 U800 ( .A(KEYINPUT63), .B(n1113), .ZN(n1103) );
OR2_X1 U801 ( .A1(n1112), .A2(n1111), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1111) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1114) );
NAND2_X1 U804 ( .A1(KEYINPUT39), .A2(n1118), .ZN(n1116) );
INV_X1 U805 ( .A(n1119), .ZN(n1118) );
NAND2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(n1112) );
NAND2_X1 U807 ( .A1(KEYINPUT16), .A2(n1122), .ZN(n1121) );
OR3_X1 U808 ( .A1(n1123), .A2(G125), .A3(KEYINPUT16), .ZN(n1120) );
NAND2_X1 U809 ( .A1(n1106), .A2(n1124), .ZN(n1099) );
OR2_X1 U810 ( .A1(n1108), .A2(G227), .ZN(n1124) );
INV_X1 U811 ( .A(n1125), .ZN(n1106) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1108), .ZN(n1127) );
AND2_X1 U814 ( .A1(G224), .A2(G898), .ZN(n1128) );
NOR2_X1 U815 ( .A1(KEYINPUT58), .A2(n1129), .ZN(n1126) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U817 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U818 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U819 ( .A(n1136), .B(n1137), .ZN(n1135) );
XOR2_X1 U820 ( .A(KEYINPUT49), .B(n1138), .Z(n1134) );
NOR2_X1 U821 ( .A1(KEYINPUT3), .A2(n1139), .ZN(n1138) );
NOR2_X1 U822 ( .A1(G898), .A2(n1108), .ZN(n1132) );
NAND2_X1 U823 ( .A1(n1108), .A2(n1140), .ZN(n1130) );
NOR2_X1 U824 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
AND2_X1 U826 ( .A1(G217), .A2(n1145), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1141), .A2(n1146), .ZN(G63) );
XNOR2_X1 U828 ( .A(n1147), .B(n1148), .ZN(n1146) );
AND2_X1 U829 ( .A1(G478), .A2(n1145), .ZN(n1148) );
NOR2_X1 U830 ( .A1(n1141), .A2(n1149), .ZN(G60) );
XOR2_X1 U831 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U832 ( .A1(KEYINPUT61), .A2(n1152), .ZN(n1150) );
NAND2_X1 U833 ( .A1(n1145), .A2(G475), .ZN(n1152) );
XNOR2_X1 U834 ( .A(n1153), .B(n1154), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1141), .A2(n1155), .ZN(G57) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U837 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U838 ( .A1(n1098), .A2(n1160), .ZN(n1159) );
NOR2_X1 U839 ( .A1(KEYINPUT44), .A2(n1161), .ZN(n1158) );
XNOR2_X1 U840 ( .A(n1162), .B(n1163), .ZN(n1161) );
XNOR2_X1 U841 ( .A(n1164), .B(KEYINPUT7), .ZN(n1163) );
NOR2_X1 U842 ( .A1(n1141), .A2(n1165), .ZN(G54) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U844 ( .A(n1168), .B(n1169), .Z(n1167) );
AND2_X1 U845 ( .A1(G469), .A2(n1145), .ZN(n1169) );
NOR2_X1 U846 ( .A1(KEYINPUT9), .A2(n1170), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U848 ( .A1(KEYINPUT28), .A2(n1173), .ZN(n1172) );
NOR2_X1 U849 ( .A1(n1141), .A2(n1174), .ZN(G51) );
XNOR2_X1 U850 ( .A(n1175), .B(n1176), .ZN(n1174) );
XNOR2_X1 U851 ( .A(n1177), .B(n1178), .ZN(n1176) );
NAND2_X1 U852 ( .A1(KEYINPUT50), .A2(n1179), .ZN(n1178) );
NAND2_X1 U853 ( .A1(KEYINPUT37), .A2(n1180), .ZN(n1177) );
NAND2_X1 U854 ( .A1(n1145), .A2(n1086), .ZN(n1180) );
INV_X1 U855 ( .A(n1181), .ZN(n1086) );
INV_X1 U856 ( .A(n1160), .ZN(n1145) );
NAND2_X1 U857 ( .A1(G902), .A2(n1182), .ZN(n1160) );
NAND3_X1 U858 ( .A1(n1183), .A2(n1038), .A3(n1037), .ZN(n1182) );
AND4_X1 U859 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1037) );
NAND4_X1 U860 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1056), .ZN(n1184) );
XNOR2_X1 U861 ( .A(n1055), .B(KEYINPUT23), .ZN(n1189) );
XNOR2_X1 U862 ( .A(n1071), .B(KEYINPUT30), .ZN(n1188) );
INV_X1 U863 ( .A(n1140), .ZN(n1038) );
NAND4_X1 U864 ( .A1(n1191), .A2(n1031), .A3(n1192), .A4(n1193), .ZN(n1140) );
NOR4_X1 U865 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1154), .ZN(n1193) );
AND3_X1 U866 ( .A1(n1197), .A2(n1045), .A3(n1056), .ZN(n1154) );
NOR3_X1 U867 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1192) );
NOR3_X1 U868 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
NAND3_X1 U869 ( .A1(n1044), .A2(n1204), .A3(n1050), .ZN(n1203) );
NAND3_X1 U870 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1202) );
INV_X1 U871 ( .A(KEYINPUT57), .ZN(n1201) );
NOR2_X1 U872 ( .A1(KEYINPUT57), .A2(n1208), .ZN(n1199) );
NAND3_X1 U873 ( .A1(n1060), .A2(n1045), .A3(n1197), .ZN(n1031) );
INV_X1 U874 ( .A(n1035), .ZN(n1183) );
XOR2_X1 U875 ( .A(n1110), .B(KEYINPUT62), .Z(n1035) );
AND3_X1 U876 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1110) );
NAND2_X1 U877 ( .A1(n1051), .A2(n1212), .ZN(n1211) );
NAND2_X1 U878 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U879 ( .A(KEYINPUT0), .B(n1215), .ZN(n1213) );
NOR2_X1 U880 ( .A1(n1108), .A2(G952), .ZN(n1141) );
XNOR2_X1 U881 ( .A(n1216), .B(n1217), .ZN(G48) );
NOR3_X1 U882 ( .A1(n1215), .A2(KEYINPUT4), .A3(n1206), .ZN(n1217) );
NAND2_X1 U883 ( .A1(n1218), .A2(n1056), .ZN(n1215) );
XNOR2_X1 U884 ( .A(G143), .B(n1219), .ZN(G45) );
NAND2_X1 U885 ( .A1(n1220), .A2(n1051), .ZN(n1219) );
XOR2_X1 U886 ( .A(n1214), .B(KEYINPUT43), .Z(n1220) );
NAND4_X1 U887 ( .A1(n1071), .A2(n1190), .A3(n1221), .A4(n1222), .ZN(n1214) );
XNOR2_X1 U888 ( .A(G140), .B(n1209), .ZN(G42) );
NAND4_X1 U889 ( .A1(n1055), .A2(n1190), .A3(n1056), .A4(n1070), .ZN(n1209) );
XNOR2_X1 U890 ( .A(G137), .B(n1210), .ZN(G39) );
NAND3_X1 U891 ( .A1(n1055), .A2(n1218), .A3(n1050), .ZN(n1210) );
XNOR2_X1 U892 ( .A(G134), .B(n1185), .ZN(G36) );
NAND4_X1 U893 ( .A1(n1071), .A2(n1055), .A3(n1190), .A4(n1060), .ZN(n1185) );
XOR2_X1 U894 ( .A(n1223), .B(G131), .Z(G33) );
NAND2_X1 U895 ( .A1(KEYINPUT32), .A2(n1224), .ZN(n1223) );
NAND4_X1 U896 ( .A1(n1071), .A2(n1055), .A3(n1190), .A4(n1056), .ZN(n1224) );
NOR2_X1 U897 ( .A1(n1225), .A2(n1054), .ZN(n1055) );
XNOR2_X1 U898 ( .A(G128), .B(n1186), .ZN(G30) );
NAND3_X1 U899 ( .A1(n1060), .A2(n1051), .A3(n1218), .ZN(n1186) );
AND3_X1 U900 ( .A1(n1204), .A2(n1207), .A3(n1190), .ZN(n1218) );
NOR3_X1 U901 ( .A1(n1226), .A2(n1068), .A3(n1227), .ZN(n1190) );
XNOR2_X1 U902 ( .A(n1228), .B(n1198), .ZN(G3) );
AND3_X1 U903 ( .A1(n1071), .A2(n1197), .A3(n1050), .ZN(n1198) );
XNOR2_X1 U904 ( .A(n1179), .B(n1229), .ZN(G27) );
NOR2_X1 U905 ( .A1(KEYINPUT14), .A2(n1187), .ZN(n1229) );
NAND4_X1 U906 ( .A1(n1056), .A2(n1044), .A3(n1230), .A4(n1070), .ZN(n1187) );
NOR2_X1 U907 ( .A1(n1226), .A2(n1206), .ZN(n1230) );
INV_X1 U908 ( .A(n1051), .ZN(n1206) );
AND2_X1 U909 ( .A1(n1062), .A2(n1231), .ZN(n1226) );
NAND3_X1 U910 ( .A1(G902), .A2(n1232), .A3(n1125), .ZN(n1231) );
NOR2_X1 U911 ( .A1(G900), .A2(n1108), .ZN(n1125) );
XOR2_X1 U912 ( .A(n1191), .B(n1233), .Z(G24) );
XNOR2_X1 U913 ( .A(G122), .B(KEYINPUT11), .ZN(n1233) );
NAND4_X1 U914 ( .A1(n1234), .A2(n1045), .A3(n1221), .A4(n1222), .ZN(n1191) );
NOR2_X1 U915 ( .A1(n1207), .A2(n1204), .ZN(n1045) );
NAND2_X1 U916 ( .A1(n1235), .A2(n1236), .ZN(G21) );
NAND2_X1 U917 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U918 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
NAND2_X1 U919 ( .A1(KEYINPUT35), .A2(n1208), .ZN(n1240) );
NAND2_X1 U920 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
INV_X1 U921 ( .A(KEYINPUT35), .ZN(n1242) );
OR2_X1 U922 ( .A1(n1241), .A2(n1238), .ZN(n1235) );
NAND2_X1 U923 ( .A1(KEYINPUT33), .A2(n1208), .ZN(n1241) );
NAND4_X1 U924 ( .A1(n1234), .A2(n1050), .A3(n1204), .A4(n1207), .ZN(n1208) );
XOR2_X1 U925 ( .A(G116), .B(n1196), .Z(G18) );
AND3_X1 U926 ( .A1(n1071), .A2(n1060), .A3(n1234), .ZN(n1196) );
NOR2_X1 U927 ( .A1(n1221), .A2(n1243), .ZN(n1060) );
XOR2_X1 U928 ( .A(G113), .B(n1195), .Z(G15) );
AND3_X1 U929 ( .A1(n1071), .A2(n1056), .A3(n1234), .ZN(n1195) );
AND3_X1 U930 ( .A1(n1051), .A2(n1205), .A3(n1044), .ZN(n1234) );
NOR2_X1 U931 ( .A1(n1069), .A2(n1068), .ZN(n1044) );
AND2_X1 U932 ( .A1(n1243), .A2(n1221), .ZN(n1056) );
AND2_X1 U933 ( .A1(n1090), .A2(n1207), .ZN(n1071) );
XOR2_X1 U934 ( .A(G110), .B(n1194), .Z(G12) );
AND3_X1 U935 ( .A1(n1070), .A2(n1197), .A3(n1050), .ZN(n1194) );
NOR2_X1 U936 ( .A1(n1222), .A2(n1221), .ZN(n1050) );
XNOR2_X1 U937 ( .A(n1084), .B(n1093), .ZN(n1221) );
XNOR2_X1 U938 ( .A(G475), .B(KEYINPUT20), .ZN(n1093) );
NOR2_X1 U939 ( .A1(n1151), .A2(G902), .ZN(n1084) );
XNOR2_X1 U940 ( .A(n1244), .B(n1245), .ZN(n1151) );
XOR2_X1 U941 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U942 ( .A(n1248), .B(G122), .Z(n1247) );
NAND2_X1 U943 ( .A1(n1249), .A2(G214), .ZN(n1248) );
XNOR2_X1 U944 ( .A(G131), .B(G143), .ZN(n1246) );
XOR2_X1 U945 ( .A(n1250), .B(n1251), .Z(n1244) );
XNOR2_X1 U946 ( .A(n1252), .B(n1122), .ZN(n1251) );
NOR2_X1 U947 ( .A1(KEYINPUT21), .A2(n1153), .ZN(n1252) );
INV_X1 U948 ( .A(G104), .ZN(n1153) );
XOR2_X1 U949 ( .A(n1253), .B(n1254), .Z(n1250) );
NOR2_X1 U950 ( .A1(G113), .A2(KEYINPUT45), .ZN(n1254) );
NAND2_X1 U951 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1253) );
INV_X1 U952 ( .A(n1243), .ZN(n1222) );
NOR2_X1 U953 ( .A1(n1255), .A2(n1095), .ZN(n1243) );
NOR3_X1 U954 ( .A1(G478), .A2(G902), .A3(n1256), .ZN(n1095) );
INV_X1 U955 ( .A(n1147), .ZN(n1256) );
XOR2_X1 U956 ( .A(n1094), .B(KEYINPUT26), .Z(n1255) );
AND2_X1 U957 ( .A1(G478), .A2(n1257), .ZN(n1094) );
NAND2_X1 U958 ( .A1(n1147), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U959 ( .A(n1259), .B(n1260), .ZN(n1147) );
XOR2_X1 U960 ( .A(G116), .B(n1261), .Z(n1260) );
XOR2_X1 U961 ( .A(G134), .B(G122), .Z(n1261) );
XOR2_X1 U962 ( .A(n1262), .B(n1263), .Z(n1259) );
XOR2_X1 U963 ( .A(n1264), .B(n1265), .Z(n1262) );
AND3_X1 U964 ( .A1(G217), .A2(n1108), .A3(G234), .ZN(n1265) );
NAND2_X1 U965 ( .A1(KEYINPUT38), .A2(n1266), .ZN(n1264) );
XNOR2_X1 U966 ( .A(n1267), .B(G128), .ZN(n1266) );
AND4_X1 U967 ( .A1(n1051), .A2(n1069), .A3(n1205), .A4(n1073), .ZN(n1197) );
INV_X1 U968 ( .A(n1068), .ZN(n1073) );
NOR2_X1 U969 ( .A1(n1268), .A2(n1269), .ZN(n1068) );
NAND2_X1 U970 ( .A1(n1062), .A2(n1270), .ZN(n1205) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1232), .A4(n1271), .ZN(n1270) );
INV_X1 U972 ( .A(G898), .ZN(n1271) );
NAND3_X1 U973 ( .A1(n1232), .A2(n1108), .A3(G952), .ZN(n1062) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1232) );
INV_X1 U975 ( .A(n1227), .ZN(n1069) );
XNOR2_X1 U976 ( .A(n1092), .B(G469), .ZN(n1227) );
AND3_X1 U977 ( .A1(n1272), .A2(n1273), .A3(n1258), .ZN(n1092) );
NAND2_X1 U978 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
NAND2_X1 U979 ( .A1(n1171), .A2(n1276), .ZN(n1272) );
XOR2_X1 U980 ( .A(n1274), .B(KEYINPUT8), .Z(n1276) );
XNOR2_X1 U981 ( .A(n1173), .B(n1166), .ZN(n1274) );
XNOR2_X1 U982 ( .A(n1277), .B(n1278), .ZN(n1166) );
XNOR2_X1 U983 ( .A(n1123), .B(G110), .ZN(n1278) );
NAND2_X1 U984 ( .A1(G227), .A2(n1108), .ZN(n1277) );
XNOR2_X1 U985 ( .A(n1279), .B(n1115), .ZN(n1173) );
XNOR2_X1 U986 ( .A(n1280), .B(n1281), .ZN(n1115) );
NOR2_X1 U987 ( .A1(KEYINPUT24), .A2(n1282), .ZN(n1281) );
NAND3_X1 U988 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1279) );
NAND2_X1 U989 ( .A1(n1286), .A2(G101), .ZN(n1285) );
NAND2_X1 U990 ( .A1(KEYINPUT29), .A2(n1287), .ZN(n1284) );
NAND2_X1 U991 ( .A1(n1288), .A2(n1228), .ZN(n1287) );
XNOR2_X1 U992 ( .A(KEYINPUT12), .B(n1286), .ZN(n1288) );
NAND2_X1 U993 ( .A1(n1289), .A2(n1290), .ZN(n1283) );
INV_X1 U994 ( .A(KEYINPUT29), .ZN(n1290) );
NAND2_X1 U995 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
NAND2_X1 U996 ( .A1(KEYINPUT12), .A2(n1286), .ZN(n1292) );
OR3_X1 U997 ( .A1(G101), .A2(KEYINPUT12), .A3(n1286), .ZN(n1291) );
XOR2_X1 U998 ( .A(n1293), .B(KEYINPUT1), .Z(n1286) );
NOR2_X1 U999 ( .A1(n1052), .A2(n1054), .ZN(n1051) );
AND2_X1 U1000 ( .A1(G214), .A2(n1294), .ZN(n1054) );
INV_X1 U1001 ( .A(n1225), .ZN(n1052) );
XOR2_X1 U1002 ( .A(n1295), .B(n1181), .Z(n1225) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1294), .ZN(n1181) );
NAND2_X1 U1004 ( .A1(n1296), .A2(n1258), .ZN(n1294) );
INV_X1 U1005 ( .A(G237), .ZN(n1296) );
NAND2_X1 U1006 ( .A1(KEYINPUT10), .A2(n1297), .ZN(n1295) );
INV_X1 U1007 ( .A(n1087), .ZN(n1297) );
NAND2_X1 U1008 ( .A1(n1298), .A2(n1258), .ZN(n1087) );
XNOR2_X1 U1009 ( .A(G125), .B(n1175), .ZN(n1298) );
XNOR2_X1 U1010 ( .A(n1299), .B(n1300), .ZN(n1175) );
XNOR2_X1 U1011 ( .A(n1301), .B(n1137), .ZN(n1300) );
XOR2_X1 U1012 ( .A(n1302), .B(G110), .Z(n1137) );
NAND2_X1 U1013 ( .A1(KEYINPUT17), .A2(G122), .ZN(n1302) );
XOR2_X1 U1014 ( .A(n1303), .B(n1304), .Z(n1299) );
NOR2_X1 U1015 ( .A1(KEYINPUT36), .A2(n1305), .ZN(n1304) );
NOR2_X1 U1016 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1017 ( .A(KEYINPUT60), .B(n1308), .Z(n1307) );
AND2_X1 U1018 ( .A1(n1136), .A2(n1139), .ZN(n1308) );
NOR2_X1 U1019 ( .A1(n1139), .A2(n1136), .ZN(n1306) );
XOR2_X1 U1020 ( .A(n1293), .B(n1228), .Z(n1136) );
XNOR2_X1 U1021 ( .A(G104), .B(n1263), .ZN(n1293) );
XOR2_X1 U1022 ( .A(G107), .B(KEYINPUT47), .Z(n1263) );
XOR2_X1 U1023 ( .A(n1309), .B(n1310), .Z(n1139) );
NAND2_X1 U1024 ( .A1(G224), .A2(n1108), .ZN(n1303) );
INV_X1 U1025 ( .A(G953), .ZN(n1108) );
NOR2_X1 U1026 ( .A1(n1207), .A2(n1090), .ZN(n1070) );
INV_X1 U1027 ( .A(n1204), .ZN(n1090) );
XNOR2_X1 U1028 ( .A(n1311), .B(n1312), .ZN(n1204) );
NOR2_X1 U1029 ( .A1(n1269), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1030 ( .A(KEYINPUT34), .B(G217), .Z(n1313) );
AND2_X1 U1031 ( .A1(G234), .A2(n1258), .ZN(n1269) );
OR2_X1 U1032 ( .A1(n1144), .A2(G902), .ZN(n1311) );
XNOR2_X1 U1033 ( .A(n1314), .B(n1315), .ZN(n1144) );
NOR3_X1 U1034 ( .A1(n1316), .A2(G953), .A3(n1268), .ZN(n1315) );
INV_X1 U1035 ( .A(G221), .ZN(n1268) );
XOR2_X1 U1036 ( .A(KEYINPUT19), .B(G234), .Z(n1316) );
XOR2_X1 U1037 ( .A(n1317), .B(G137), .Z(n1314) );
NAND2_X1 U1038 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1039 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XOR2_X1 U1040 ( .A(KEYINPUT55), .B(n1322), .Z(n1318) );
NOR2_X1 U1041 ( .A1(n1323), .A2(n1321), .ZN(n1322) );
XNOR2_X1 U1042 ( .A(n1324), .B(G110), .ZN(n1321) );
NAND2_X1 U1043 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1044 ( .A1(G119), .A2(n1280), .ZN(n1326) );
INV_X1 U1045 ( .A(G128), .ZN(n1280) );
XOR2_X1 U1046 ( .A(n1327), .B(KEYINPUT5), .Z(n1325) );
NAND2_X1 U1047 ( .A1(G128), .A2(n1238), .ZN(n1327) );
XOR2_X1 U1048 ( .A(n1320), .B(KEYINPUT46), .Z(n1323) );
XNOR2_X1 U1049 ( .A(n1328), .B(n1122), .ZN(n1320) );
XNOR2_X1 U1050 ( .A(n1179), .B(n1123), .ZN(n1122) );
INV_X1 U1051 ( .A(G140), .ZN(n1123) );
INV_X1 U1052 ( .A(G125), .ZN(n1179) );
XNOR2_X1 U1053 ( .A(G146), .B(KEYINPUT51), .ZN(n1328) );
XOR2_X1 U1054 ( .A(n1096), .B(n1098), .Z(n1207) );
INV_X1 U1055 ( .A(G472), .ZN(n1098) );
NAND2_X1 U1056 ( .A1(n1258), .A2(n1329), .ZN(n1096) );
NAND2_X1 U1057 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1058 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1059 ( .A(KEYINPUT52), .B(n1156), .Z(n1333) );
XNOR2_X1 U1060 ( .A(n1334), .B(n1164), .ZN(n1332) );
XOR2_X1 U1061 ( .A(n1335), .B(KEYINPUT27), .Z(n1330) );
NAND2_X1 U1062 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1063 ( .A(n1334), .B(n1338), .ZN(n1337) );
INV_X1 U1064 ( .A(n1164), .ZN(n1338) );
XNOR2_X1 U1065 ( .A(n1309), .B(n1339), .ZN(n1164) );
NOR2_X1 U1066 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
AND3_X1 U1067 ( .A1(KEYINPUT15), .A2(n1238), .A3(G116), .ZN(n1341) );
NOR2_X1 U1068 ( .A1(KEYINPUT15), .A2(n1310), .ZN(n1340) );
XNOR2_X1 U1069 ( .A(G116), .B(n1238), .ZN(n1310) );
INV_X1 U1070 ( .A(G119), .ZN(n1238) );
XNOR2_X1 U1071 ( .A(G113), .B(KEYINPUT48), .ZN(n1309) );
NAND2_X1 U1072 ( .A1(KEYINPUT59), .A2(n1162), .ZN(n1334) );
XOR2_X1 U1073 ( .A(n1342), .B(n1343), .Z(n1162) );
INV_X1 U1074 ( .A(n1301), .ZN(n1343) );
XOR2_X1 U1075 ( .A(n1344), .B(n1282), .Z(n1301) );
XNOR2_X1 U1076 ( .A(n1267), .B(n1216), .ZN(n1282) );
INV_X1 U1077 ( .A(G146), .ZN(n1216) );
INV_X1 U1078 ( .A(G143), .ZN(n1267) );
NAND2_X1 U1079 ( .A1(KEYINPUT53), .A2(G128), .ZN(n1344) );
XNOR2_X1 U1080 ( .A(n1171), .B(KEYINPUT22), .ZN(n1342) );
INV_X1 U1081 ( .A(n1275), .ZN(n1171) );
NAND2_X1 U1082 ( .A1(n1345), .A2(n1346), .ZN(n1275) );
NAND2_X1 U1083 ( .A1(n1117), .A2(n1119), .ZN(n1346) );
XOR2_X1 U1084 ( .A(KEYINPUT54), .B(n1347), .Z(n1345) );
NOR2_X1 U1085 ( .A1(n1117), .A2(n1119), .ZN(n1347) );
XOR2_X1 U1086 ( .A(G131), .B(KEYINPUT2), .Z(n1119) );
XOR2_X1 U1087 ( .A(G134), .B(G137), .Z(n1117) );
XNOR2_X1 U1088 ( .A(n1156), .B(KEYINPUT52), .ZN(n1336) );
XOR2_X1 U1089 ( .A(n1348), .B(n1228), .Z(n1156) );
INV_X1 U1090 ( .A(G101), .ZN(n1228) );
NAND2_X1 U1091 ( .A1(n1249), .A2(G210), .ZN(n1348) );
NOR2_X1 U1092 ( .A1(G953), .A2(G237), .ZN(n1249) );
INV_X1 U1093 ( .A(G902), .ZN(n1258) );
endmodule


