//Key = 0101101001001000011011001110110000010001110110101101000011000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419;

XNOR2_X1 U784 ( .A(G107), .B(n1078), .ZN(G9) );
NAND4_X1 U785 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
XOR2_X1 U786 ( .A(KEYINPUT7), .B(KEYINPUT56), .Z(n1082) );
NOR2_X1 U787 ( .A1(n1083), .A2(n1084), .ZN(G75) );
NOR3_X1 U788 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND3_X1 U789 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1085) );
NAND2_X1 U790 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U791 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND4_X1 U792 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
NAND2_X1 U793 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
OR2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U796 ( .A1(n1081), .A2(n1105), .ZN(n1099) );
NAND2_X1 U797 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U798 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND4_X1 U799 ( .A1(n1101), .A2(n1081), .A3(n1110), .A4(n1111), .ZN(n1093) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U801 ( .A1(n1095), .A2(n1096), .ZN(n1113) );
NAND2_X1 U802 ( .A1(n1114), .A2(n1098), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
OR2_X1 U804 ( .A1(n1095), .A2(n1096), .ZN(n1116) );
OR3_X1 U805 ( .A1(n1080), .A2(n1117), .A3(n1118), .ZN(n1115) );
INV_X1 U806 ( .A(n1119), .ZN(n1091) );
AND3_X1 U807 ( .A1(n1088), .A2(n1089), .A3(n1120), .ZN(n1083) );
NAND4_X1 U808 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1088) );
NOR4_X1 U809 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1124) );
XOR2_X1 U810 ( .A(KEYINPUT0), .B(n1129), .Z(n1128) );
NOR3_X1 U811 ( .A1(n1112), .A2(n1130), .A3(n1131), .ZN(n1123) );
INV_X1 U812 ( .A(n1132), .ZN(n1131) );
NAND2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1122) );
XNOR2_X1 U814 ( .A(KEYINPUT17), .B(n1135), .ZN(n1134) );
XOR2_X1 U815 ( .A(KEYINPUT11), .B(G472), .Z(n1133) );
OR2_X1 U816 ( .A1(n1135), .A2(G472), .ZN(n1121) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(G72) );
NOR2_X1 U818 ( .A1(n1138), .A2(n1089), .ZN(n1137) );
AND2_X1 U819 ( .A1(G227), .A2(G900), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U821 ( .A1(n1141), .A2(n1089), .ZN(n1140) );
XNOR2_X1 U822 ( .A(n1086), .B(n1142), .ZN(n1141) );
OR3_X1 U823 ( .A1(n1143), .A2(n1142), .A3(n1089), .ZN(n1139) );
XNOR2_X1 U824 ( .A(n1144), .B(n1145), .ZN(n1142) );
XNOR2_X1 U825 ( .A(G131), .B(n1146), .ZN(n1145) );
XOR2_X1 U826 ( .A(n1147), .B(n1148), .Z(n1144) );
NAND2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
NAND2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U829 ( .A(KEYINPUT4), .B(n1153), .Z(n1149) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1151), .ZN(n1153) );
XOR2_X1 U831 ( .A(n1154), .B(n1155), .Z(G69) );
XOR2_X1 U832 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U833 ( .A1(n1158), .A2(n1089), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U835 ( .A1(n1161), .A2(n1162), .ZN(n1156) );
NAND2_X1 U836 ( .A1(G953), .A2(n1160), .ZN(n1162) );
XOR2_X1 U837 ( .A(n1163), .B(KEYINPUT28), .Z(n1161) );
NAND2_X1 U838 ( .A1(n1089), .A2(n1087), .ZN(n1154) );
NOR2_X1 U839 ( .A1(n1164), .A2(n1165), .ZN(G66) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U841 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NOR2_X1 U842 ( .A1(n1164), .A2(n1170), .ZN(G63) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U844 ( .A(KEYINPUT58), .B(n1173), .Z(n1172) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
AND2_X1 U846 ( .A1(n1175), .A2(n1174), .ZN(n1171) );
NAND2_X1 U847 ( .A1(n1168), .A2(G478), .ZN(n1175) );
NOR3_X1 U848 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(G60) );
AND2_X1 U849 ( .A1(KEYINPUT9), .A2(n1164), .ZN(n1178) );
NOR3_X1 U850 ( .A1(KEYINPUT9), .A2(n1120), .A3(n1089), .ZN(n1177) );
INV_X1 U851 ( .A(G952), .ZN(n1120) );
XOR2_X1 U852 ( .A(n1179), .B(n1180), .Z(n1176) );
NAND3_X1 U853 ( .A1(n1168), .A2(G475), .A3(KEYINPUT24), .ZN(n1179) );
XNOR2_X1 U854 ( .A(G104), .B(n1181), .ZN(G6) );
NOR2_X1 U855 ( .A1(n1164), .A2(n1182), .ZN(G57) );
NOR2_X1 U856 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U857 ( .A(KEYINPUT16), .B(n1185), .Z(n1184) );
NOR2_X1 U858 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U859 ( .A(G101), .B(n1188), .ZN(n1187) );
NOR2_X1 U860 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
XNOR2_X1 U861 ( .A(n1188), .B(n1191), .ZN(n1190) );
INV_X1 U862 ( .A(n1186), .ZN(n1189) );
XNOR2_X1 U863 ( .A(n1192), .B(n1193), .ZN(n1186) );
NOR2_X1 U864 ( .A1(KEYINPUT30), .A2(n1194), .ZN(n1193) );
NOR3_X1 U865 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
NOR2_X1 U866 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR3_X1 U867 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1196) );
INV_X1 U868 ( .A(n1199), .ZN(n1200) );
NAND2_X1 U869 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
XNOR2_X1 U870 ( .A(KEYINPUT2), .B(n1205), .ZN(n1203) );
INV_X1 U871 ( .A(n1206), .ZN(n1195) );
NAND2_X1 U872 ( .A1(n1168), .A2(G472), .ZN(n1192) );
NOR2_X1 U873 ( .A1(n1164), .A2(n1207), .ZN(G54) );
XOR2_X1 U874 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U875 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U876 ( .A(KEYINPUT38), .B(n1212), .ZN(n1211) );
NOR2_X1 U877 ( .A1(KEYINPUT45), .A2(n1213), .ZN(n1212) );
XNOR2_X1 U878 ( .A(n1146), .B(n1214), .ZN(n1213) );
NOR2_X1 U879 ( .A1(KEYINPUT55), .A2(n1215), .ZN(n1214) );
NAND2_X1 U880 ( .A1(n1216), .A2(n1168), .ZN(n1210) );
XNOR2_X1 U881 ( .A(G469), .B(KEYINPUT48), .ZN(n1216) );
XNOR2_X1 U882 ( .A(n1217), .B(n1218), .ZN(n1208) );
XNOR2_X1 U883 ( .A(n1219), .B(n1220), .ZN(n1217) );
NAND3_X1 U884 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1219) );
NAND2_X1 U885 ( .A1(KEYINPUT32), .A2(n1224), .ZN(n1222) );
NAND2_X1 U886 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
INV_X1 U887 ( .A(KEYINPUT32), .ZN(n1226) );
NOR2_X1 U888 ( .A1(n1164), .A2(n1227), .ZN(G51) );
NOR2_X1 U889 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XOR2_X1 U890 ( .A(n1230), .B(KEYINPUT20), .Z(n1229) );
NAND2_X1 U891 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(n1228) );
AND2_X1 U893 ( .A1(n1168), .A2(n1233), .ZN(n1231) );
AND2_X1 U894 ( .A1(G902), .A2(n1234), .ZN(n1168) );
OR2_X1 U895 ( .A1(n1087), .A2(n1086), .ZN(n1234) );
NAND4_X1 U896 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1086) );
AND4_X1 U897 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1238) );
NOR2_X1 U898 ( .A1(n1243), .A2(n1244), .ZN(n1237) );
NOR2_X1 U899 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
INV_X1 U900 ( .A(KEYINPUT41), .ZN(n1246) );
NOR3_X1 U901 ( .A1(n1247), .A2(n1248), .A3(n1106), .ZN(n1243) );
NOR2_X1 U902 ( .A1(n1249), .A2(n1080), .ZN(n1248) );
NOR2_X1 U903 ( .A1(KEYINPUT41), .A2(n1117), .ZN(n1249) );
NAND4_X1 U904 ( .A1(n1250), .A2(n1117), .A3(n1103), .A4(n1101), .ZN(n1235) );
NAND4_X1 U905 ( .A1(n1181), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1087) );
NOR4_X1 U906 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1253) );
INV_X1 U907 ( .A(n1258), .ZN(n1257) );
NAND2_X1 U908 ( .A1(n1081), .A2(n1259), .ZN(n1252) );
NAND2_X1 U909 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U910 ( .A1(n1129), .A2(n1126), .A3(n1262), .ZN(n1261) );
NAND3_X1 U911 ( .A1(n1263), .A2(n1264), .A3(n1080), .ZN(n1260) );
OR2_X1 U912 ( .A1(n1079), .A2(KEYINPUT63), .ZN(n1264) );
NAND2_X1 U913 ( .A1(KEYINPUT63), .A2(n1265), .ZN(n1263) );
NAND3_X1 U914 ( .A1(n1266), .A2(n1118), .A3(n1267), .ZN(n1265) );
NAND3_X1 U915 ( .A1(n1079), .A2(n1081), .A3(n1117), .ZN(n1181) );
NOR2_X1 U916 ( .A1(n1089), .A2(G952), .ZN(n1164) );
NAND2_X1 U917 ( .A1(n1268), .A2(n1269), .ZN(G48) );
NAND2_X1 U918 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U919 ( .A(n1245), .B(KEYINPUT46), .Z(n1270) );
NAND2_X1 U920 ( .A1(n1272), .A2(G146), .ZN(n1268) );
XOR2_X1 U921 ( .A(n1245), .B(KEYINPUT13), .Z(n1272) );
NAND3_X1 U922 ( .A1(n1117), .A2(n1273), .A3(n1274), .ZN(n1245) );
NAND2_X1 U923 ( .A1(n1275), .A2(n1276), .ZN(G45) );
NAND2_X1 U924 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U925 ( .A(KEYINPUT21), .B(n1279), .Z(n1275) );
NOR2_X1 U926 ( .A1(n1277), .A2(n1278), .ZN(n1279) );
INV_X1 U927 ( .A(n1236), .ZN(n1277) );
NAND4_X1 U928 ( .A1(n1280), .A2(n1273), .A3(n1129), .A4(n1126), .ZN(n1236) );
XOR2_X1 U929 ( .A(n1281), .B(n1282), .Z(G42) );
NAND2_X1 U930 ( .A1(KEYINPUT26), .A2(G140), .ZN(n1282) );
NAND4_X1 U931 ( .A1(n1283), .A2(n1250), .A3(n1117), .A4(n1284), .ZN(n1281) );
XNOR2_X1 U932 ( .A(KEYINPUT59), .B(n1127), .ZN(n1284) );
XNOR2_X1 U933 ( .A(n1103), .B(KEYINPUT35), .ZN(n1283) );
XNOR2_X1 U934 ( .A(G137), .B(n1242), .ZN(G39) );
NAND3_X1 U935 ( .A1(n1096), .A2(n1101), .A3(n1274), .ZN(n1242) );
XOR2_X1 U936 ( .A(n1241), .B(n1285), .Z(G36) );
XNOR2_X1 U937 ( .A(G134), .B(KEYINPUT60), .ZN(n1285) );
NAND3_X1 U938 ( .A1(n1101), .A2(n1080), .A3(n1280), .ZN(n1241) );
XNOR2_X1 U939 ( .A(G131), .B(n1240), .ZN(G33) );
NAND3_X1 U940 ( .A1(n1117), .A2(n1101), .A3(n1280), .ZN(n1240) );
AND2_X1 U941 ( .A1(n1250), .A2(n1104), .ZN(n1280) );
INV_X1 U942 ( .A(n1127), .ZN(n1101) );
NAND2_X1 U943 ( .A1(n1109), .A2(n1286), .ZN(n1127) );
XOR2_X1 U944 ( .A(n1287), .B(n1288), .Z(G30) );
NAND2_X1 U945 ( .A1(KEYINPUT62), .A2(G128), .ZN(n1288) );
NAND2_X1 U946 ( .A1(n1289), .A2(n1273), .ZN(n1287) );
XOR2_X1 U947 ( .A(n1290), .B(KEYINPUT18), .Z(n1289) );
NAND2_X1 U948 ( .A1(n1274), .A2(n1080), .ZN(n1290) );
INV_X1 U949 ( .A(n1247), .ZN(n1274) );
NAND3_X1 U950 ( .A1(n1291), .A2(n1125), .A3(n1250), .ZN(n1247) );
NOR3_X1 U951 ( .A1(n1095), .A2(n1292), .A3(n1112), .ZN(n1250) );
XNOR2_X1 U952 ( .A(G101), .B(n1258), .ZN(G3) );
NAND3_X1 U953 ( .A1(n1096), .A2(n1079), .A3(n1104), .ZN(n1258) );
XNOR2_X1 U954 ( .A(G125), .B(n1239), .ZN(G27) );
NAND4_X1 U955 ( .A1(n1117), .A2(n1095), .A3(n1293), .A4(n1103), .ZN(n1239) );
NOR2_X1 U956 ( .A1(n1292), .A2(n1294), .ZN(n1293) );
AND2_X1 U957 ( .A1(n1295), .A2(n1119), .ZN(n1292) );
NAND2_X1 U958 ( .A1(n1296), .A2(n1143), .ZN(n1295) );
INV_X1 U959 ( .A(G900), .ZN(n1143) );
XNOR2_X1 U960 ( .A(G122), .B(n1297), .ZN(G24) );
NAND3_X1 U961 ( .A1(KEYINPUT51), .A2(n1262), .A3(n1298), .ZN(n1297) );
AND3_X1 U962 ( .A1(n1081), .A2(n1126), .A3(n1129), .ZN(n1298) );
NOR2_X1 U963 ( .A1(n1125), .A2(n1291), .ZN(n1081) );
XNOR2_X1 U964 ( .A(G119), .B(n1251), .ZN(G21) );
NAND4_X1 U965 ( .A1(n1262), .A2(n1096), .A3(n1291), .A4(n1125), .ZN(n1251) );
XOR2_X1 U966 ( .A(G116), .B(n1256), .Z(G18) );
AND3_X1 U967 ( .A1(n1104), .A2(n1080), .A3(n1262), .ZN(n1256) );
AND2_X1 U968 ( .A1(n1299), .A2(n1129), .ZN(n1080) );
XOR2_X1 U969 ( .A(n1255), .B(n1300), .Z(G15) );
NOR2_X1 U970 ( .A1(KEYINPUT42), .A2(n1301), .ZN(n1300) );
INV_X1 U971 ( .A(G113), .ZN(n1301) );
AND3_X1 U972 ( .A1(n1117), .A2(n1104), .A3(n1262), .ZN(n1255) );
NOR3_X1 U973 ( .A1(n1294), .A2(n1267), .A3(n1118), .ZN(n1262) );
AND2_X1 U974 ( .A1(n1302), .A2(n1291), .ZN(n1104) );
NOR2_X1 U975 ( .A1(n1129), .A2(n1299), .ZN(n1117) );
INV_X1 U976 ( .A(n1126), .ZN(n1299) );
XNOR2_X1 U977 ( .A(G110), .B(n1303), .ZN(G12) );
NOR2_X1 U978 ( .A1(n1254), .A2(KEYINPUT10), .ZN(n1303) );
AND3_X1 U979 ( .A1(n1103), .A2(n1079), .A3(n1096), .ZN(n1254) );
NOR2_X1 U980 ( .A1(n1129), .A2(n1126), .ZN(n1096) );
XNOR2_X1 U981 ( .A(n1304), .B(G475), .ZN(n1126) );
NAND2_X1 U982 ( .A1(n1180), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U983 ( .A(n1306), .B(n1307), .ZN(n1180) );
XNOR2_X1 U984 ( .A(n1308), .B(n1309), .ZN(n1307) );
NAND2_X1 U985 ( .A1(KEYINPUT3), .A2(n1310), .ZN(n1308) );
INV_X1 U986 ( .A(G104), .ZN(n1310) );
XOR2_X1 U987 ( .A(n1311), .B(n1312), .Z(n1306) );
XNOR2_X1 U988 ( .A(G131), .B(n1313), .ZN(n1312) );
NAND2_X1 U989 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
OR2_X1 U990 ( .A1(n1316), .A2(G146), .ZN(n1315) );
XOR2_X1 U991 ( .A(n1317), .B(KEYINPUT14), .Z(n1314) );
NAND2_X1 U992 ( .A1(G146), .A2(n1316), .ZN(n1317) );
XOR2_X1 U993 ( .A(n1148), .B(KEYINPUT31), .Z(n1316) );
XNOR2_X1 U994 ( .A(G125), .B(n1224), .ZN(n1148) );
NAND2_X1 U995 ( .A1(n1318), .A2(KEYINPUT57), .ZN(n1311) );
XNOR2_X1 U996 ( .A(n1319), .B(n1278), .ZN(n1318) );
NAND2_X1 U997 ( .A1(n1320), .A2(G214), .ZN(n1319) );
XNOR2_X1 U998 ( .A(n1321), .B(G478), .ZN(n1129) );
NAND2_X1 U999 ( .A1(n1174), .A2(n1305), .ZN(n1321) );
XOR2_X1 U1000 ( .A(n1322), .B(n1323), .Z(n1174) );
XOR2_X1 U1001 ( .A(n1324), .B(n1325), .Z(n1323) );
AND3_X1 U1002 ( .A1(G217), .A2(n1089), .A3(G234), .ZN(n1325) );
NOR2_X1 U1003 ( .A1(KEYINPUT54), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1004 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1005 ( .A(n1329), .B(G107), .ZN(n1328) );
NOR2_X1 U1006 ( .A1(G116), .A2(KEYINPUT37), .ZN(n1327) );
NAND3_X1 U1007 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1322) );
NAND2_X1 U1008 ( .A1(KEYINPUT33), .A2(n1333), .ZN(n1332) );
NAND3_X1 U1009 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1331) );
INV_X1 U1010 ( .A(KEYINPUT33), .ZN(n1335) );
OR2_X1 U1011 ( .A1(n1336), .A2(n1334), .ZN(n1330) );
NOR2_X1 U1012 ( .A1(n1333), .A2(KEYINPUT50), .ZN(n1334) );
AND2_X1 U1013 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
NAND2_X1 U1014 ( .A1(G143), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1015 ( .A(n1340), .B(KEYINPUT8), .Z(n1337) );
NAND2_X1 U1016 ( .A1(G128), .A2(n1278), .ZN(n1340) );
INV_X1 U1017 ( .A(G143), .ZN(n1278) );
NOR3_X1 U1018 ( .A1(n1095), .A2(n1267), .A3(n1294), .ZN(n1079) );
INV_X1 U1019 ( .A(n1266), .ZN(n1294) );
NOR2_X1 U1020 ( .A1(n1106), .A2(n1112), .ZN(n1266) );
INV_X1 U1021 ( .A(n1098), .ZN(n1112) );
NAND2_X1 U1022 ( .A1(G221), .A2(n1341), .ZN(n1098) );
INV_X1 U1023 ( .A(n1273), .ZN(n1106) );
NOR2_X1 U1024 ( .A1(n1109), .A2(n1108), .ZN(n1273) );
INV_X1 U1025 ( .A(n1286), .ZN(n1108) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1342), .ZN(n1286) );
XOR2_X1 U1027 ( .A(n1343), .B(n1233), .Z(n1109) );
AND2_X1 U1028 ( .A1(G210), .A2(n1342), .ZN(n1233) );
NAND2_X1 U1029 ( .A1(n1344), .A2(n1305), .ZN(n1342) );
INV_X1 U1030 ( .A(G237), .ZN(n1344) );
NAND2_X1 U1031 ( .A1(n1345), .A2(n1305), .ZN(n1343) );
XOR2_X1 U1032 ( .A(KEYINPUT44), .B(n1232), .Z(n1345) );
XNOR2_X1 U1033 ( .A(n1346), .B(n1347), .ZN(n1232) );
XNOR2_X1 U1034 ( .A(n1348), .B(n1349), .ZN(n1347) );
NOR2_X1 U1035 ( .A1(G953), .A2(n1159), .ZN(n1349) );
INV_X1 U1036 ( .A(G224), .ZN(n1159) );
XNOR2_X1 U1037 ( .A(n1163), .B(n1205), .ZN(n1346) );
XOR2_X1 U1038 ( .A(n1350), .B(n1351), .Z(n1163) );
XOR2_X1 U1039 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1040 ( .A(G116), .B(G110), .Z(n1353) );
XNOR2_X1 U1041 ( .A(KEYINPUT12), .B(n1354), .ZN(n1352) );
XOR2_X1 U1042 ( .A(n1355), .B(n1356), .Z(n1350) );
XNOR2_X1 U1043 ( .A(n1357), .B(G104), .ZN(n1356) );
XNOR2_X1 U1044 ( .A(G101), .B(n1309), .ZN(n1355) );
XNOR2_X1 U1045 ( .A(G113), .B(n1329), .ZN(n1309) );
INV_X1 U1046 ( .A(G122), .ZN(n1329) );
AND2_X1 U1047 ( .A1(n1358), .A2(n1119), .ZN(n1267) );
NAND3_X1 U1048 ( .A1(n1359), .A2(n1089), .A3(G952), .ZN(n1119) );
NAND2_X1 U1049 ( .A1(n1296), .A2(n1160), .ZN(n1358) );
INV_X1 U1050 ( .A(G898), .ZN(n1160) );
AND3_X1 U1051 ( .A1(G902), .A2(n1359), .A3(G953), .ZN(n1296) );
NAND2_X1 U1052 ( .A1(G237), .A2(G234), .ZN(n1359) );
INV_X1 U1053 ( .A(n1118), .ZN(n1095) );
NAND2_X1 U1054 ( .A1(n1360), .A2(n1132), .ZN(n1118) );
NAND2_X1 U1055 ( .A1(G469), .A2(n1361), .ZN(n1132) );
OR2_X1 U1056 ( .A1(n1362), .A2(G902), .ZN(n1361) );
XOR2_X1 U1057 ( .A(KEYINPUT49), .B(n1130), .Z(n1360) );
NOR3_X1 U1058 ( .A1(G469), .A2(G902), .A3(n1362), .ZN(n1130) );
XNOR2_X1 U1059 ( .A(n1363), .B(n1364), .ZN(n1362) );
NOR2_X1 U1060 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1061 ( .A(KEYINPUT52), .B(n1367), .Z(n1366) );
NOR3_X1 U1062 ( .A1(n1220), .A2(n1225), .A3(n1368), .ZN(n1367) );
NOR2_X1 U1063 ( .A1(n1369), .A2(n1370), .ZN(n1365) );
INV_X1 U1064 ( .A(n1220), .ZN(n1370) );
NAND2_X1 U1065 ( .A1(G227), .A2(n1089), .ZN(n1220) );
NOR2_X1 U1066 ( .A1(n1225), .A2(n1368), .ZN(n1369) );
INV_X1 U1067 ( .A(n1223), .ZN(n1368) );
NAND2_X1 U1068 ( .A1(G110), .A2(n1224), .ZN(n1223) );
NOR2_X1 U1069 ( .A1(n1224), .A2(G110), .ZN(n1225) );
INV_X1 U1070 ( .A(G140), .ZN(n1224) );
NAND3_X1 U1071 ( .A1(n1371), .A2(n1372), .A3(n1373), .ZN(n1363) );
OR2_X1 U1072 ( .A1(n1374), .A2(KEYINPUT25), .ZN(n1373) );
NAND3_X1 U1073 ( .A1(KEYINPUT25), .A2(n1374), .A3(n1204), .ZN(n1372) );
NAND2_X1 U1074 ( .A1(n1218), .A2(n1375), .ZN(n1371) );
NAND2_X1 U1075 ( .A1(KEYINPUT25), .A2(n1376), .ZN(n1375) );
XNOR2_X1 U1076 ( .A(KEYINPUT29), .B(n1374), .ZN(n1376) );
XOR2_X1 U1077 ( .A(n1146), .B(n1215), .Z(n1374) );
XNOR2_X1 U1078 ( .A(n1377), .B(n1378), .ZN(n1215) );
XNOR2_X1 U1079 ( .A(KEYINPUT36), .B(n1191), .ZN(n1378) );
NAND3_X1 U1080 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1377) );
NAND2_X1 U1081 ( .A1(KEYINPUT22), .A2(G104), .ZN(n1381) );
NAND3_X1 U1082 ( .A1(n1382), .A2(n1383), .A3(n1357), .ZN(n1380) );
INV_X1 U1083 ( .A(KEYINPUT22), .ZN(n1383) );
OR2_X1 U1084 ( .A1(n1357), .A2(n1382), .ZN(n1379) );
NOR2_X1 U1085 ( .A1(G104), .A2(KEYINPUT27), .ZN(n1382) );
INV_X1 U1086 ( .A(G107), .ZN(n1357) );
NAND3_X1 U1087 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n1146) );
NAND2_X1 U1088 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
INV_X1 U1089 ( .A(KEYINPUT43), .ZN(n1388) );
NAND3_X1 U1090 ( .A1(KEYINPUT43), .A2(n1389), .A3(n1339), .ZN(n1385) );
OR2_X1 U1091 ( .A1(n1339), .A2(n1389), .ZN(n1384) );
NOR2_X1 U1092 ( .A1(n1390), .A2(n1387), .ZN(n1389) );
XOR2_X1 U1093 ( .A(G143), .B(n1391), .Z(n1387) );
XNOR2_X1 U1094 ( .A(KEYINPUT39), .B(n1271), .ZN(n1391) );
INV_X1 U1095 ( .A(KEYINPUT6), .ZN(n1390) );
INV_X1 U1096 ( .A(G128), .ZN(n1339) );
INV_X1 U1097 ( .A(n1204), .ZN(n1218) );
NOR2_X1 U1098 ( .A1(n1291), .A2(n1302), .ZN(n1103) );
INV_X1 U1099 ( .A(n1125), .ZN(n1302) );
XNOR2_X1 U1100 ( .A(n1392), .B(n1169), .ZN(n1125) );
AND2_X1 U1101 ( .A1(G217), .A2(n1341), .ZN(n1169) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1305), .ZN(n1341) );
NAND2_X1 U1103 ( .A1(n1167), .A2(n1305), .ZN(n1392) );
XNOR2_X1 U1104 ( .A(n1393), .B(n1394), .ZN(n1167) );
XOR2_X1 U1105 ( .A(n1395), .B(n1396), .Z(n1394) );
XOR2_X1 U1106 ( .A(n1397), .B(n1398), .Z(n1396) );
AND3_X1 U1107 ( .A1(G221), .A2(n1089), .A3(G234), .ZN(n1398) );
INV_X1 U1108 ( .A(G953), .ZN(n1089) );
NAND2_X1 U1109 ( .A1(KEYINPUT40), .A2(n1348), .ZN(n1397) );
INV_X1 U1110 ( .A(G125), .ZN(n1348) );
XOR2_X1 U1111 ( .A(n1399), .B(G110), .Z(n1395) );
NAND2_X1 U1112 ( .A1(KEYINPUT1), .A2(n1354), .ZN(n1399) );
INV_X1 U1113 ( .A(G119), .ZN(n1354) );
XOR2_X1 U1114 ( .A(n1400), .B(n1401), .Z(n1393) );
XNOR2_X1 U1115 ( .A(n1271), .B(G140), .ZN(n1401) );
XNOR2_X1 U1116 ( .A(G137), .B(G128), .ZN(n1400) );
XNOR2_X1 U1117 ( .A(n1135), .B(G472), .ZN(n1291) );
NAND2_X1 U1118 ( .A1(n1402), .A2(n1305), .ZN(n1135) );
INV_X1 U1119 ( .A(G902), .ZN(n1305) );
XOR2_X1 U1120 ( .A(n1403), .B(n1404), .Z(n1402) );
NAND2_X1 U1121 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
OR2_X1 U1122 ( .A1(n1188), .A2(n1191), .ZN(n1406) );
XOR2_X1 U1123 ( .A(n1407), .B(KEYINPUT34), .Z(n1405) );
NAND2_X1 U1124 ( .A1(n1191), .A2(n1188), .ZN(n1407) );
NAND2_X1 U1125 ( .A1(n1320), .A2(n1408), .ZN(n1188) );
XOR2_X1 U1126 ( .A(KEYINPUT5), .B(G210), .Z(n1408) );
NOR2_X1 U1127 ( .A1(G953), .A2(G237), .ZN(n1320) );
INV_X1 U1128 ( .A(G101), .ZN(n1191) );
NAND3_X1 U1129 ( .A1(n1409), .A2(n1410), .A3(n1206), .ZN(n1403) );
NAND2_X1 U1130 ( .A1(n1201), .A2(n1202), .ZN(n1206) );
NOR2_X1 U1131 ( .A1(n1204), .A2(n1411), .ZN(n1201) );
NAND2_X1 U1132 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
XNOR2_X1 U1133 ( .A(n1202), .B(n1204), .ZN(n1412) );
NAND3_X1 U1134 ( .A1(n1204), .A2(n1198), .A3(n1205), .ZN(n1409) );
INV_X1 U1135 ( .A(n1411), .ZN(n1205) );
XOR2_X1 U1136 ( .A(G128), .B(n1413), .Z(n1411) );
NOR2_X1 U1137 ( .A1(KEYINPUT19), .A2(n1414), .ZN(n1413) );
XNOR2_X1 U1138 ( .A(G143), .B(n1415), .ZN(n1414) );
NOR2_X1 U1139 ( .A1(KEYINPUT47), .A2(n1271), .ZN(n1415) );
INV_X1 U1140 ( .A(G146), .ZN(n1271) );
INV_X1 U1141 ( .A(n1202), .ZN(n1198) );
XNOR2_X1 U1142 ( .A(n1416), .B(n1417), .ZN(n1202) );
NOR2_X1 U1143 ( .A1(KEYINPUT23), .A2(G116), .ZN(n1417) );
XNOR2_X1 U1144 ( .A(G113), .B(G119), .ZN(n1416) );
XNOR2_X1 U1145 ( .A(n1418), .B(n1419), .ZN(n1204) );
XNOR2_X1 U1146 ( .A(n1152), .B(G131), .ZN(n1419) );
INV_X1 U1147 ( .A(G137), .ZN(n1152) );
NAND2_X1 U1148 ( .A1(KEYINPUT61), .A2(n1151), .ZN(n1418) );
XNOR2_X1 U1149 ( .A(n1336), .B(KEYINPUT53), .ZN(n1151) );
XNOR2_X1 U1150 ( .A(G134), .B(KEYINPUT15), .ZN(n1336) );
endmodule


