//Key = 1110111000110000011101111001100011000110110100011000001111111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333;

XNOR2_X1 U732 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U733 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR3_X1 U734 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR4_X1 U735 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1022) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR3_X1 U738 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1028) );
NOR3_X1 U739 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1033) );
NAND3_X1 U741 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1021) );
NAND4_X1 U742 ( .A1(n1043), .A2(n1044), .A3(n1038), .A4(n1045), .ZN(n1042) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1032), .ZN(n1045) );
NAND2_X1 U744 ( .A1(n1046), .A2(n1027), .ZN(n1044) );
OR3_X1 U745 ( .A1(n1025), .A2(KEYINPUT28), .A3(n1047), .ZN(n1046) );
INV_X1 U746 ( .A(n1048), .ZN(n1025) );
NAND3_X1 U747 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1043) );
INV_X1 U748 ( .A(n1027), .ZN(n1051) );
NAND2_X1 U749 ( .A1(n1048), .A2(n1052), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U751 ( .A1(KEYINPUT28), .A2(n1055), .ZN(n1054) );
NAND2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1049) );
NAND3_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
OR2_X1 U754 ( .A1(n1061), .A2(KEYINPUT6), .ZN(n1059) );
NAND3_X1 U755 ( .A1(n1062), .A2(n1061), .A3(KEYINPUT6), .ZN(n1058) );
NOR3_X1 U756 ( .A1(n1063), .A2(G953), .A3(G952), .ZN(n1019) );
INV_X1 U757 ( .A(n1040), .ZN(n1063) );
NAND4_X1 U758 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1040) );
NOR4_X1 U759 ( .A1(n1035), .A2(n1062), .A3(n1068), .A4(n1069), .ZN(n1067) );
NOR2_X1 U760 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
XNOR2_X1 U761 ( .A(n1072), .B(n1073), .ZN(n1071) );
NOR2_X1 U762 ( .A1(KEYINPUT31), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U763 ( .A(n1075), .B(G478), .ZN(n1065) );
XNOR2_X1 U764 ( .A(G469), .B(n1076), .ZN(n1064) );
XOR2_X1 U765 ( .A(n1077), .B(n1078), .Z(G72) );
XOR2_X1 U766 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U767 ( .A1(n1041), .A2(n1081), .ZN(n1080) );
NAND3_X1 U768 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR3_X1 U769 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
INV_X1 U770 ( .A(n1088), .ZN(n1085) );
XOR2_X1 U771 ( .A(KEYINPUT60), .B(n1089), .Z(n1083) );
NAND2_X1 U772 ( .A1(n1090), .A2(n1091), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U774 ( .A(n1094), .B(n1095), .Z(n1090) );
XNOR2_X1 U775 ( .A(n1096), .B(n1097), .ZN(n1095) );
XNOR2_X1 U776 ( .A(n1098), .B(n1099), .ZN(n1094) );
NOR2_X1 U777 ( .A1(KEYINPUT7), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U778 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND2_X1 U779 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U780 ( .A1(G134), .A2(n1105), .ZN(n1104) );
XOR2_X1 U781 ( .A(KEYINPUT11), .B(n1106), .Z(n1103) );
NOR2_X1 U782 ( .A1(G134), .A2(n1105), .ZN(n1106) );
NOR2_X1 U783 ( .A1(n1107), .A2(n1108), .ZN(n1077) );
NOR2_X1 U784 ( .A1(n1109), .A2(n1093), .ZN(n1107) );
XOR2_X1 U785 ( .A(n1110), .B(n1111), .Z(G69) );
XOR2_X1 U786 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U787 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U788 ( .A(n1116), .B(KEYINPUT23), .Z(n1115) );
AND2_X1 U789 ( .A1(n1117), .A2(n1092), .ZN(n1114) );
NOR2_X1 U790 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
XNOR2_X1 U791 ( .A(G953), .B(KEYINPUT41), .ZN(n1119) );
NOR3_X1 U792 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1118) );
XNOR2_X1 U793 ( .A(n1123), .B(KEYINPUT5), .ZN(n1122) );
NOR2_X1 U794 ( .A1(n1124), .A2(n1108), .ZN(n1110) );
XNOR2_X1 U795 ( .A(n1041), .B(KEYINPUT4), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1125), .A2(n1117), .ZN(n1124) );
NOR2_X1 U797 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XNOR2_X1 U798 ( .A(n1128), .B(n1129), .ZN(n1127) );
NOR2_X1 U799 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U800 ( .A1(n1126), .A2(n1132), .ZN(G63) );
NOR3_X1 U801 ( .A1(n1075), .A2(n1133), .A3(n1134), .ZN(n1132) );
AND3_X1 U802 ( .A1(n1135), .A2(G478), .A3(n1136), .ZN(n1134) );
NOR2_X1 U803 ( .A1(n1137), .A2(n1135), .ZN(n1133) );
AND2_X1 U804 ( .A1(n1023), .A2(G478), .ZN(n1137) );
NOR2_X1 U805 ( .A1(n1126), .A2(n1138), .ZN(G60) );
XOR2_X1 U806 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U807 ( .A1(n1141), .A2(KEYINPUT26), .ZN(n1140) );
AND2_X1 U808 ( .A1(G475), .A2(n1136), .ZN(n1141) );
XNOR2_X1 U809 ( .A(G104), .B(n1142), .ZN(G6) );
NAND2_X1 U810 ( .A1(KEYINPUT1), .A2(n1123), .ZN(n1142) );
NOR2_X1 U811 ( .A1(n1126), .A2(n1143), .ZN(G57) );
XOR2_X1 U812 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U813 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U814 ( .A1(KEYINPUT35), .A2(n1148), .ZN(n1147) );
XOR2_X1 U815 ( .A(G101), .B(n1149), .Z(n1148) );
NAND3_X1 U816 ( .A1(n1136), .A2(G472), .A3(KEYINPUT57), .ZN(n1146) );
NAND2_X1 U817 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
OR3_X1 U818 ( .A1(n1152), .A2(n1153), .A3(KEYINPUT0), .ZN(n1151) );
NAND2_X1 U819 ( .A1(n1154), .A2(KEYINPUT0), .ZN(n1150) );
NOR2_X1 U820 ( .A1(n1126), .A2(n1155), .ZN(G54) );
NOR2_X1 U821 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U822 ( .A(KEYINPUT44), .B(n1158), .Z(n1157) );
NOR2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND2_X1 U824 ( .A1(n1160), .A2(n1159), .ZN(n1156) );
XNOR2_X1 U825 ( .A(n1161), .B(n1162), .ZN(n1159) );
NAND2_X1 U826 ( .A1(KEYINPUT22), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U827 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U828 ( .A1(KEYINPUT14), .A2(n1166), .ZN(n1164) );
NAND2_X1 U829 ( .A1(n1136), .A2(G469), .ZN(n1160) );
INV_X1 U830 ( .A(n1131), .ZN(n1136) );
NOR2_X1 U831 ( .A1(n1126), .A2(n1167), .ZN(G51) );
XOR2_X1 U832 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U833 ( .A(KEYINPUT62), .B(n1170), .Z(n1169) );
NOR2_X1 U834 ( .A1(n1072), .A2(n1131), .ZN(n1170) );
NAND2_X1 U835 ( .A1(G902), .A2(n1023), .ZN(n1131) );
NAND4_X1 U836 ( .A1(n1171), .A2(n1088), .A3(n1172), .A4(n1173), .ZN(n1023) );
NOR4_X1 U837 ( .A1(n1089), .A2(n1123), .A3(n1086), .A4(n1087), .ZN(n1173) );
NOR3_X1 U838 ( .A1(n1174), .A2(n1031), .A3(n1047), .ZN(n1123) );
NOR2_X1 U839 ( .A1(n1120), .A2(n1175), .ZN(n1172) );
XOR2_X1 U840 ( .A(KEYINPUT42), .B(n1121), .Z(n1175) );
NAND4_X1 U841 ( .A1(n1176), .A2(n1018), .A3(n1177), .A4(n1178), .ZN(n1120) );
NOR3_X1 U842 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
NOR3_X1 U843 ( .A1(n1026), .A2(n1174), .A3(n1182), .ZN(n1181) );
NOR2_X1 U844 ( .A1(n1183), .A2(n1030), .ZN(n1179) );
XOR2_X1 U845 ( .A(n1184), .B(KEYINPUT50), .Z(n1183) );
OR3_X1 U846 ( .A1(n1174), .A2(n1031), .A3(n1053), .ZN(n1018) );
NAND3_X1 U847 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1088) );
XOR2_X1 U848 ( .A(KEYINPUT9), .B(n1082), .Z(n1171) );
AND4_X1 U849 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1082) );
NAND3_X1 U850 ( .A1(n1055), .A2(n1037), .A3(n1192), .ZN(n1188) );
NAND2_X1 U851 ( .A1(n1193), .A2(n1194), .ZN(n1168) );
NAND3_X1 U852 ( .A1(n1195), .A2(n1116), .A3(n1196), .ZN(n1194) );
INV_X1 U853 ( .A(KEYINPUT56), .ZN(n1196) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1116) );
XNOR2_X1 U855 ( .A(n1199), .B(n1200), .ZN(n1195) );
NAND2_X1 U856 ( .A1(n1201), .A2(KEYINPUT56), .ZN(n1193) );
NOR2_X1 U857 ( .A1(n1041), .A2(G952), .ZN(n1126) );
XNOR2_X1 U858 ( .A(n1202), .B(n1087), .ZN(G48) );
AND2_X1 U859 ( .A1(n1203), .A2(n1055), .ZN(n1087) );
XOR2_X1 U860 ( .A(n1204), .B(n1205), .Z(G45) );
NOR2_X1 U861 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1205) );
NAND3_X1 U862 ( .A1(n1187), .A2(n1185), .A3(n1206), .ZN(n1204) );
XOR2_X1 U863 ( .A(n1186), .B(KEYINPUT51), .Z(n1206) );
AND3_X1 U864 ( .A1(n1207), .A2(n1069), .A3(n1037), .ZN(n1187) );
XOR2_X1 U865 ( .A(G140), .B(n1089), .Z(G42) );
NOR3_X1 U866 ( .A1(n1182), .A2(n1047), .A3(n1208), .ZN(n1089) );
XNOR2_X1 U867 ( .A(n1105), .B(n1086), .ZN(G39) );
AND3_X1 U868 ( .A1(n1192), .A2(n1209), .A3(n1056), .ZN(n1086) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(G36) );
NAND2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
NAND2_X1 U872 ( .A1(n1189), .A2(n1216), .ZN(n1215) );
INV_X1 U873 ( .A(n1217), .ZN(n1189) );
OR2_X1 U874 ( .A1(n1216), .A2(n1218), .ZN(n1214) );
INV_X1 U875 ( .A(KEYINPUT58), .ZN(n1216) );
NAND2_X1 U876 ( .A1(n1218), .A2(G134), .ZN(n1210) );
NOR2_X1 U877 ( .A1(n1217), .A2(KEYINPUT20), .ZN(n1218) );
NOR3_X1 U878 ( .A1(n1053), .A2(n1219), .A3(n1208), .ZN(n1217) );
XNOR2_X1 U879 ( .A(n1102), .B(n1220), .ZN(G33) );
NOR3_X1 U880 ( .A1(n1221), .A2(n1219), .A3(n1208), .ZN(n1220) );
INV_X1 U881 ( .A(n1192), .ZN(n1208) );
NOR4_X1 U882 ( .A1(n1060), .A2(n1032), .A3(n1222), .A4(n1035), .ZN(n1192) );
INV_X1 U883 ( .A(n1039), .ZN(n1035) );
INV_X1 U884 ( .A(n1186), .ZN(n1222) );
XNOR2_X1 U885 ( .A(KEYINPUT32), .B(n1047), .ZN(n1221) );
XNOR2_X1 U886 ( .A(n1223), .B(n1190), .ZN(G30) );
NAND2_X1 U887 ( .A1(n1203), .A2(n1224), .ZN(n1190) );
AND3_X1 U888 ( .A1(n1209), .A2(n1186), .A3(n1185), .ZN(n1203) );
XNOR2_X1 U889 ( .A(G128), .B(KEYINPUT55), .ZN(n1223) );
XOR2_X1 U890 ( .A(G101), .B(n1180), .Z(G3) );
NOR3_X1 U891 ( .A1(n1174), .A2(n1219), .A3(n1026), .ZN(n1180) );
INV_X1 U892 ( .A(n1037), .ZN(n1219) );
XNOR2_X1 U893 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U894 ( .A1(n1048), .A2(n1186), .A3(n1225), .A4(n1226), .ZN(n1191) );
NOR2_X1 U895 ( .A1(n1047), .A2(n1182), .ZN(n1226) );
NAND2_X1 U896 ( .A1(n1027), .A2(n1227), .ZN(n1186) );
NAND4_X1 U897 ( .A1(n1092), .A2(G902), .A3(n1228), .A4(n1093), .ZN(n1227) );
INV_X1 U898 ( .A(G900), .ZN(n1093) );
XOR2_X1 U899 ( .A(G122), .B(n1121), .Z(G24) );
AND4_X1 U900 ( .A1(n1229), .A2(n1038), .A3(n1207), .A4(n1069), .ZN(n1121) );
XOR2_X1 U901 ( .A(G119), .B(n1230), .Z(G21) );
NOR2_X1 U902 ( .A1(n1184), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U903 ( .A(KEYINPUT37), .B(n1030), .ZN(n1231) );
NAND4_X1 U904 ( .A1(n1056), .A2(n1209), .A3(n1048), .A4(n1232), .ZN(n1184) );
NAND2_X1 U905 ( .A1(n1233), .A2(n1234), .ZN(n1209) );
NAND2_X1 U906 ( .A1(n1036), .A2(n1235), .ZN(n1234) );
INV_X1 U907 ( .A(n1182), .ZN(n1036) );
NAND3_X1 U908 ( .A1(n1236), .A2(n1070), .A3(KEYINPUT21), .ZN(n1233) );
INV_X1 U909 ( .A(n1026), .ZN(n1056) );
XOR2_X1 U910 ( .A(n1237), .B(G116), .Z(G18) );
NAND2_X1 U911 ( .A1(KEYINPUT38), .A2(n1177), .ZN(n1237) );
NAND3_X1 U912 ( .A1(n1224), .A2(n1037), .A3(n1229), .ZN(n1177) );
INV_X1 U913 ( .A(n1053), .ZN(n1224) );
NAND2_X1 U914 ( .A1(n1238), .A2(n1207), .ZN(n1053) );
XOR2_X1 U915 ( .A(n1239), .B(KEYINPUT33), .Z(n1207) );
XNOR2_X1 U916 ( .A(G113), .B(n1176), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1055), .A2(n1037), .A3(n1229), .ZN(n1176) );
AND3_X1 U918 ( .A1(n1048), .A2(n1232), .A3(n1225), .ZN(n1229) );
INV_X1 U919 ( .A(n1030), .ZN(n1225) );
NAND2_X1 U920 ( .A1(n1240), .A2(n1241), .ZN(n1048) );
OR2_X1 U921 ( .A1(n1060), .A2(KEYINPUT6), .ZN(n1241) );
NAND3_X1 U922 ( .A1(n1061), .A2(n1242), .A3(KEYINPUT6), .ZN(n1240) );
NAND2_X1 U923 ( .A1(n1243), .A2(n1244), .ZN(n1037) );
NAND2_X1 U924 ( .A1(n1038), .A2(n1235), .ZN(n1244) );
INV_X1 U925 ( .A(KEYINPUT21), .ZN(n1235) );
INV_X1 U926 ( .A(n1031), .ZN(n1038) );
NAND2_X1 U927 ( .A1(n1245), .A2(n1246), .ZN(n1031) );
NAND3_X1 U928 ( .A1(n1070), .A2(n1245), .A3(KEYINPUT21), .ZN(n1243) );
INV_X1 U929 ( .A(n1047), .ZN(n1055) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1069), .ZN(n1047) );
XNOR2_X1 U931 ( .A(n1247), .B(n1248), .ZN(G12) );
NOR4_X1 U932 ( .A1(KEYINPUT34), .A2(n1174), .A3(n1182), .A4(n1026), .ZN(n1248) );
NAND2_X1 U933 ( .A1(n1238), .A2(n1239), .ZN(n1026) );
XOR2_X1 U934 ( .A(n1075), .B(n1249), .Z(n1239) );
NOR2_X1 U935 ( .A1(G478), .A2(KEYINPUT49), .ZN(n1249) );
NOR2_X1 U936 ( .A1(n1135), .A2(G902), .ZN(n1075) );
XNOR2_X1 U937 ( .A(n1250), .B(n1251), .ZN(n1135) );
XOR2_X1 U938 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U939 ( .A(G134), .B(G143), .ZN(n1253) );
NAND2_X1 U940 ( .A1(G217), .A2(n1254), .ZN(n1252) );
XNOR2_X1 U941 ( .A(n1255), .B(n1256), .ZN(n1250) );
NAND2_X1 U942 ( .A1(n1257), .A2(KEYINPUT10), .ZN(n1256) );
XOR2_X1 U943 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U944 ( .A(G107), .B(G116), .ZN(n1258) );
NAND2_X1 U945 ( .A1(KEYINPUT43), .A2(G128), .ZN(n1255) );
INV_X1 U946 ( .A(n1069), .ZN(n1238) );
XNOR2_X1 U947 ( .A(n1260), .B(G475), .ZN(n1069) );
NAND2_X1 U948 ( .A1(n1139), .A2(n1261), .ZN(n1260) );
XOR2_X1 U949 ( .A(n1262), .B(n1263), .Z(n1139) );
XOR2_X1 U950 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U951 ( .A(n1266), .B(n1267), .Z(n1265) );
AND3_X1 U952 ( .A1(G214), .A2(n1041), .A3(n1268), .ZN(n1267) );
NAND2_X1 U953 ( .A1(KEYINPUT18), .A2(n1102), .ZN(n1266) );
XNOR2_X1 U954 ( .A(G143), .B(G146), .ZN(n1264) );
XOR2_X1 U955 ( .A(n1269), .B(n1270), .Z(n1262) );
XNOR2_X1 U956 ( .A(n1271), .B(n1259), .ZN(n1270) );
NAND2_X1 U957 ( .A1(n1246), .A2(n1236), .ZN(n1182) );
XNOR2_X1 U958 ( .A(n1245), .B(KEYINPUT39), .ZN(n1236) );
XNOR2_X1 U959 ( .A(n1068), .B(KEYINPUT52), .ZN(n1245) );
XOR2_X1 U960 ( .A(n1272), .B(n1130), .Z(n1068) );
NAND2_X1 U961 ( .A1(G217), .A2(n1273), .ZN(n1130) );
NAND2_X1 U962 ( .A1(n1128), .A2(n1261), .ZN(n1272) );
XNOR2_X1 U963 ( .A(n1274), .B(n1275), .ZN(n1128) );
XOR2_X1 U964 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U965 ( .A(G119), .B(n1247), .ZN(n1277) );
XNOR2_X1 U966 ( .A(KEYINPUT8), .B(n1105), .ZN(n1276) );
INV_X1 U967 ( .A(G137), .ZN(n1105) );
XOR2_X1 U968 ( .A(n1278), .B(n1279), .Z(n1274) );
XNOR2_X1 U969 ( .A(n1280), .B(n1271), .ZN(n1279) );
INV_X1 U970 ( .A(n1096), .ZN(n1271) );
XOR2_X1 U971 ( .A(G125), .B(G140), .Z(n1096) );
NOR2_X1 U972 ( .A1(G146), .A2(KEYINPUT36), .ZN(n1280) );
XOR2_X1 U973 ( .A(n1281), .B(n1282), .Z(n1278) );
NOR2_X1 U974 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1282) );
NAND2_X1 U975 ( .A1(G221), .A2(n1254), .ZN(n1281) );
AND2_X1 U976 ( .A1(G234), .A2(n1041), .ZN(n1254) );
INV_X1 U977 ( .A(n1070), .ZN(n1246) );
XNOR2_X1 U978 ( .A(n1283), .B(G472), .ZN(n1070) );
NAND2_X1 U979 ( .A1(n1284), .A2(n1261), .ZN(n1283) );
XOR2_X1 U980 ( .A(n1285), .B(n1154), .Z(n1284) );
XOR2_X1 U981 ( .A(n1153), .B(n1152), .Z(n1154) );
XOR2_X1 U982 ( .A(n1286), .B(n1287), .Z(n1152) );
INV_X1 U983 ( .A(n1199), .ZN(n1287) );
XOR2_X1 U984 ( .A(n1288), .B(n1098), .Z(n1199) );
INV_X1 U985 ( .A(G128), .ZN(n1098) );
XNOR2_X1 U986 ( .A(n1166), .B(KEYINPUT45), .ZN(n1286) );
XNOR2_X1 U987 ( .A(n1289), .B(n1290), .ZN(n1153) );
XNOR2_X1 U988 ( .A(G113), .B(KEYINPUT29), .ZN(n1289) );
NOR2_X1 U989 ( .A1(n1291), .A2(n1292), .ZN(n1285) );
XOR2_X1 U990 ( .A(n1293), .B(KEYINPUT47), .Z(n1292) );
NAND2_X1 U991 ( .A1(n1149), .A2(G101), .ZN(n1293) );
NOR2_X1 U992 ( .A1(G101), .A2(n1149), .ZN(n1291) );
AND3_X1 U993 ( .A1(G210), .A2(n1041), .A3(n1294), .ZN(n1149) );
XNOR2_X1 U994 ( .A(G237), .B(KEYINPUT16), .ZN(n1294) );
NAND2_X1 U995 ( .A1(n1185), .A2(n1232), .ZN(n1174) );
NAND2_X1 U996 ( .A1(n1027), .A2(n1295), .ZN(n1232) );
NAND4_X1 U997 ( .A1(n1092), .A2(G902), .A3(n1228), .A4(n1117), .ZN(n1295) );
INV_X1 U998 ( .A(G898), .ZN(n1117) );
XNOR2_X1 U999 ( .A(G953), .B(KEYINPUT54), .ZN(n1092) );
NAND3_X1 U1000 ( .A1(n1228), .A2(n1041), .A3(G952), .ZN(n1027) );
INV_X1 U1001 ( .A(G953), .ZN(n1041) );
NAND2_X1 U1002 ( .A1(n1296), .A2(G234), .ZN(n1228) );
XNOR2_X1 U1003 ( .A(G237), .B(KEYINPUT63), .ZN(n1296) );
NOR2_X1 U1004 ( .A1(n1030), .A2(n1060), .ZN(n1185) );
OR2_X1 U1005 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U1006 ( .A(n1242), .ZN(n1062) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1273), .ZN(n1242) );
NAND2_X1 U1008 ( .A1(G234), .A2(n1261), .ZN(n1273) );
XOR2_X1 U1009 ( .A(G469), .B(n1297), .Z(n1061) );
NOR2_X1 U1010 ( .A1(n1076), .A2(KEYINPUT15), .ZN(n1297) );
AND2_X1 U1011 ( .A1(n1298), .A2(n1299), .ZN(n1076) );
XNOR2_X1 U1012 ( .A(n1162), .B(n1300), .ZN(n1299) );
NOR3_X1 U1013 ( .A1(n1301), .A2(KEYINPUT13), .A3(n1302), .ZN(n1300) );
NOR2_X1 U1014 ( .A1(n1303), .A2(n1165), .ZN(n1302) );
XOR2_X1 U1015 ( .A(n1304), .B(KEYINPUT48), .Z(n1301) );
NAND2_X1 U1016 ( .A1(n1303), .A2(n1165), .ZN(n1304) );
XOR2_X1 U1017 ( .A(n1305), .B(n1306), .Z(n1165) );
XNOR2_X1 U1018 ( .A(n1307), .B(KEYINPUT46), .ZN(n1306) );
NAND2_X1 U1019 ( .A1(KEYINPUT24), .A2(n1308), .ZN(n1307) );
INV_X1 U1020 ( .A(G104), .ZN(n1308) );
XOR2_X1 U1021 ( .A(n1097), .B(n1309), .Z(n1305) );
XOR2_X1 U1022 ( .A(n1310), .B(n1311), .Z(n1097) );
XNOR2_X1 U1023 ( .A(KEYINPUT2), .B(n1202), .ZN(n1311) );
NAND2_X1 U1024 ( .A1(KEYINPUT17), .A2(n1312), .ZN(n1310) );
INV_X1 U1025 ( .A(G143), .ZN(n1312) );
INV_X1 U1026 ( .A(n1166), .ZN(n1303) );
XOR2_X1 U1027 ( .A(n1313), .B(n1102), .Z(n1166) );
INV_X1 U1028 ( .A(G131), .ZN(n1102) );
NAND2_X1 U1029 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1030 ( .A1(G137), .A2(n1213), .ZN(n1315) );
XOR2_X1 U1031 ( .A(KEYINPUT40), .B(n1316), .Z(n1314) );
NOR2_X1 U1032 ( .A1(G137), .A2(n1213), .ZN(n1316) );
INV_X1 U1033 ( .A(G134), .ZN(n1213) );
XNOR2_X1 U1034 ( .A(n1317), .B(n1318), .ZN(n1162) );
XNOR2_X1 U1035 ( .A(n1247), .B(n1319), .ZN(n1318) );
NOR2_X1 U1036 ( .A1(G953), .A2(n1109), .ZN(n1319) );
INV_X1 U1037 ( .A(G227), .ZN(n1109) );
XNOR2_X1 U1038 ( .A(G140), .B(KEYINPUT61), .ZN(n1317) );
XNOR2_X1 U1039 ( .A(G902), .B(KEYINPUT12), .ZN(n1298) );
NAND2_X1 U1040 ( .A1(n1032), .A2(n1039), .ZN(n1030) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1320), .ZN(n1039) );
XNOR2_X1 U1042 ( .A(n1321), .B(n1072), .ZN(n1032) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1320), .ZN(n1072) );
NAND2_X1 U1044 ( .A1(n1268), .A2(n1261), .ZN(n1320) );
INV_X1 U1045 ( .A(G902), .ZN(n1261) );
INV_X1 U1046 ( .A(G237), .ZN(n1268) );
NAND2_X1 U1047 ( .A1(KEYINPUT59), .A2(n1074), .ZN(n1321) );
OR2_X1 U1048 ( .A1(n1201), .A2(G902), .ZN(n1074) );
XNOR2_X1 U1049 ( .A(n1322), .B(n1323), .ZN(n1201) );
XNOR2_X1 U1050 ( .A(n1288), .B(n1309), .ZN(n1323) );
XOR2_X1 U1051 ( .A(G128), .B(n1198), .Z(n1309) );
XOR2_X1 U1052 ( .A(G107), .B(G101), .Z(n1198) );
NAND2_X1 U1053 ( .A1(n1324), .A2(n1325), .ZN(n1288) );
NAND2_X1 U1054 ( .A1(G143), .A2(n1202), .ZN(n1325) );
XOR2_X1 U1055 ( .A(KEYINPUT19), .B(n1326), .Z(n1324) );
NOR2_X1 U1056 ( .A1(G143), .A2(n1202), .ZN(n1326) );
INV_X1 U1057 ( .A(G146), .ZN(n1202) );
XOR2_X1 U1058 ( .A(n1197), .B(n1200), .Z(n1322) );
XOR2_X1 U1059 ( .A(G125), .B(n1327), .Z(n1200) );
NOR2_X1 U1060 ( .A1(G953), .A2(n1125), .ZN(n1327) );
INV_X1 U1061 ( .A(G224), .ZN(n1125) );
XOR2_X1 U1062 ( .A(n1328), .B(n1329), .Z(n1197) );
XOR2_X1 U1063 ( .A(KEYINPUT27), .B(n1330), .Z(n1329) );
NOR2_X1 U1064 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1065 ( .A(KEYINPUT3), .B(n1333), .Z(n1332) );
NOR2_X1 U1066 ( .A1(n1259), .A2(n1247), .ZN(n1333) );
AND2_X1 U1067 ( .A1(n1247), .A2(n1259), .ZN(n1331) );
XOR2_X1 U1068 ( .A(G122), .B(KEYINPUT53), .Z(n1259) );
XOR2_X1 U1069 ( .A(n1269), .B(n1290), .Z(n1328) );
XOR2_X1 U1070 ( .A(G116), .B(G119), .Z(n1290) );
XNOR2_X1 U1071 ( .A(G104), .B(G113), .ZN(n1269) );
INV_X1 U1072 ( .A(G110), .ZN(n1247) );
endmodule


