//Key = 0010011101111001011110001010000011010001001101101001010010010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;

XOR2_X1 U716 ( .A(G107), .B(n990), .Z(G9) );
NOR2_X1 U717 ( .A1(n991), .A2(n992), .ZN(n990) );
XNOR2_X1 U718 ( .A(n993), .B(KEYINPUT4), .ZN(n991) );
NOR2_X1 U719 ( .A1(n994), .A2(n995), .ZN(G75) );
NOR4_X1 U720 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(n995) );
INV_X1 U721 ( .A(G952), .ZN(n998) );
NAND2_X1 U722 ( .A1(n1000), .A2(n1001), .ZN(n997) );
NOR3_X1 U723 ( .A1(n1002), .A2(KEYINPUT36), .A3(n1003), .ZN(n996) );
INV_X1 U724 ( .A(n1004), .ZN(n1003) );
NOR2_X1 U725 ( .A1(n1005), .A2(n1006), .ZN(n1002) );
NOR3_X1 U726 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NOR2_X1 U727 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR3_X1 U729 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1010) );
NOR3_X1 U730 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NOR2_X1 U731 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
XOR2_X1 U732 ( .A(n1022), .B(KEYINPUT10), .Z(n1020) );
NOR2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1015) );
NOR3_X1 U734 ( .A1(n1012), .A2(n1025), .A3(n1026), .ZN(n1005) );
INV_X1 U735 ( .A(n1027), .ZN(n1026) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1009), .ZN(n1029) );
INV_X1 U738 ( .A(n1031), .ZN(n1009) );
NOR2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U741 ( .A1(n1036), .A2(n1007), .ZN(n1028) );
NOR2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR3_X1 U743 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n994) );
NOR2_X1 U744 ( .A1(KEYINPUT1), .A2(n1042), .ZN(n1041) );
NOR2_X1 U745 ( .A1(G953), .A2(G952), .ZN(n1042) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
INV_X1 U747 ( .A(KEYINPUT1), .ZN(n1044) );
INV_X1 U748 ( .A(n1000), .ZN(n1039) );
NAND4_X1 U749 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1000) );
NOR4_X1 U750 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XNOR2_X1 U751 ( .A(G472), .B(n1053), .ZN(n1052) );
XOR2_X1 U752 ( .A(G478), .B(n1054), .Z(n1051) );
AND2_X1 U753 ( .A1(n1021), .A2(n1035), .ZN(n1047) );
XNOR2_X1 U754 ( .A(KEYINPUT24), .B(n1024), .ZN(n1046) );
INV_X1 U755 ( .A(n1017), .ZN(n1024) );
XNOR2_X1 U756 ( .A(KEYINPUT18), .B(n1055), .ZN(n1045) );
XOR2_X1 U757 ( .A(n1056), .B(n1057), .Z(G72) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1001), .ZN(n1057) );
AND2_X1 U759 ( .A1(G227), .A2(G900), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U762 ( .A(KEYINPUT33), .ZN(n1062) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(n1059) );
AND3_X1 U765 ( .A1(KEYINPUT33), .A2(n1064), .A3(n1063), .ZN(n1066) );
XNOR2_X1 U766 ( .A(n1067), .B(n1068), .ZN(n1063) );
XOR2_X1 U767 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
XOR2_X1 U769 ( .A(n1073), .B(KEYINPUT26), .Z(n1072) );
NAND2_X1 U770 ( .A1(G125), .A2(n1074), .ZN(n1073) );
NOR2_X1 U771 ( .A1(G125), .A2(n1074), .ZN(n1071) );
XOR2_X1 U772 ( .A(n1075), .B(n1076), .Z(n1067) );
NOR2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U774 ( .A(KEYINPUT16), .B(n1079), .Z(n1078) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
AND2_X1 U776 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
XOR2_X1 U777 ( .A(G134), .B(KEYINPUT49), .Z(n1081) );
XNOR2_X1 U778 ( .A(G131), .B(KEYINPUT63), .ZN(n1075) );
INV_X1 U779 ( .A(n1082), .ZN(n1064) );
NAND2_X1 U780 ( .A1(n1001), .A2(n1083), .ZN(n1065) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(G69) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(n1085) );
OR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U784 ( .A1(KEYINPUT56), .A2(n1001), .A3(n1090), .ZN(n1086) );
XOR2_X1 U785 ( .A(n1091), .B(KEYINPUT44), .Z(n1090) );
NAND3_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
XOR2_X1 U787 ( .A(n1095), .B(KEYINPUT61), .Z(n1094) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1001), .ZN(n1084) );
AND2_X1 U789 ( .A1(G224), .A2(G898), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1043), .A2(n1097), .ZN(G66) );
XOR2_X1 U791 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U792 ( .A1(n1100), .A2(n1101), .A3(KEYINPUT6), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1043), .A2(n1102), .ZN(G63) );
XOR2_X1 U794 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U795 ( .A1(KEYINPUT17), .A2(n1105), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1100), .A2(G478), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1043), .A2(n1106), .ZN(G60) );
XOR2_X1 U798 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U799 ( .A1(KEYINPUT27), .A2(n1109), .ZN(n1108) );
NAND2_X1 U800 ( .A1(n1100), .A2(G475), .ZN(n1107) );
XNOR2_X1 U801 ( .A(G104), .B(n1095), .ZN(G6) );
NOR2_X1 U802 ( .A1(n1043), .A2(n1110), .ZN(G57) );
XOR2_X1 U803 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U804 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR3_X1 U806 ( .A1(n1117), .A2(KEYINPUT31), .A3(n1118), .ZN(n1113) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
XNOR2_X1 U808 ( .A(KEYINPUT38), .B(n1121), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1043), .A2(n1122), .ZN(G54) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U812 ( .A(n1127), .B(n1128), .Z(n1126) );
AND2_X1 U813 ( .A1(G469), .A2(n1100), .ZN(n1127) );
INV_X1 U814 ( .A(n1116), .ZN(n1100) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1123) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U817 ( .A(KEYINPUT58), .B(G140), .ZN(n1129) );
NOR2_X1 U818 ( .A1(n1043), .A2(n1133), .ZN(G51) );
XOR2_X1 U819 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U820 ( .A(n1136), .B(n1137), .ZN(n1135) );
XNOR2_X1 U821 ( .A(KEYINPUT51), .B(n1138), .ZN(n1137) );
NOR3_X1 U822 ( .A1(n1116), .A2(KEYINPUT40), .A3(n1139), .ZN(n1138) );
NAND2_X1 U823 ( .A1(G902), .A2(n999), .ZN(n1116) );
NAND4_X1 U824 ( .A1(n1140), .A2(n1141), .A3(n1092), .A4(n1095), .ZN(n999) );
NAND3_X1 U825 ( .A1(n1037), .A2(n1027), .A3(n1142), .ZN(n1095) );
AND3_X1 U826 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1092) );
NAND2_X1 U827 ( .A1(n1018), .A2(n993), .ZN(n1145) );
AND4_X1 U828 ( .A1(n1146), .A2(n1033), .A3(n1038), .A4(n1027), .ZN(n993) );
INV_X1 U829 ( .A(n1083), .ZN(n1141) );
NAND4_X1 U830 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1083) );
NOR4_X1 U831 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
INV_X1 U832 ( .A(n1155), .ZN(n1154) );
AND2_X1 U833 ( .A1(n1156), .A2(n1157), .ZN(n1149) );
XNOR2_X1 U834 ( .A(n1093), .B(KEYINPUT53), .ZN(n1140) );
AND4_X1 U835 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1093) );
NAND3_X1 U836 ( .A1(n1162), .A2(n1038), .A3(n1163), .ZN(n1158) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1134) );
NOR2_X1 U838 ( .A1(n1001), .A2(G952), .ZN(n1043) );
NAND3_X1 U839 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(G48) );
OR2_X1 U840 ( .A1(n1147), .A2(G146), .ZN(n1168) );
NAND2_X1 U841 ( .A1(KEYINPUT21), .A2(n1169), .ZN(n1167) );
NAND2_X1 U842 ( .A1(G146), .A2(n1170), .ZN(n1169) );
XNOR2_X1 U843 ( .A(KEYINPUT15), .B(n1147), .ZN(n1170) );
NAND2_X1 U844 ( .A1(n1171), .A2(n1172), .ZN(n1166) );
INV_X1 U845 ( .A(KEYINPUT21), .ZN(n1172) );
NAND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
OR2_X1 U847 ( .A1(n1147), .A2(KEYINPUT15), .ZN(n1174) );
NAND3_X1 U848 ( .A1(G146), .A2(n1147), .A3(KEYINPUT15), .ZN(n1173) );
NAND3_X1 U849 ( .A1(n1175), .A2(n1018), .A3(n1037), .ZN(n1147) );
XOR2_X1 U850 ( .A(n1148), .B(n1176), .Z(G45) );
XNOR2_X1 U851 ( .A(G143), .B(KEYINPUT14), .ZN(n1176) );
NAND4_X1 U852 ( .A1(n1177), .A2(n1018), .A3(n1178), .A4(n1049), .ZN(n1148) );
XNOR2_X1 U853 ( .A(G140), .B(n1157), .ZN(G42) );
NAND3_X1 U854 ( .A1(n1023), .A2(n1033), .A3(n1179), .ZN(n1157) );
XNOR2_X1 U855 ( .A(n1080), .B(n1152), .ZN(G39) );
AND3_X1 U856 ( .A1(n1175), .A2(n1031), .A3(n1023), .ZN(n1152) );
XNOR2_X1 U857 ( .A(G134), .B(n1156), .ZN(G36) );
NAND3_X1 U858 ( .A1(n1023), .A2(n1038), .A3(n1177), .ZN(n1156) );
XNOR2_X1 U859 ( .A(G131), .B(n1155), .ZN(G33) );
NAND3_X1 U860 ( .A1(n1037), .A2(n1023), .A3(n1177), .ZN(n1155) );
AND3_X1 U861 ( .A1(n1033), .A2(n1180), .A3(n1162), .ZN(n1177) );
INV_X1 U862 ( .A(n1012), .ZN(n1023) );
NAND2_X1 U863 ( .A1(n1022), .A2(n1021), .ZN(n1012) );
XNOR2_X1 U864 ( .A(n1181), .B(KEYINPUT30), .ZN(n1022) );
XOR2_X1 U865 ( .A(n1151), .B(n1182), .Z(G30) );
NOR2_X1 U866 ( .A1(KEYINPUT52), .A2(n1183), .ZN(n1182) );
AND3_X1 U867 ( .A1(n1018), .A2(n1038), .A3(n1175), .ZN(n1151) );
AND4_X1 U868 ( .A1(n1014), .A2(n1033), .A3(n1017), .A4(n1180), .ZN(n1175) );
XNOR2_X1 U869 ( .A(G101), .B(n1143), .ZN(G3) );
NAND3_X1 U870 ( .A1(n1162), .A2(n1031), .A3(n1142), .ZN(n1143) );
XOR2_X1 U871 ( .A(G125), .B(n1153), .Z(G27) );
AND3_X1 U872 ( .A1(n1179), .A2(n1018), .A3(n1184), .ZN(n1153) );
AND4_X1 U873 ( .A1(n1037), .A2(n1017), .A3(n1185), .A4(n1180), .ZN(n1179) );
NAND2_X1 U874 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NAND3_X1 U875 ( .A1(G902), .A2(n1188), .A3(n1082), .ZN(n1187) );
NOR2_X1 U876 ( .A1(n1001), .A2(G900), .ZN(n1082) );
XNOR2_X1 U877 ( .A(KEYINPUT2), .B(n1004), .ZN(n1188) );
NAND3_X1 U878 ( .A1(n1004), .A2(n1001), .A3(G952), .ZN(n1186) );
NAND3_X1 U879 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(G24) );
OR2_X1 U880 ( .A1(n1192), .A2(KEYINPUT45), .ZN(n1191) );
NAND3_X1 U881 ( .A1(KEYINPUT45), .A2(n1192), .A3(n1193), .ZN(n1190) );
NAND2_X1 U882 ( .A1(n1194), .A2(n1195), .ZN(n1189) );
NAND2_X1 U883 ( .A1(n1196), .A2(KEYINPUT45), .ZN(n1195) );
XNOR2_X1 U884 ( .A(n1192), .B(KEYINPUT39), .ZN(n1196) );
INV_X1 U885 ( .A(n1159), .ZN(n1192) );
NAND4_X1 U886 ( .A1(n1163), .A2(n1027), .A3(n1178), .A4(n1049), .ZN(n1159) );
NOR2_X1 U887 ( .A1(n1017), .A2(n1014), .ZN(n1027) );
INV_X1 U888 ( .A(n1193), .ZN(n1194) );
XOR2_X1 U889 ( .A(G122), .B(KEYINPUT9), .Z(n1193) );
XNOR2_X1 U890 ( .A(n1160), .B(n1197), .ZN(G21) );
NOR2_X1 U891 ( .A1(KEYINPUT34), .A2(n1198), .ZN(n1197) );
NAND4_X1 U892 ( .A1(n1014), .A2(n1163), .A3(n1031), .A4(n1017), .ZN(n1160) );
INV_X1 U893 ( .A(n1185), .ZN(n1014) );
XNOR2_X1 U894 ( .A(G116), .B(n1199), .ZN(G18) );
NAND4_X1 U895 ( .A1(n1038), .A2(n1200), .A3(n1146), .A4(n1201), .ZN(n1199) );
NOR2_X1 U896 ( .A1(n992), .A2(n1013), .ZN(n1201) );
INV_X1 U897 ( .A(n1162), .ZN(n1013) );
XNOR2_X1 U898 ( .A(KEYINPUT57), .B(n1007), .ZN(n1200) );
XNOR2_X1 U899 ( .A(G113), .B(n1161), .ZN(G15) );
NAND3_X1 U900 ( .A1(n1162), .A2(n1037), .A3(n1163), .ZN(n1161) );
AND3_X1 U901 ( .A1(n1018), .A2(n1146), .A3(n1184), .ZN(n1163) );
INV_X1 U902 ( .A(n1007), .ZN(n1184) );
NAND2_X1 U903 ( .A1(n1055), .A2(n1035), .ZN(n1007) );
INV_X1 U904 ( .A(n1034), .ZN(n1055) );
NOR2_X1 U905 ( .A1(n1178), .A2(n1202), .ZN(n1037) );
INV_X1 U906 ( .A(n1203), .ZN(n1178) );
NOR2_X1 U907 ( .A1(n1185), .A2(n1017), .ZN(n1162) );
XNOR2_X1 U908 ( .A(G110), .B(n1144), .ZN(G12) );
NAND4_X1 U909 ( .A1(n1142), .A2(n1031), .A3(n1017), .A4(n1185), .ZN(n1144) );
XOR2_X1 U910 ( .A(n1204), .B(n1053), .Z(n1185) );
NAND2_X1 U911 ( .A1(n1205), .A2(n1206), .ZN(n1053) );
XNOR2_X1 U912 ( .A(n1111), .B(n1207), .ZN(n1205) );
NOR3_X1 U913 ( .A1(n1208), .A2(KEYINPUT47), .A3(n1118), .ZN(n1207) );
AND2_X1 U914 ( .A1(n1119), .A2(G101), .ZN(n1118) );
NOR2_X1 U915 ( .A1(G101), .A2(n1119), .ZN(n1208) );
AND2_X1 U916 ( .A1(n1209), .A2(G210), .ZN(n1119) );
XOR2_X1 U917 ( .A(n1128), .B(n1210), .Z(n1111) );
NOR2_X1 U918 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U919 ( .A(n1213), .B(KEYINPUT42), .Z(n1212) );
NAND2_X1 U920 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U921 ( .A1(n1215), .A2(n1214), .ZN(n1211) );
NAND2_X1 U922 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND2_X1 U923 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U924 ( .A(KEYINPUT60), .ZN(n1219) );
NAND3_X1 U925 ( .A1(G119), .A2(n1220), .A3(KEYINPUT60), .ZN(n1216) );
INV_X1 U926 ( .A(G116), .ZN(n1220) );
XNOR2_X1 U927 ( .A(n1221), .B(n1070), .ZN(n1128) );
NAND2_X1 U928 ( .A1(KEYINPUT35), .A2(n1115), .ZN(n1204) );
INV_X1 U929 ( .A(G472), .ZN(n1115) );
XNOR2_X1 U930 ( .A(n1222), .B(n1101), .ZN(n1017) );
AND2_X1 U931 ( .A1(G217), .A2(n1223), .ZN(n1101) );
NAND2_X1 U932 ( .A1(n1099), .A2(n1206), .ZN(n1222) );
XOR2_X1 U933 ( .A(n1224), .B(n1225), .Z(n1099) );
XOR2_X1 U934 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U935 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U936 ( .A1(G146), .A2(KEYINPUT25), .ZN(n1229) );
NAND2_X1 U937 ( .A1(KEYINPUT32), .A2(n1230), .ZN(n1228) );
XOR2_X1 U938 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U939 ( .A(n1198), .B(G110), .ZN(n1232) );
INV_X1 U940 ( .A(G119), .ZN(n1198) );
XNOR2_X1 U941 ( .A(KEYINPUT5), .B(n1183), .ZN(n1231) );
NOR2_X1 U942 ( .A1(n1233), .A2(n1234), .ZN(n1226) );
INV_X1 U943 ( .A(G221), .ZN(n1233) );
XOR2_X1 U944 ( .A(n1235), .B(n1236), .Z(n1224) );
XNOR2_X1 U945 ( .A(KEYINPUT19), .B(n1074), .ZN(n1236) );
INV_X1 U946 ( .A(G140), .ZN(n1074) );
XNOR2_X1 U947 ( .A(G137), .B(G125), .ZN(n1235) );
NAND2_X1 U948 ( .A1(n1237), .A2(n1238), .ZN(n1031) );
NAND2_X1 U949 ( .A1(n1038), .A2(n1239), .ZN(n1238) );
INV_X1 U950 ( .A(KEYINPUT20), .ZN(n1239) );
NOR2_X1 U951 ( .A1(n1049), .A2(n1203), .ZN(n1038) );
NAND3_X1 U952 ( .A1(n1203), .A2(n1202), .A3(KEYINPUT20), .ZN(n1237) );
INV_X1 U953 ( .A(n1049), .ZN(n1202) );
XNOR2_X1 U954 ( .A(n1240), .B(G475), .ZN(n1049) );
OR2_X1 U955 ( .A1(n1109), .A2(G902), .ZN(n1240) );
XNOR2_X1 U956 ( .A(n1241), .B(n1242), .ZN(n1109) );
XOR2_X1 U957 ( .A(n1136), .B(n1243), .Z(n1242) );
XNOR2_X1 U958 ( .A(G104), .B(n1244), .ZN(n1243) );
NAND2_X1 U959 ( .A1(KEYINPUT48), .A2(n1245), .ZN(n1244) );
NAND2_X1 U960 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND3_X1 U961 ( .A1(G214), .A2(n1248), .A3(n1209), .ZN(n1247) );
XNOR2_X1 U962 ( .A(KEYINPUT3), .B(n1249), .ZN(n1248) );
XOR2_X1 U963 ( .A(n1250), .B(KEYINPUT28), .Z(n1246) );
NAND2_X1 U964 ( .A1(n1249), .A2(n1251), .ZN(n1250) );
NAND2_X1 U965 ( .A1(n1209), .A2(G214), .ZN(n1251) );
NOR2_X1 U966 ( .A1(G237), .A2(G953), .ZN(n1209) );
INV_X1 U967 ( .A(G143), .ZN(n1249) );
XOR2_X1 U968 ( .A(G125), .B(n1252), .Z(n1136) );
XOR2_X1 U969 ( .A(n1253), .B(n1254), .Z(n1241) );
XOR2_X1 U970 ( .A(KEYINPUT13), .B(G146), .Z(n1254) );
XNOR2_X1 U971 ( .A(G131), .B(G140), .ZN(n1253) );
XOR2_X1 U972 ( .A(G478), .B(n1255), .Z(n1203) );
NOR2_X1 U973 ( .A1(KEYINPUT54), .A2(n1256), .ZN(n1255) );
XOR2_X1 U974 ( .A(KEYINPUT8), .B(n1054), .Z(n1256) );
NOR2_X1 U975 ( .A1(n1257), .A2(n1105), .ZN(n1054) );
XOR2_X1 U976 ( .A(n1258), .B(n1259), .Z(n1105) );
XOR2_X1 U977 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U978 ( .A(G107), .B(n1262), .Z(n1261) );
NOR2_X1 U979 ( .A1(n1234), .A2(n1263), .ZN(n1262) );
INV_X1 U980 ( .A(G217), .ZN(n1263) );
NAND2_X1 U981 ( .A1(n1264), .A2(n1001), .ZN(n1234) );
XNOR2_X1 U982 ( .A(G234), .B(KEYINPUT12), .ZN(n1264) );
XNOR2_X1 U983 ( .A(G116), .B(n1265), .ZN(n1258) );
XNOR2_X1 U984 ( .A(n1266), .B(G122), .ZN(n1265) );
INV_X1 U985 ( .A(G134), .ZN(n1266) );
XNOR2_X1 U986 ( .A(KEYINPUT7), .B(G902), .ZN(n1257) );
AND3_X1 U987 ( .A1(n1146), .A2(n1033), .A3(n1018), .ZN(n1142) );
INV_X1 U988 ( .A(n992), .ZN(n1018) );
NAND2_X1 U989 ( .A1(n1181), .A2(n1021), .ZN(n992) );
NAND2_X1 U990 ( .A1(G214), .A2(n1267), .ZN(n1021) );
XOR2_X1 U991 ( .A(n1050), .B(KEYINPUT37), .Z(n1181) );
XOR2_X1 U992 ( .A(n1268), .B(n1139), .Z(n1050) );
NAND2_X1 U993 ( .A1(G210), .A2(n1267), .ZN(n1139) );
NAND2_X1 U994 ( .A1(n1269), .A2(n1206), .ZN(n1267) );
INV_X1 U995 ( .A(G237), .ZN(n1269) );
NAND3_X1 U996 ( .A1(n1270), .A2(n1206), .A3(n1271), .ZN(n1268) );
XOR2_X1 U997 ( .A(KEYINPUT11), .B(n1272), .Z(n1271) );
NOR2_X1 U998 ( .A1(n1273), .A2(n1088), .ZN(n1272) );
NAND2_X1 U999 ( .A1(n1273), .A2(n1088), .ZN(n1270) );
XNOR2_X1 U1000 ( .A(n1252), .B(n1165), .ZN(n1088) );
XNOR2_X1 U1001 ( .A(n1274), .B(n1125), .ZN(n1165) );
XNOR2_X1 U1002 ( .A(n1275), .B(G101), .ZN(n1125) );
INV_X1 U1003 ( .A(G110), .ZN(n1275) );
XOR2_X1 U1004 ( .A(n1218), .B(n1276), .Z(n1274) );
NOR2_X1 U1005 ( .A1(KEYINPUT22), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U1006 ( .A(G107), .B(n1278), .ZN(n1277) );
INV_X1 U1007 ( .A(G104), .ZN(n1278) );
XNOR2_X1 U1008 ( .A(G116), .B(G119), .ZN(n1218) );
XNOR2_X1 U1009 ( .A(G122), .B(n1215), .ZN(n1252) );
INV_X1 U1010 ( .A(G113), .ZN(n1215) );
XOR2_X1 U1011 ( .A(n1164), .B(n1279), .Z(n1273) );
NOR2_X1 U1012 ( .A1(G125), .A2(KEYINPUT62), .ZN(n1279) );
XOR2_X1 U1013 ( .A(n1280), .B(n1070), .Z(n1164) );
NAND2_X1 U1014 ( .A1(G224), .A2(n1001), .ZN(n1280) );
AND2_X1 U1015 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1223), .ZN(n1035) );
NAND2_X1 U1017 ( .A1(G234), .A2(n1206), .ZN(n1223) );
XNOR2_X1 U1018 ( .A(n1281), .B(G469), .ZN(n1034) );
NAND2_X1 U1019 ( .A1(n1282), .A2(n1206), .ZN(n1281) );
INV_X1 U1020 ( .A(G902), .ZN(n1206) );
XOR2_X1 U1021 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1022 ( .A(n1221), .B(n1285), .Z(n1284) );
NOR2_X1 U1023 ( .A1(KEYINPUT50), .A2(n1131), .ZN(n1285) );
NAND2_X1 U1024 ( .A1(G227), .A2(n1001), .ZN(n1131) );
XOR2_X1 U1025 ( .A(n1286), .B(KEYINPUT46), .Z(n1221) );
NAND3_X1 U1026 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1286) );
OR2_X1 U1027 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND3_X1 U1028 ( .A1(n1291), .A2(n1290), .A3(G131), .ZN(n1288) );
NAND2_X1 U1029 ( .A1(n1292), .A2(n1293), .ZN(n1287) );
INV_X1 U1030 ( .A(G131), .ZN(n1293) );
NAND2_X1 U1031 ( .A1(n1294), .A2(n1290), .ZN(n1292) );
INV_X1 U1032 ( .A(KEYINPUT0), .ZN(n1290) );
XNOR2_X1 U1033 ( .A(n1291), .B(KEYINPUT59), .ZN(n1294) );
XNOR2_X1 U1034 ( .A(G134), .B(n1080), .ZN(n1291) );
INV_X1 U1035 ( .A(G137), .ZN(n1080) );
XOR2_X1 U1036 ( .A(n1295), .B(n1296), .Z(n1283) );
NOR2_X1 U1037 ( .A1(KEYINPUT29), .A2(n1297), .ZN(n1296) );
NOR2_X1 U1038 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U1039 ( .A(KEYINPUT23), .B(n1300), .Z(n1299) );
NOR2_X1 U1040 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XNOR2_X1 U1041 ( .A(n1121), .B(n1132), .ZN(n1302) );
INV_X1 U1042 ( .A(G101), .ZN(n1121) );
XNOR2_X1 U1043 ( .A(n1303), .B(KEYINPUT41), .ZN(n1301) );
NOR2_X1 U1044 ( .A1(n1304), .A2(n1303), .ZN(n1298) );
XNOR2_X1 U1045 ( .A(n1305), .B(n1070), .ZN(n1303) );
XOR2_X1 U1046 ( .A(G146), .B(n1260), .Z(n1070) );
XNOR2_X1 U1047 ( .A(n1183), .B(G143), .ZN(n1260) );
INV_X1 U1048 ( .A(G128), .ZN(n1183) );
XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(KEYINPUT43), .ZN(n1305) );
XNOR2_X1 U1050 ( .A(G101), .B(n1132), .ZN(n1304) );
NOR2_X1 U1051 ( .A1(KEYINPUT55), .A2(n1306), .ZN(n1132) );
XNOR2_X1 U1052 ( .A(G104), .B(G107), .ZN(n1306) );
XNOR2_X1 U1053 ( .A(G110), .B(G140), .ZN(n1295) );
AND2_X1 U1054 ( .A1(n1307), .A2(n1004), .ZN(n1146) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1004) );
NAND2_X1 U1056 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1057 ( .A1(G902), .A2(n1089), .ZN(n1309) );
NOR2_X1 U1058 ( .A1(n1001), .A2(G898), .ZN(n1089) );
NAND2_X1 U1059 ( .A1(G952), .A2(n1001), .ZN(n1308) );
INV_X1 U1060 ( .A(G953), .ZN(n1001) );
endmodule


