//Key = 0010101001001101000011011110011011000111010111111110100111101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396;

XNOR2_X1 U775 ( .A(G107), .B(n1063), .ZN(G9) );
NAND4_X1 U776 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(G75) );
NAND3_X1 U777 ( .A1(KEYINPUT31), .A2(n1068), .A3(n1069), .ZN(n1067) );
NAND2_X1 U778 ( .A1(G952), .A2(n1070), .ZN(n1066) );
NAND3_X1 U779 ( .A1(n1071), .A2(n1068), .A3(n1072), .ZN(n1070) );
NAND2_X1 U780 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NAND2_X1 U781 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND4_X1 U782 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
NAND2_X1 U783 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U785 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U786 ( .A1(n1085), .A2(n1087), .ZN(n1081) );
OR2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND4_X1 U788 ( .A1(n1085), .A2(n1083), .A3(n1090), .A4(n1091), .ZN(n1075) );
NAND2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND3_X1 U790 ( .A1(n1078), .A2(n1086), .A3(n1077), .ZN(n1093) );
INV_X1 U791 ( .A(KEYINPUT3), .ZN(n1086) );
INV_X1 U792 ( .A(n1080), .ZN(n1092) );
NAND3_X1 U793 ( .A1(n1094), .A2(n1095), .A3(n1080), .ZN(n1090) );
NAND2_X1 U794 ( .A1(n1077), .A2(n1096), .ZN(n1095) );
OR2_X1 U795 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U796 ( .A1(n1078), .A2(n1099), .ZN(n1094) );
NAND2_X1 U797 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U799 ( .A(n1104), .ZN(n1073) );
OR2_X1 U800 ( .A1(n1068), .A2(KEYINPUT31), .ZN(n1064) );
NAND2_X1 U801 ( .A1(n1105), .A2(n1106), .ZN(n1068) );
NOR4_X1 U802 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1106) );
XOR2_X1 U803 ( .A(n1080), .B(KEYINPUT33), .Z(n1110) );
XOR2_X1 U804 ( .A(n1111), .B(n1112), .Z(n1109) );
XOR2_X1 U805 ( .A(KEYINPUT56), .B(G478), .Z(n1112) );
NOR2_X1 U806 ( .A1(n1113), .A2(n1114), .ZN(n1108) );
INV_X1 U807 ( .A(n1115), .ZN(n1107) );
NOR4_X1 U808 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1105) );
XNOR2_X1 U809 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR2_X1 U810 ( .A1(KEYINPUT63), .A2(n1122), .ZN(n1121) );
INV_X1 U811 ( .A(G475), .ZN(n1122) );
INV_X1 U812 ( .A(n1077), .ZN(n1118) );
XOR2_X1 U813 ( .A(n1123), .B(n1124), .Z(G72) );
XOR2_X1 U814 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U815 ( .A1(n1065), .A2(n1127), .ZN(n1126) );
NAND2_X1 U816 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND2_X1 U817 ( .A1(G953), .A2(n1130), .ZN(n1129) );
XNOR2_X1 U818 ( .A(KEYINPUT39), .B(n1131), .ZN(n1130) );
XOR2_X1 U819 ( .A(n1132), .B(n1133), .Z(n1128) );
XOR2_X1 U820 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U821 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U822 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
INV_X1 U823 ( .A(n1140), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U826 ( .A1(n1140), .A2(n1145), .ZN(n1136) );
NAND2_X1 U827 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1148), .A2(n1144), .ZN(n1147) );
NAND2_X1 U829 ( .A1(G134), .A2(n1143), .ZN(n1146) );
XOR2_X1 U830 ( .A(G131), .B(KEYINPUT18), .Z(n1143) );
NOR2_X1 U831 ( .A1(G137), .A2(KEYINPUT35), .ZN(n1140) );
XNOR2_X1 U832 ( .A(n1149), .B(KEYINPUT52), .ZN(n1132) );
NAND2_X1 U833 ( .A1(KEYINPUT58), .A2(n1150), .ZN(n1149) );
NAND3_X1 U834 ( .A1(n1151), .A2(n1152), .A3(KEYINPUT38), .ZN(n1123) );
NAND2_X1 U835 ( .A1(G900), .A2(G227), .ZN(n1152) );
XOR2_X1 U836 ( .A(KEYINPUT5), .B(G953), .Z(n1151) );
XOR2_X1 U837 ( .A(n1153), .B(n1154), .Z(G69) );
XOR2_X1 U838 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U839 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U840 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U841 ( .A1(KEYINPUT37), .A2(n1161), .ZN(n1159) );
NAND2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1155) );
XOR2_X1 U843 ( .A(KEYINPUT45), .B(G953), .Z(n1162) );
NAND2_X1 U844 ( .A1(G953), .A2(n1164), .ZN(n1153) );
NAND2_X1 U845 ( .A1(G898), .A2(G224), .ZN(n1164) );
NOR2_X1 U846 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XOR2_X1 U847 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U848 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
XOR2_X1 U849 ( .A(KEYINPUT43), .B(G217), .Z(n1170) );
NOR2_X1 U850 ( .A1(n1171), .A2(n1172), .ZN(G63) );
XNOR2_X1 U851 ( .A(n1165), .B(KEYINPUT6), .ZN(n1172) );
NOR3_X1 U852 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1171) );
NOR2_X1 U853 ( .A1(KEYINPUT26), .A2(n1176), .ZN(n1175) );
NOR2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1174) );
NOR2_X1 U855 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NOR2_X1 U856 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NOR2_X1 U857 ( .A1(n1072), .A2(n1183), .ZN(n1181) );
NOR3_X1 U858 ( .A1(n1169), .A2(n1184), .A3(n1183), .ZN(n1173) );
NOR2_X1 U859 ( .A1(n1182), .A2(n1178), .ZN(n1184) );
INV_X1 U860 ( .A(KEYINPUT26), .ZN(n1178) );
NOR2_X1 U861 ( .A1(n1165), .A2(n1185), .ZN(G60) );
XOR2_X1 U862 ( .A(n1186), .B(n1187), .Z(n1185) );
NAND4_X1 U863 ( .A1(n1188), .A2(KEYINPUT55), .A3(G475), .A4(n1189), .ZN(n1187) );
XOR2_X1 U864 ( .A(n1190), .B(KEYINPUT57), .Z(n1188) );
NAND2_X1 U865 ( .A1(n1191), .A2(n1192), .ZN(G6) );
OR2_X1 U866 ( .A1(n1193), .A2(G104), .ZN(n1192) );
NAND2_X1 U867 ( .A1(G104), .A2(n1194), .ZN(n1191) );
NAND2_X1 U868 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U869 ( .A1(KEYINPUT19), .A2(n1197), .ZN(n1196) );
NAND2_X1 U870 ( .A1(n1193), .A2(n1198), .ZN(n1195) );
INV_X1 U871 ( .A(KEYINPUT19), .ZN(n1198) );
NAND2_X1 U872 ( .A1(KEYINPUT46), .A2(n1197), .ZN(n1193) );
NOR2_X1 U873 ( .A1(n1165), .A2(n1199), .ZN(G57) );
XNOR2_X1 U874 ( .A(n1200), .B(n1201), .ZN(n1199) );
XOR2_X1 U875 ( .A(G101), .B(n1202), .Z(n1201) );
NOR2_X1 U876 ( .A1(KEYINPUT14), .A2(n1203), .ZN(n1202) );
XNOR2_X1 U877 ( .A(n1204), .B(n1205), .ZN(n1203) );
XOR2_X1 U878 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR3_X1 U879 ( .A1(n1169), .A2(KEYINPUT1), .A3(n1208), .ZN(n1206) );
INV_X1 U880 ( .A(G472), .ZN(n1208) );
NOR2_X1 U881 ( .A1(n1165), .A2(n1209), .ZN(G54) );
XOR2_X1 U882 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U883 ( .A(n1212), .B(n1213), .Z(n1211) );
NAND3_X1 U884 ( .A1(G227), .A2(n1065), .A3(KEYINPUT50), .ZN(n1212) );
XOR2_X1 U885 ( .A(n1214), .B(n1215), .Z(n1210) );
NOR2_X1 U886 ( .A1(n1216), .A2(n1169), .ZN(n1215) );
INV_X1 U887 ( .A(G469), .ZN(n1216) );
NAND2_X1 U888 ( .A1(n1217), .A2(KEYINPUT47), .ZN(n1214) );
XOR2_X1 U889 ( .A(n1218), .B(n1219), .Z(n1217) );
NAND2_X1 U890 ( .A1(KEYINPUT49), .A2(n1220), .ZN(n1218) );
NOR2_X1 U891 ( .A1(n1165), .A2(n1221), .ZN(G51) );
XOR2_X1 U892 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U893 ( .A(n1224), .B(n1225), .Z(n1223) );
NOR2_X1 U894 ( .A1(n1114), .A2(n1169), .ZN(n1224) );
NAND2_X1 U895 ( .A1(G902), .A2(n1189), .ZN(n1169) );
INV_X1 U896 ( .A(n1072), .ZN(n1189) );
NOR2_X1 U897 ( .A1(n1163), .A2(n1127), .ZN(n1072) );
NAND2_X1 U898 ( .A1(n1226), .A2(n1227), .ZN(n1127) );
AND4_X1 U899 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
AND4_X1 U900 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1226) );
NAND3_X1 U901 ( .A1(n1236), .A2(n1088), .A3(n1098), .ZN(n1235) );
NAND4_X1 U902 ( .A1(n1237), .A2(n1063), .A3(n1238), .A4(n1239), .ZN(n1163) );
NOR4_X1 U903 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1197), .ZN(n1239) );
AND2_X1 U904 ( .A1(n1098), .A2(n1243), .ZN(n1197) );
NOR3_X1 U905 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1238) );
AND2_X1 U906 ( .A1(KEYINPUT4), .A2(n1247), .ZN(n1246) );
NOR3_X1 U907 ( .A1(KEYINPUT4), .A2(n1083), .A3(n1248), .ZN(n1245) );
INV_X1 U908 ( .A(n1249), .ZN(n1244) );
NAND2_X1 U909 ( .A1(n1243), .A2(n1097), .ZN(n1063) );
AND3_X1 U910 ( .A1(n1250), .A2(n1251), .A3(n1083), .ZN(n1243) );
INV_X1 U911 ( .A(n1252), .ZN(n1083) );
XOR2_X1 U912 ( .A(n1253), .B(n1254), .Z(n1222) );
XOR2_X1 U913 ( .A(KEYINPUT28), .B(n1255), .Z(n1254) );
NOR2_X1 U914 ( .A1(KEYINPUT59), .A2(n1256), .ZN(n1253) );
NOR2_X1 U915 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U916 ( .A(n1259), .B(KEYINPUT62), .Z(n1258) );
NAND2_X1 U917 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NOR2_X1 U918 ( .A1(n1261), .A2(n1260), .ZN(n1257) );
XOR2_X1 U919 ( .A(n1262), .B(KEYINPUT51), .Z(n1260) );
NOR2_X1 U920 ( .A1(n1065), .A2(G952), .ZN(n1165) );
XOR2_X1 U921 ( .A(n1232), .B(n1263), .Z(G48) );
XOR2_X1 U922 ( .A(n1264), .B(KEYINPUT11), .Z(n1263) );
NAND3_X1 U923 ( .A1(n1265), .A2(n1098), .A3(n1266), .ZN(n1232) );
XOR2_X1 U924 ( .A(n1267), .B(n1234), .Z(G45) );
NAND4_X1 U925 ( .A1(n1266), .A2(n1088), .A3(n1268), .A4(n1269), .ZN(n1234) );
XNOR2_X1 U926 ( .A(G140), .B(n1233), .ZN(G42) );
NAND3_X1 U927 ( .A1(n1089), .A2(n1098), .A3(n1236), .ZN(n1233) );
XNOR2_X1 U928 ( .A(G137), .B(n1231), .ZN(G39) );
NAND3_X1 U929 ( .A1(n1265), .A2(n1078), .A3(n1236), .ZN(n1231) );
XOR2_X1 U930 ( .A(n1144), .B(n1230), .Z(G36) );
NAND3_X1 U931 ( .A1(n1088), .A2(n1097), .A3(n1236), .ZN(n1230) );
XOR2_X1 U932 ( .A(n1148), .B(n1270), .Z(G33) );
NAND3_X1 U933 ( .A1(n1098), .A2(n1271), .A3(n1236), .ZN(n1270) );
AND4_X1 U934 ( .A1(n1085), .A2(n1251), .A3(n1080), .A4(n1272), .ZN(n1236) );
INV_X1 U935 ( .A(n1273), .ZN(n1085) );
XOR2_X1 U936 ( .A(KEYINPUT22), .B(n1088), .Z(n1271) );
XOR2_X1 U937 ( .A(n1274), .B(n1229), .Z(G30) );
NAND3_X1 U938 ( .A1(n1265), .A2(n1097), .A3(n1266), .ZN(n1229) );
AND2_X1 U939 ( .A1(n1275), .A2(n1251), .ZN(n1266) );
XOR2_X1 U940 ( .A(n1276), .B(n1249), .Z(G3) );
NAND2_X1 U941 ( .A1(n1277), .A2(n1088), .ZN(n1249) );
XOR2_X1 U942 ( .A(n1262), .B(n1228), .Z(G27) );
NAND4_X1 U943 ( .A1(n1275), .A2(n1089), .A3(n1098), .A4(n1077), .ZN(n1228) );
AND3_X1 U944 ( .A1(n1080), .A2(n1272), .A3(n1273), .ZN(n1275) );
NAND2_X1 U945 ( .A1(n1278), .A2(n1104), .ZN(n1272) );
NAND4_X1 U946 ( .A1(n1131), .A2(G953), .A3(G902), .A4(n1279), .ZN(n1278) );
XNOR2_X1 U947 ( .A(KEYINPUT32), .B(n1280), .ZN(n1279) );
XNOR2_X1 U948 ( .A(G900), .B(KEYINPUT54), .ZN(n1131) );
XOR2_X1 U949 ( .A(G122), .B(n1247), .Z(G24) );
NOR2_X1 U950 ( .A1(n1248), .A2(n1252), .ZN(n1247) );
NAND2_X1 U951 ( .A1(n1281), .A2(n1282), .ZN(n1252) );
NAND3_X1 U952 ( .A1(n1268), .A2(n1269), .A3(n1283), .ZN(n1248) );
NAND2_X1 U953 ( .A1(n1284), .A2(n1285), .ZN(G21) );
NAND2_X1 U954 ( .A1(n1242), .A2(n1286), .ZN(n1285) );
XOR2_X1 U955 ( .A(KEYINPUT20), .B(n1287), .Z(n1284) );
NOR2_X1 U956 ( .A1(n1242), .A2(n1286), .ZN(n1287) );
INV_X1 U957 ( .A(G119), .ZN(n1286) );
AND3_X1 U958 ( .A1(n1283), .A2(n1078), .A3(n1265), .ZN(n1242) );
NOR2_X1 U959 ( .A1(n1282), .A2(n1281), .ZN(n1265) );
XNOR2_X1 U960 ( .A(n1241), .B(n1288), .ZN(G18) );
XOR2_X1 U961 ( .A(KEYINPUT2), .B(G116), .Z(n1288) );
AND3_X1 U962 ( .A1(n1283), .A2(n1097), .A3(n1088), .ZN(n1241) );
NAND2_X1 U963 ( .A1(n1289), .A2(n1290), .ZN(n1097) );
NAND2_X1 U964 ( .A1(n1078), .A2(n1291), .ZN(n1290) );
INV_X1 U965 ( .A(KEYINPUT21), .ZN(n1291) );
NAND3_X1 U966 ( .A1(n1292), .A2(n1269), .A3(KEYINPUT21), .ZN(n1289) );
XOR2_X1 U967 ( .A(n1240), .B(n1293), .Z(G15) );
NOR2_X1 U968 ( .A1(KEYINPUT40), .A2(n1294), .ZN(n1293) );
INV_X1 U969 ( .A(G113), .ZN(n1294) );
AND3_X1 U970 ( .A1(n1088), .A2(n1283), .A3(n1098), .ZN(n1240) );
NOR2_X1 U971 ( .A1(n1269), .A2(n1292), .ZN(n1098) );
AND2_X1 U972 ( .A1(n1077), .A2(n1250), .ZN(n1283) );
NOR2_X1 U973 ( .A1(n1295), .A2(n1103), .ZN(n1077) );
NOR2_X1 U974 ( .A1(n1296), .A2(n1281), .ZN(n1088) );
XNOR2_X1 U975 ( .A(G110), .B(n1237), .ZN(G12) );
NAND2_X1 U976 ( .A1(n1277), .A2(n1089), .ZN(n1237) );
NOR2_X1 U977 ( .A1(n1282), .A2(n1117), .ZN(n1089) );
INV_X1 U978 ( .A(n1281), .ZN(n1117) );
XOR2_X1 U979 ( .A(n1297), .B(G472), .Z(n1281) );
NAND3_X1 U980 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
XOR2_X1 U981 ( .A(n1190), .B(KEYINPUT36), .Z(n1300) );
NAND2_X1 U982 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND2_X1 U983 ( .A1(KEYINPUT23), .A2(n1276), .ZN(n1302) );
XOR2_X1 U984 ( .A(n1303), .B(n1304), .Z(n1301) );
AND2_X1 U985 ( .A1(n1200), .A2(KEYINPUT60), .ZN(n1303) );
NAND3_X1 U986 ( .A1(n1305), .A2(n1276), .A3(KEYINPUT23), .ZN(n1298) );
XOR2_X1 U987 ( .A(n1306), .B(n1304), .Z(n1305) );
XNOR2_X1 U988 ( .A(n1307), .B(n1204), .ZN(n1304) );
XNOR2_X1 U989 ( .A(n1308), .B(n1309), .ZN(n1204) );
XOR2_X1 U990 ( .A(n1310), .B(n1311), .Z(n1308) );
NAND2_X1 U991 ( .A1(KEYINPUT25), .A2(n1207), .ZN(n1307) );
INV_X1 U992 ( .A(n1261), .ZN(n1207) );
NOR2_X1 U993 ( .A1(n1312), .A2(n1200), .ZN(n1306) );
NAND2_X1 U994 ( .A1(G210), .A2(n1313), .ZN(n1200) );
INV_X1 U995 ( .A(KEYINPUT60), .ZN(n1312) );
INV_X1 U996 ( .A(n1296), .ZN(n1282) );
XNOR2_X1 U997 ( .A(n1116), .B(KEYINPUT41), .ZN(n1296) );
XNOR2_X1 U998 ( .A(n1314), .B(n1315), .ZN(n1116) );
NOR2_X1 U999 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
OR2_X1 U1000 ( .A1(n1168), .A2(G902), .ZN(n1314) );
XNOR2_X1 U1001 ( .A(n1318), .B(n1319), .ZN(n1168) );
XNOR2_X1 U1002 ( .A(n1320), .B(n1321), .ZN(n1319) );
XOR2_X1 U1003 ( .A(n1150), .B(n1322), .Z(n1321) );
NOR4_X1 U1004 ( .A1(KEYINPUT34), .A2(G953), .A3(n1323), .A4(n1324), .ZN(n1322) );
INV_X1 U1005 ( .A(n1325), .ZN(n1150) );
XOR2_X1 U1006 ( .A(n1326), .B(n1327), .Z(n1318) );
NOR2_X1 U1007 ( .A1(KEYINPUT53), .A2(G119), .ZN(n1327) );
XNOR2_X1 U1008 ( .A(G110), .B(G137), .ZN(n1326) );
AND3_X1 U1009 ( .A1(n1250), .A2(n1251), .A3(n1078), .ZN(n1277) );
NOR2_X1 U1010 ( .A1(n1269), .A2(n1268), .ZN(n1078) );
INV_X1 U1011 ( .A(n1292), .ZN(n1268) );
XOR2_X1 U1012 ( .A(n1120), .B(G475), .Z(n1292) );
NAND2_X1 U1013 ( .A1(n1190), .A2(n1186), .ZN(n1120) );
NAND3_X1 U1014 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1186) );
NAND2_X1 U1015 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1016 ( .A1(KEYINPUT8), .A2(n1333), .ZN(n1329) );
NAND2_X1 U1017 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1018 ( .A(n1332), .B(KEYINPUT42), .ZN(n1334) );
NAND2_X1 U1019 ( .A1(n1336), .A2(n1337), .ZN(n1328) );
INV_X1 U1020 ( .A(KEYINPUT8), .ZN(n1337) );
NAND2_X1 U1021 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
OR3_X1 U1022 ( .A1(n1331), .A2(n1332), .A3(KEYINPUT42), .ZN(n1339) );
INV_X1 U1023 ( .A(n1335), .ZN(n1331) );
XOR2_X1 U1024 ( .A(n1340), .B(n1341), .Z(n1335) );
XOR2_X1 U1025 ( .A(n1342), .B(n1325), .Z(n1341) );
XOR2_X1 U1026 ( .A(G140), .B(G125), .Z(n1325) );
NOR2_X1 U1027 ( .A1(G131), .A2(KEYINPUT10), .ZN(n1342) );
XOR2_X1 U1028 ( .A(n1343), .B(n1344), .Z(n1340) );
XOR2_X1 U1029 ( .A(G146), .B(G143), .Z(n1344) );
NAND2_X1 U1030 ( .A1(G214), .A2(n1313), .ZN(n1343) );
NOR2_X1 U1031 ( .A1(G953), .A2(G237), .ZN(n1313) );
NAND2_X1 U1032 ( .A1(KEYINPUT42), .A2(n1332), .ZN(n1338) );
XOR2_X1 U1033 ( .A(G104), .B(n1345), .Z(n1332) );
XOR2_X1 U1034 ( .A(G122), .B(G113), .Z(n1345) );
NAND3_X1 U1035 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1269) );
NAND2_X1 U1036 ( .A1(G478), .A2(n1111), .ZN(n1348) );
NAND2_X1 U1037 ( .A1(n1349), .A2(n1350), .ZN(n1347) );
INV_X1 U1038 ( .A(KEYINPUT12), .ZN(n1350) );
NAND2_X1 U1039 ( .A1(n1351), .A2(n1183), .ZN(n1349) );
INV_X1 U1040 ( .A(G478), .ZN(n1183) );
XOR2_X1 U1041 ( .A(KEYINPUT16), .B(n1180), .Z(n1351) );
INV_X1 U1042 ( .A(n1111), .ZN(n1180) );
NAND2_X1 U1043 ( .A1(KEYINPUT12), .A2(n1352), .ZN(n1346) );
NAND2_X1 U1044 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1045 ( .A1(KEYINPUT16), .A2(n1111), .ZN(n1354) );
OR3_X1 U1046 ( .A1(G478), .A2(KEYINPUT16), .A3(n1111), .ZN(n1353) );
NAND2_X1 U1047 ( .A1(n1176), .A2(n1190), .ZN(n1111) );
INV_X1 U1048 ( .A(n1182), .ZN(n1176) );
XOR2_X1 U1049 ( .A(n1355), .B(n1356), .Z(n1182) );
XNOR2_X1 U1050 ( .A(n1357), .B(n1358), .ZN(n1356) );
XOR2_X1 U1051 ( .A(n1359), .B(n1360), .Z(n1358) );
NOR3_X1 U1052 ( .A1(n1317), .A2(G953), .A3(n1323), .ZN(n1360) );
INV_X1 U1053 ( .A(G217), .ZN(n1317) );
NAND2_X1 U1054 ( .A1(KEYINPUT30), .A2(n1267), .ZN(n1359) );
XOR2_X1 U1055 ( .A(n1361), .B(n1362), .Z(n1355) );
XOR2_X1 U1056 ( .A(G134), .B(G128), .Z(n1362) );
XOR2_X1 U1057 ( .A(n1311), .B(G122), .Z(n1361) );
INV_X1 U1058 ( .A(n1100), .ZN(n1251) );
NAND2_X1 U1059 ( .A1(n1363), .A2(n1295), .ZN(n1100) );
INV_X1 U1060 ( .A(n1102), .ZN(n1295) );
XOR2_X1 U1061 ( .A(n1364), .B(G469), .Z(n1102) );
NAND2_X1 U1062 ( .A1(n1365), .A2(n1190), .ZN(n1364) );
XOR2_X1 U1063 ( .A(n1366), .B(n1367), .Z(n1365) );
XOR2_X1 U1064 ( .A(n1219), .B(n1213), .Z(n1367) );
XOR2_X1 U1065 ( .A(G140), .B(G110), .Z(n1213) );
XNOR2_X1 U1066 ( .A(n1134), .B(n1310), .ZN(n1219) );
XNOR2_X1 U1067 ( .A(n1368), .B(n1369), .ZN(n1310) );
XOR2_X1 U1068 ( .A(KEYINPUT9), .B(G137), .Z(n1369) );
NAND2_X1 U1069 ( .A1(n1141), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1070 ( .A1(G131), .A2(n1144), .ZN(n1370) );
INV_X1 U1071 ( .A(G134), .ZN(n1144) );
NAND2_X1 U1072 ( .A1(G134), .A2(n1148), .ZN(n1141) );
INV_X1 U1073 ( .A(G131), .ZN(n1148) );
XOR2_X1 U1074 ( .A(n1371), .B(G128), .Z(n1134) );
NAND3_X1 U1075 ( .A1(n1372), .A2(n1373), .A3(n1374), .ZN(n1371) );
NAND2_X1 U1076 ( .A1(KEYINPUT7), .A2(G143), .ZN(n1374) );
NAND3_X1 U1077 ( .A1(n1267), .A2(n1375), .A3(G146), .ZN(n1373) );
NAND2_X1 U1078 ( .A1(n1376), .A2(n1264), .ZN(n1372) );
INV_X1 U1079 ( .A(G146), .ZN(n1264) );
NAND2_X1 U1080 ( .A1(n1377), .A2(n1375), .ZN(n1376) );
INV_X1 U1081 ( .A(KEYINPUT7), .ZN(n1375) );
XOR2_X1 U1082 ( .A(n1267), .B(KEYINPUT27), .Z(n1377) );
XOR2_X1 U1083 ( .A(n1220), .B(n1378), .Z(n1366) );
XOR2_X1 U1084 ( .A(KEYINPUT17), .B(G227), .Z(n1378) );
XNOR2_X1 U1085 ( .A(n1103), .B(KEYINPUT0), .ZN(n1363) );
NOR2_X1 U1086 ( .A1(n1324), .A2(n1316), .ZN(n1103) );
NOR2_X1 U1087 ( .A1(n1323), .A2(G902), .ZN(n1316) );
INV_X1 U1088 ( .A(G234), .ZN(n1323) );
INV_X1 U1089 ( .A(G221), .ZN(n1324) );
AND3_X1 U1090 ( .A1(n1273), .A2(n1080), .A3(n1379), .ZN(n1250) );
NAND2_X1 U1091 ( .A1(n1380), .A2(n1104), .ZN(n1379) );
NAND3_X1 U1092 ( .A1(n1280), .A2(n1065), .A3(n1381), .ZN(n1104) );
XOR2_X1 U1093 ( .A(n1069), .B(KEYINPUT48), .Z(n1381) );
INV_X1 U1094 ( .A(G952), .ZN(n1069) );
NAND3_X1 U1095 ( .A1(G902), .A2(n1280), .A3(n1157), .ZN(n1380) );
NOR2_X1 U1096 ( .A1(n1065), .A2(G898), .ZN(n1157) );
NAND2_X1 U1097 ( .A1(G237), .A2(G234), .ZN(n1280) );
NAND2_X1 U1098 ( .A1(G214), .A2(n1382), .ZN(n1080) );
NAND3_X1 U1099 ( .A1(n1383), .A2(n1384), .A3(n1115), .ZN(n1273) );
NAND2_X1 U1100 ( .A1(n1113), .A2(n1114), .ZN(n1115) );
NAND2_X1 U1101 ( .A1(n1114), .A2(n1385), .ZN(n1384) );
OR3_X1 U1102 ( .A1(n1114), .A2(n1113), .A3(n1385), .ZN(n1383) );
INV_X1 U1103 ( .A(KEYINPUT15), .ZN(n1385) );
AND2_X1 U1104 ( .A1(n1386), .A2(n1190), .ZN(n1113) );
XOR2_X1 U1105 ( .A(n1387), .B(n1388), .Z(n1386) );
XOR2_X1 U1106 ( .A(n1225), .B(n1261), .Z(n1388) );
XOR2_X1 U1107 ( .A(n1389), .B(n1320), .Z(n1261) );
XNOR2_X1 U1108 ( .A(n1274), .B(G146), .ZN(n1320) );
INV_X1 U1109 ( .A(G128), .ZN(n1274) );
NAND2_X1 U1110 ( .A1(KEYINPUT44), .A2(n1267), .ZN(n1389) );
INV_X1 U1111 ( .A(G143), .ZN(n1267) );
XOR2_X1 U1112 ( .A(n1160), .B(n1161), .Z(n1225) );
XNOR2_X1 U1113 ( .A(n1390), .B(n1309), .ZN(n1161) );
XOR2_X1 U1114 ( .A(G113), .B(G119), .Z(n1309) );
NAND2_X1 U1115 ( .A1(KEYINPUT24), .A2(n1311), .ZN(n1390) );
INV_X1 U1116 ( .A(G116), .ZN(n1311) );
XNOR2_X1 U1117 ( .A(n1391), .B(n1392), .ZN(n1160) );
XOR2_X1 U1118 ( .A(n1393), .B(n1220), .Z(n1392) );
XNOR2_X1 U1119 ( .A(n1394), .B(n1357), .ZN(n1220) );
XOR2_X1 U1120 ( .A(G107), .B(KEYINPUT29), .Z(n1357) );
XOR2_X1 U1121 ( .A(n1276), .B(G104), .Z(n1394) );
INV_X1 U1122 ( .A(G101), .ZN(n1276) );
NOR2_X1 U1123 ( .A1(KEYINPUT61), .A2(n1395), .ZN(n1393) );
INV_X1 U1124 ( .A(G122), .ZN(n1395) );
XNOR2_X1 U1125 ( .A(G110), .B(KEYINPUT13), .ZN(n1391) );
XOR2_X1 U1126 ( .A(n1262), .B(n1255), .Z(n1387) );
AND2_X1 U1127 ( .A1(G224), .A2(n1065), .ZN(n1255) );
INV_X1 U1128 ( .A(G953), .ZN(n1065) );
INV_X1 U1129 ( .A(G125), .ZN(n1262) );
NAND2_X1 U1130 ( .A1(G210), .A2(n1382), .ZN(n1114) );
NAND2_X1 U1131 ( .A1(n1396), .A2(n1190), .ZN(n1382) );
INV_X1 U1132 ( .A(G902), .ZN(n1190) );
INV_X1 U1133 ( .A(G237), .ZN(n1396) );
endmodule


