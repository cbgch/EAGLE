//Key = 1110101010101101100110011000100111100000101001010111000000110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;

NAND2_X1 U714 ( .A1(n977), .A2(n978), .ZN(G9) );
OR2_X1 U715 ( .A1(n979), .A2(G107), .ZN(n978) );
NAND2_X1 U716 ( .A1(G107), .A2(n980), .ZN(n977) );
NAND2_X1 U717 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND2_X1 U718 ( .A1(n983), .A2(n984), .ZN(n982) );
INV_X1 U719 ( .A(KEYINPUT10), .ZN(n984) );
NAND2_X1 U720 ( .A1(KEYINPUT10), .A2(n979), .ZN(n981) );
NAND2_X1 U721 ( .A1(KEYINPUT19), .A2(n983), .ZN(n979) );
NOR2_X1 U722 ( .A1(n985), .A2(n986), .ZN(G75) );
NOR3_X1 U723 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND3_X1 U724 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n987) );
NAND2_X1 U725 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U726 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND3_X1 U727 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NAND2_X1 U728 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NAND2_X1 U729 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
OR2_X1 U730 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U731 ( .A1(n1006), .A2(n1007), .ZN(n1000) );
OR2_X1 U732 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND3_X1 U733 ( .A1(n1002), .A2(n1010), .A3(n1006), .ZN(n995) );
NAND3_X1 U734 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NAND2_X1 U735 ( .A1(n999), .A2(n1014), .ZN(n1013) );
NAND3_X1 U736 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1012) );
XOR2_X1 U737 ( .A(KEYINPUT18), .B(n999), .Z(n1016) );
NAND2_X1 U738 ( .A1(n997), .A2(n1018), .ZN(n1011) );
NAND2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
INV_X1 U741 ( .A(n1023), .ZN(n993) );
NOR3_X1 U742 ( .A1(n1024), .A2(G953), .A3(G952), .ZN(n985) );
INV_X1 U743 ( .A(n990), .ZN(n1024) );
NAND4_X1 U744 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n990) );
NOR4_X1 U745 ( .A1(n1017), .A2(n1021), .A3(n1029), .A4(n1030), .ZN(n1028) );
XOR2_X1 U746 ( .A(n1031), .B(n1032), .Z(n1029) );
NOR2_X1 U747 ( .A1(G475), .A2(KEYINPUT56), .ZN(n1032) );
NOR3_X1 U748 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1027) );
AND2_X1 U749 ( .A1(n1036), .A2(KEYINPUT13), .ZN(n1035) );
NOR2_X1 U750 ( .A1(KEYINPUT13), .A2(n1037), .ZN(n1034) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U752 ( .A(n1040), .B(n1041), .Z(n1033) );
XOR2_X1 U753 ( .A(n1042), .B(n1043), .Z(n1025) );
XNOR2_X1 U754 ( .A(KEYINPUT2), .B(KEYINPUT0), .ZN(n1042) );
XOR2_X1 U755 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U756 ( .A1(n1046), .A2(n991), .ZN(n1045) );
AND2_X1 U757 ( .A1(G227), .A2(G900), .ZN(n1046) );
NOR3_X1 U758 ( .A1(KEYINPUT60), .A2(n1047), .A3(n1048), .ZN(n1044) );
NOR2_X1 U759 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U761 ( .A(n1053), .B(KEYINPUT59), .Z(n1052) );
AND2_X1 U762 ( .A1(n1050), .A2(n1053), .ZN(n1047) );
NAND2_X1 U763 ( .A1(n991), .A2(n988), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
NAND2_X1 U765 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U766 ( .A(n1058), .B(KEYINPUT17), .Z(n1054) );
OR2_X1 U767 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
XOR2_X1 U768 ( .A(G125), .B(n1059), .Z(n1056) );
NAND2_X1 U769 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
NAND2_X1 U770 ( .A1(G131), .A2(n1062), .ZN(n1061) );
NAND2_X1 U771 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
XNOR2_X1 U772 ( .A(KEYINPUT52), .B(n1062), .ZN(n1063) );
NAND2_X1 U773 ( .A1(n1065), .A2(n1066), .ZN(G69) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U775 ( .A(n1069), .B(n1070), .Z(n1065) );
NAND2_X1 U776 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U777 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
XOR2_X1 U778 ( .A(n1076), .B(KEYINPUT29), .Z(n1075) );
NAND2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1071) );
NAND2_X1 U780 ( .A1(n1073), .A2(n1074), .ZN(n1078) );
INV_X1 U781 ( .A(n1079), .ZN(n1074) );
XNOR2_X1 U782 ( .A(n1080), .B(n1081), .ZN(n1073) );
XNOR2_X1 U783 ( .A(KEYINPUT39), .B(n1076), .ZN(n1077) );
NAND2_X1 U784 ( .A1(n991), .A2(n989), .ZN(n1076) );
OR2_X1 U785 ( .A1(n1068), .A2(n1067), .ZN(n1069) );
NAND2_X1 U786 ( .A1(G953), .A2(n1082), .ZN(n1067) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1082) );
INV_X1 U788 ( .A(KEYINPUT28), .ZN(n1068) );
NOR2_X1 U789 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U790 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U791 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U792 ( .A1(n1083), .A2(n1089), .ZN(G63) );
XOR2_X1 U793 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U794 ( .A1(n1092), .A2(n1088), .ZN(n1090) );
INV_X1 U795 ( .A(G478), .ZN(n1092) );
NOR2_X1 U796 ( .A1(n1083), .A2(n1093), .ZN(G60) );
XOR2_X1 U797 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U798 ( .A(KEYINPUT1), .B(n1096), .Z(n1095) );
NOR2_X1 U799 ( .A1(n1097), .A2(n1088), .ZN(n1096) );
INV_X1 U800 ( .A(G475), .ZN(n1097) );
NAND2_X1 U801 ( .A1(n1098), .A2(n1099), .ZN(G6) );
NAND2_X1 U802 ( .A1(G104), .A2(n1100), .ZN(n1099) );
XOR2_X1 U803 ( .A(n1101), .B(KEYINPUT11), .Z(n1098) );
OR2_X1 U804 ( .A1(n1100), .A2(G104), .ZN(n1101) );
NOR2_X1 U805 ( .A1(n1083), .A2(n1102), .ZN(G57) );
XOR2_X1 U806 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U807 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U808 ( .A(KEYINPUT46), .B(n1107), .Z(n1106) );
NOR2_X1 U809 ( .A1(KEYINPUT61), .A2(n1108), .ZN(n1107) );
NOR2_X1 U810 ( .A1(n1039), .A2(n1088), .ZN(n1105) );
INV_X1 U811 ( .A(G472), .ZN(n1039) );
XOR2_X1 U812 ( .A(n1109), .B(n1110), .Z(n1103) );
NOR2_X1 U813 ( .A1(n1083), .A2(n1111), .ZN(G54) );
XOR2_X1 U814 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U815 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U816 ( .A1(n1040), .A2(n1088), .ZN(n1114) );
INV_X1 U817 ( .A(G469), .ZN(n1040) );
XOR2_X1 U818 ( .A(n1116), .B(n1117), .Z(n1112) );
XOR2_X1 U819 ( .A(G140), .B(n1118), .Z(n1117) );
NAND2_X1 U820 ( .A1(KEYINPUT32), .A2(G110), .ZN(n1116) );
NOR2_X1 U821 ( .A1(n1083), .A2(n1119), .ZN(G51) );
XOR2_X1 U822 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U823 ( .A(KEYINPUT4), .B(n1122), .Z(n1121) );
NOR2_X1 U824 ( .A1(n1123), .A2(n1088), .ZN(n1122) );
NAND2_X1 U825 ( .A1(n1124), .A2(n1125), .ZN(n1088) );
OR2_X1 U826 ( .A1(n989), .A2(n988), .ZN(n1125) );
NAND4_X1 U827 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n988) );
AND4_X1 U828 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
AND2_X1 U829 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
OR2_X1 U830 ( .A1(n1136), .A2(n1019), .ZN(n1126) );
NAND2_X1 U831 ( .A1(n1137), .A2(n1138), .ZN(n989) );
NOR4_X1 U832 ( .A1(n1139), .A2(n1140), .A3(n983), .A4(n1141), .ZN(n1138) );
INV_X1 U833 ( .A(n1142), .ZN(n1141) );
AND3_X1 U834 ( .A1(n1005), .A2(n1002), .A3(n1143), .ZN(n983) );
AND4_X1 U835 ( .A1(n1144), .A2(n1145), .A3(n1100), .A4(n1146), .ZN(n1137) );
NAND3_X1 U836 ( .A1(n1008), .A2(n1005), .A3(n1147), .ZN(n1146) );
NAND3_X1 U837 ( .A1(n1143), .A2(n1002), .A3(n1004), .ZN(n1100) );
XOR2_X1 U838 ( .A(n1148), .B(KEYINPUT47), .Z(n1124) );
XOR2_X1 U839 ( .A(n1149), .B(n1150), .Z(n1120) );
NOR2_X1 U840 ( .A1(n991), .A2(G952), .ZN(n1083) );
NAND2_X1 U841 ( .A1(n1151), .A2(n1152), .ZN(G48) );
OR2_X1 U842 ( .A1(n1127), .A2(G146), .ZN(n1152) );
XOR2_X1 U843 ( .A(n1153), .B(KEYINPUT27), .Z(n1151) );
NAND2_X1 U844 ( .A1(G146), .A2(n1127), .ZN(n1153) );
NAND3_X1 U845 ( .A1(n1014), .A2(n1154), .A3(n1155), .ZN(n1127) );
XOR2_X1 U846 ( .A(n1156), .B(n1135), .Z(G45) );
NAND4_X1 U847 ( .A1(n1157), .A2(n1014), .A3(n1008), .A4(n1158), .ZN(n1135) );
AND3_X1 U848 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
XOR2_X1 U849 ( .A(n1059), .B(n1134), .Z(G42) );
NAND3_X1 U850 ( .A1(n1004), .A2(n1009), .A3(n1162), .ZN(n1134) );
XNOR2_X1 U851 ( .A(G137), .B(n1133), .ZN(G39) );
NAND3_X1 U852 ( .A1(n1006), .A2(n1154), .A3(n1162), .ZN(n1133) );
XOR2_X1 U853 ( .A(n1163), .B(G134), .Z(G36) );
NAND2_X1 U854 ( .A1(KEYINPUT23), .A2(n1132), .ZN(n1163) );
NAND3_X1 U855 ( .A1(n1008), .A2(n1005), .A3(n1162), .ZN(n1132) );
XOR2_X1 U856 ( .A(n1064), .B(n1131), .Z(G33) );
NAND3_X1 U857 ( .A1(n1004), .A2(n1008), .A3(n1162), .ZN(n1131) );
AND3_X1 U858 ( .A1(n1014), .A2(n1160), .A3(n999), .ZN(n1162) );
NOR2_X1 U859 ( .A1(n1043), .A2(n1021), .ZN(n999) );
INV_X1 U860 ( .A(n1022), .ZN(n1043) );
INV_X1 U861 ( .A(G131), .ZN(n1064) );
XOR2_X1 U862 ( .A(G128), .B(n1164), .Z(G30) );
NOR2_X1 U863 ( .A1(n1165), .A2(n1019), .ZN(n1164) );
INV_X1 U864 ( .A(n1157), .ZN(n1019) );
XOR2_X1 U865 ( .A(n1136), .B(KEYINPUT54), .Z(n1165) );
NAND4_X1 U866 ( .A1(n1005), .A2(n1154), .A3(n1166), .A4(n1160), .ZN(n1136) );
XOR2_X1 U867 ( .A(G101), .B(n1140), .Z(G3) );
AND3_X1 U868 ( .A1(n1008), .A2(n1143), .A3(n1006), .ZN(n1140) );
XOR2_X1 U869 ( .A(n1167), .B(n1130), .Z(G27) );
NAND3_X1 U870 ( .A1(n1009), .A2(n997), .A3(n1155), .ZN(n1130) );
AND3_X1 U871 ( .A1(n1157), .A2(n1160), .A3(n1004), .ZN(n1155) );
NAND2_X1 U872 ( .A1(n1168), .A2(n1023), .ZN(n1160) );
XOR2_X1 U873 ( .A(n1169), .B(KEYINPUT36), .Z(n1168) );
NAND3_X1 U874 ( .A1(G902), .A2(n1170), .A3(n1051), .ZN(n1169) );
NOR2_X1 U875 ( .A1(n991), .A2(G900), .ZN(n1051) );
NAND2_X1 U876 ( .A1(n1171), .A2(n1172), .ZN(G24) );
NAND2_X1 U877 ( .A1(n1139), .A2(n1173), .ZN(n1172) );
XOR2_X1 U878 ( .A(KEYINPUT12), .B(n1174), .Z(n1171) );
NOR2_X1 U879 ( .A1(n1139), .A2(n1173), .ZN(n1174) );
AND4_X1 U880 ( .A1(n1147), .A2(n1002), .A3(n1159), .A4(n1161), .ZN(n1139) );
NOR2_X1 U881 ( .A1(n1030), .A2(n1036), .ZN(n1002) );
NAND2_X1 U882 ( .A1(n1175), .A2(n1176), .ZN(G21) );
NAND2_X1 U883 ( .A1(G119), .A2(n1145), .ZN(n1176) );
XOR2_X1 U884 ( .A(KEYINPUT49), .B(n1177), .Z(n1175) );
NOR2_X1 U885 ( .A1(G119), .A2(n1145), .ZN(n1177) );
NAND3_X1 U886 ( .A1(n1147), .A2(n1154), .A3(n1006), .ZN(n1145) );
NAND2_X1 U887 ( .A1(n1178), .A2(n1179), .ZN(n1154) );
NAND3_X1 U888 ( .A1(n1036), .A2(n1030), .A3(n1180), .ZN(n1179) );
INV_X1 U889 ( .A(KEYINPUT53), .ZN(n1180) );
NAND2_X1 U890 ( .A1(KEYINPUT53), .A2(n1008), .ZN(n1178) );
XOR2_X1 U891 ( .A(n1181), .B(G116), .Z(G18) );
NAND2_X1 U892 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND4_X1 U893 ( .A1(n1005), .A2(n1184), .A3(n1147), .A4(n1185), .ZN(n1183) );
INV_X1 U894 ( .A(KEYINPUT3), .ZN(n1185) );
NAND3_X1 U895 ( .A1(n1157), .A2(n1186), .A3(KEYINPUT3), .ZN(n1182) );
NAND4_X1 U896 ( .A1(n997), .A2(n1005), .A3(n1184), .A4(n1187), .ZN(n1186) );
XOR2_X1 U897 ( .A(n1008), .B(KEYINPUT25), .Z(n1184) );
NOR2_X1 U898 ( .A1(n1159), .A2(n1026), .ZN(n1005) );
XNOR2_X1 U899 ( .A(G113), .B(n1144), .ZN(G15) );
NAND3_X1 U900 ( .A1(n1008), .A2(n1147), .A3(n1004), .ZN(n1144) );
AND2_X1 U901 ( .A1(n1026), .A2(n1159), .ZN(n1004) );
AND3_X1 U902 ( .A1(n1157), .A2(n1187), .A3(n997), .ZN(n1147) );
NOR2_X1 U903 ( .A1(n1188), .A2(n1017), .ZN(n997) );
INV_X1 U904 ( .A(n1015), .ZN(n1188) );
NOR2_X1 U905 ( .A1(n1030), .A2(n1189), .ZN(n1008) );
NAND2_X1 U906 ( .A1(n1190), .A2(n1191), .ZN(G12) );
NAND2_X1 U907 ( .A1(G110), .A2(n1142), .ZN(n1191) );
XOR2_X1 U908 ( .A(n1192), .B(KEYINPUT22), .Z(n1190) );
OR2_X1 U909 ( .A1(n1142), .A2(G110), .ZN(n1192) );
NAND3_X1 U910 ( .A1(n1006), .A2(n1143), .A3(n1009), .ZN(n1142) );
AND2_X1 U911 ( .A1(n1189), .A2(n1030), .ZN(n1009) );
XNOR2_X1 U912 ( .A(n1087), .B(n1193), .ZN(n1030) );
NOR2_X1 U913 ( .A1(n1085), .A2(G902), .ZN(n1193) );
AND2_X1 U914 ( .A1(n1194), .A2(n1195), .ZN(n1085) );
NAND2_X1 U915 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U916 ( .A(KEYINPUT16), .B(n1198), .Z(n1194) );
NOR2_X1 U917 ( .A1(n1196), .A2(n1197), .ZN(n1198) );
XNOR2_X1 U918 ( .A(n1199), .B(n1200), .ZN(n1197) );
XOR2_X1 U919 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND2_X1 U920 ( .A1(n1203), .A2(KEYINPUT6), .ZN(n1201) );
XOR2_X1 U921 ( .A(KEYINPUT43), .B(n1059), .Z(n1203) );
XOR2_X1 U922 ( .A(n1204), .B(G125), .Z(n1199) );
NAND2_X1 U923 ( .A1(n1205), .A2(KEYINPUT31), .ZN(n1204) );
XOR2_X1 U924 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U925 ( .A1(KEYINPUT62), .A2(G110), .ZN(n1207) );
XNOR2_X1 U926 ( .A(G119), .B(n1208), .ZN(n1206) );
NOR2_X1 U927 ( .A1(KEYINPUT14), .A2(n1209), .ZN(n1208) );
XOR2_X1 U928 ( .A(KEYINPUT8), .B(G128), .Z(n1209) );
XOR2_X1 U929 ( .A(n1210), .B(G137), .Z(n1196) );
NAND3_X1 U930 ( .A1(G234), .A2(n991), .A3(G221), .ZN(n1210) );
NAND2_X1 U931 ( .A1(G217), .A2(n1211), .ZN(n1087) );
INV_X1 U932 ( .A(n1036), .ZN(n1189) );
XOR2_X1 U933 ( .A(n1038), .B(G472), .Z(n1036) );
AND2_X1 U934 ( .A1(n1212), .A2(n1148), .ZN(n1038) );
XOR2_X1 U935 ( .A(n1213), .B(n1214), .Z(n1212) );
INV_X1 U936 ( .A(n1109), .ZN(n1214) );
XOR2_X1 U937 ( .A(n1215), .B(n1216), .Z(n1109) );
XOR2_X1 U938 ( .A(KEYINPUT33), .B(G113), .Z(n1216) );
XOR2_X1 U939 ( .A(n1217), .B(n1218), .Z(n1215) );
NOR2_X1 U940 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
INV_X1 U941 ( .A(G210), .ZN(n1219) );
NAND2_X1 U942 ( .A1(n1221), .A2(n1222), .ZN(n1213) );
OR2_X1 U943 ( .A1(n1110), .A2(n1108), .ZN(n1222) );
XOR2_X1 U944 ( .A(n1223), .B(KEYINPUT9), .Z(n1221) );
NAND2_X1 U945 ( .A1(n1108), .A2(n1110), .ZN(n1223) );
XOR2_X1 U946 ( .A(n1224), .B(G128), .Z(n1110) );
XNOR2_X1 U947 ( .A(G131), .B(n1225), .ZN(n1108) );
AND3_X1 U948 ( .A1(n1166), .A2(n1187), .A3(n1157), .ZN(n1143) );
NOR2_X1 U949 ( .A1(n1022), .A2(n1021), .ZN(n1157) );
AND2_X1 U950 ( .A1(G214), .A2(n1226), .ZN(n1021) );
XNOR2_X1 U951 ( .A(n1227), .B(n1123), .ZN(n1022) );
NAND2_X1 U952 ( .A1(G210), .A2(n1226), .ZN(n1123) );
NAND2_X1 U953 ( .A1(n1148), .A2(n1228), .ZN(n1226) );
NAND3_X1 U954 ( .A1(n1229), .A2(n1148), .A3(n1230), .ZN(n1227) );
NAND3_X1 U955 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
INV_X1 U956 ( .A(KEYINPUT7), .ZN(n1233) );
NAND2_X1 U957 ( .A1(KEYINPUT42), .A2(n1234), .ZN(n1232) );
OR2_X1 U958 ( .A1(n1150), .A2(n1149), .ZN(n1234) );
OR2_X1 U959 ( .A1(n1149), .A2(KEYINPUT42), .ZN(n1231) );
NAND2_X1 U960 ( .A1(n1150), .A2(n1235), .ZN(n1229) );
NAND2_X1 U961 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U962 ( .A1(KEYINPUT7), .A2(KEYINPUT42), .ZN(n1237) );
INV_X1 U963 ( .A(n1149), .ZN(n1236) );
XOR2_X1 U964 ( .A(n1238), .B(n1239), .Z(n1149) );
XOR2_X1 U965 ( .A(KEYINPUT41), .B(G128), .Z(n1239) );
XOR2_X1 U966 ( .A(n1240), .B(n1241), .Z(n1238) );
AND2_X1 U967 ( .A1(n991), .A2(G224), .ZN(n1241) );
XNOR2_X1 U968 ( .A(n1242), .B(n1081), .ZN(n1150) );
XOR2_X1 U969 ( .A(G122), .B(G110), .Z(n1081) );
NAND2_X1 U970 ( .A1(KEYINPUT40), .A2(n1080), .ZN(n1242) );
XNOR2_X1 U971 ( .A(n1243), .B(n1244), .ZN(n1080) );
XOR2_X1 U972 ( .A(G107), .B(n1245), .Z(n1244) );
NOR2_X1 U973 ( .A1(KEYINPUT57), .A2(n1246), .ZN(n1245) );
XOR2_X1 U974 ( .A(n1217), .B(n1247), .Z(n1243) );
NOR2_X1 U975 ( .A1(G113), .A2(KEYINPUT48), .ZN(n1247) );
XNOR2_X1 U976 ( .A(G101), .B(n1248), .ZN(n1217) );
XOR2_X1 U977 ( .A(G119), .B(G116), .Z(n1248) );
NAND2_X1 U978 ( .A1(n1249), .A2(n1250), .ZN(n1187) );
NAND3_X1 U979 ( .A1(n1079), .A2(n1170), .A3(G902), .ZN(n1250) );
NOR2_X1 U980 ( .A1(n991), .A2(G898), .ZN(n1079) );
XOR2_X1 U981 ( .A(n1023), .B(KEYINPUT26), .Z(n1249) );
NAND3_X1 U982 ( .A1(n1170), .A2(n991), .A3(G952), .ZN(n1023) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1170) );
XOR2_X1 U984 ( .A(n1014), .B(KEYINPUT63), .Z(n1166) );
NOR2_X1 U985 ( .A1(n1015), .A2(n1017), .ZN(n1014) );
AND2_X1 U986 ( .A1(G221), .A2(n1211), .ZN(n1017) );
NAND2_X1 U987 ( .A1(n1251), .A2(n1148), .ZN(n1211) );
XOR2_X1 U988 ( .A(KEYINPUT38), .B(G234), .Z(n1251) );
XOR2_X1 U989 ( .A(n1252), .B(G469), .Z(n1015) );
NAND2_X1 U990 ( .A1(KEYINPUT24), .A2(n1253), .ZN(n1252) );
INV_X1 U991 ( .A(n1041), .ZN(n1253) );
NAND2_X1 U992 ( .A1(n1254), .A2(n1148), .ZN(n1041) );
XOR2_X1 U993 ( .A(n1255), .B(n1115), .Z(n1254) );
XNOR2_X1 U994 ( .A(n1256), .B(n1257), .ZN(n1115) );
XNOR2_X1 U995 ( .A(n1258), .B(n1062), .ZN(n1257) );
XNOR2_X1 U996 ( .A(n1225), .B(n1259), .ZN(n1062) );
XOR2_X1 U997 ( .A(G128), .B(n1260), .Z(n1259) );
NOR2_X1 U998 ( .A1(KEYINPUT37), .A2(n1224), .ZN(n1260) );
XOR2_X1 U999 ( .A(G134), .B(G137), .Z(n1225) );
XOR2_X1 U1000 ( .A(n1261), .B(G107), .Z(n1256) );
NAND2_X1 U1001 ( .A1(KEYINPUT50), .A2(G101), .ZN(n1261) );
NAND2_X1 U1002 ( .A1(KEYINPUT20), .A2(n1262), .ZN(n1255) );
XOR2_X1 U1003 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U1004 ( .A(G110), .B(n1118), .ZN(n1264) );
AND2_X1 U1005 ( .A1(G227), .A2(n991), .ZN(n1118) );
NAND2_X1 U1006 ( .A1(KEYINPUT58), .A2(n1059), .ZN(n1263) );
INV_X1 U1007 ( .A(G140), .ZN(n1059) );
NOR2_X1 U1008 ( .A1(n1161), .A2(n1159), .ZN(n1006) );
XNOR2_X1 U1009 ( .A(n1031), .B(G475), .ZN(n1159) );
NAND2_X1 U1010 ( .A1(n1094), .A2(n1148), .ZN(n1031) );
INV_X1 U1011 ( .A(G902), .ZN(n1148) );
XOR2_X1 U1012 ( .A(n1265), .B(n1266), .Z(n1094) );
XOR2_X1 U1013 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U1014 ( .A(n1269), .B(n1270), .ZN(n1268) );
NOR2_X1 U1015 ( .A1(KEYINPUT21), .A2(n1271), .ZN(n1270) );
XOR2_X1 U1016 ( .A(KEYINPUT43), .B(G140), .Z(n1271) );
NAND2_X1 U1017 ( .A1(KEYINPUT34), .A2(n1173), .ZN(n1269) );
INV_X1 U1018 ( .A(G122), .ZN(n1173) );
XOR2_X1 U1019 ( .A(KEYINPUT35), .B(G113), .Z(n1267) );
XOR2_X1 U1020 ( .A(n1240), .B(n1272), .Z(n1265) );
XOR2_X1 U1021 ( .A(n1273), .B(n1258), .Z(n1272) );
XOR2_X1 U1022 ( .A(G131), .B(n1246), .Z(n1258) );
XOR2_X1 U1023 ( .A(G104), .B(KEYINPUT55), .Z(n1246) );
NOR2_X1 U1024 ( .A1(n1274), .A2(n1220), .ZN(n1273) );
NAND2_X1 U1025 ( .A1(n991), .A2(n1228), .ZN(n1220) );
INV_X1 U1026 ( .A(G237), .ZN(n1228) );
INV_X1 U1027 ( .A(G214), .ZN(n1274) );
XOR2_X1 U1028 ( .A(n1224), .B(n1167), .Z(n1240) );
INV_X1 U1029 ( .A(G125), .ZN(n1167) );
XOR2_X1 U1030 ( .A(n1156), .B(n1202), .Z(n1224) );
XNOR2_X1 U1031 ( .A(G146), .B(KEYINPUT51), .ZN(n1202) );
INV_X1 U1032 ( .A(G143), .ZN(n1156) );
INV_X1 U1033 ( .A(n1026), .ZN(n1161) );
XOR2_X1 U1034 ( .A(n1275), .B(G478), .Z(n1026) );
OR2_X1 U1035 ( .A1(n1091), .A2(G902), .ZN(n1275) );
XNOR2_X1 U1036 ( .A(n1276), .B(n1277), .ZN(n1091) );
XOR2_X1 U1037 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U1038 ( .A(KEYINPUT44), .B(G107), .Z(n1279) );
AND3_X1 U1039 ( .A1(n1280), .A2(G234), .A3(G217), .ZN(n1278) );
XOR2_X1 U1040 ( .A(KEYINPUT5), .B(n991), .Z(n1280) );
INV_X1 U1041 ( .A(G953), .ZN(n991) );
XNOR2_X1 U1042 ( .A(n1281), .B(n1282), .ZN(n1276) );
NAND2_X1 U1043 ( .A1(n1283), .A2(KEYINPUT15), .ZN(n1282) );
XNOR2_X1 U1044 ( .A(G128), .B(n1284), .ZN(n1283) );
XOR2_X1 U1045 ( .A(G143), .B(G134), .Z(n1284) );
NAND2_X1 U1046 ( .A1(KEYINPUT45), .A2(n1285), .ZN(n1281) );
XOR2_X1 U1047 ( .A(G116), .B(n1286), .Z(n1285) );
XOR2_X1 U1048 ( .A(KEYINPUT30), .B(G122), .Z(n1286) );
endmodule


