//Key = 1000010000010001011111101111000010100110111100110000111001100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381;

XNOR2_X1 U750 ( .A(G107), .B(n1040), .ZN(G9) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1042) );
XOR2_X1 U753 ( .A(n1046), .B(KEYINPUT48), .Z(n1044) );
NAND4_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NAND2_X1 U755 ( .A1(KEYINPUT8), .A2(n1051), .ZN(n1050) );
NAND4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1049) );
NOR4_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
NOR3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1058) );
NOR2_X1 U760 ( .A1(KEYINPUT8), .A2(n1065), .ZN(n1064) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1062) );
NOR4_X1 U765 ( .A1(n1074), .A2(n1075), .A3(n1067), .A4(n1073), .ZN(n1056) );
NOR4_X1 U766 ( .A1(n1061), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1075) );
NOR3_X1 U767 ( .A1(n1060), .A2(KEYINPUT16), .A3(n1079), .ZN(n1078) );
NOR3_X1 U768 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
XOR2_X1 U769 ( .A(KEYINPUT42), .B(n1054), .Z(n1080) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1059), .ZN(n1076) );
NOR2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
AND2_X1 U772 ( .A1(n1086), .A2(KEYINPUT18), .ZN(n1084) );
NOR3_X1 U773 ( .A1(n1052), .A2(n1087), .A3(n1088), .ZN(n1074) );
NOR3_X1 U774 ( .A1(n1089), .A2(KEYINPUT18), .A3(n1059), .ZN(n1088) );
AND3_X1 U775 ( .A1(KEYINPUT16), .A2(n1090), .A3(n1054), .ZN(n1087) );
INV_X1 U776 ( .A(n1061), .ZN(n1052) );
NOR3_X1 U777 ( .A1(n1091), .A2(n1043), .A3(n1092), .ZN(n1041) );
XOR2_X1 U778 ( .A(n1045), .B(KEYINPUT0), .Z(n1092) );
INV_X1 U779 ( .A(G952), .ZN(n1045) );
AND4_X1 U780 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1043) );
NOR4_X1 U781 ( .A1(n1097), .A2(n1098), .A3(n1059), .A4(n1099), .ZN(n1096) );
XNOR2_X1 U782 ( .A(n1100), .B(n1101), .ZN(n1098) );
NAND2_X1 U783 ( .A1(KEYINPUT11), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U784 ( .A(KEYINPUT41), .B(n1103), .ZN(n1102) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(n1097) );
XOR2_X1 U786 ( .A(KEYINPUT19), .B(n1106), .Z(n1105) );
NOR3_X1 U787 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1095) );
INV_X1 U788 ( .A(n1110), .ZN(n1107) );
NAND2_X1 U789 ( .A1(G475), .A2(n1111), .ZN(n1093) );
XOR2_X1 U790 ( .A(KEYINPUT43), .B(n1112), .Z(n1111) );
XOR2_X1 U791 ( .A(KEYINPUT55), .B(G953), .Z(n1091) );
NAND2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(G72) );
NAND2_X1 U793 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
INV_X1 U794 ( .A(n1117), .ZN(n1115) );
NAND2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
NAND2_X1 U796 ( .A1(n1119), .A2(n1116), .ZN(n1118) );
NAND2_X1 U797 ( .A1(G953), .A2(n1120), .ZN(n1116) );
INV_X1 U798 ( .A(n1121), .ZN(n1119) );
XOR2_X1 U799 ( .A(n1122), .B(n1123), .Z(n1117) );
NOR2_X1 U800 ( .A1(n1121), .A2(n1124), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U802 ( .A1(n1127), .A2(KEYINPUT57), .ZN(n1125) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1122) );
XOR2_X1 U805 ( .A(n1132), .B(n1133), .Z(G69) );
XOR2_X1 U806 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U807 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U808 ( .A(n1138), .ZN(n1137) );
NAND2_X1 U809 ( .A1(G953), .A2(n1139), .ZN(n1134) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1139) );
NOR2_X1 U811 ( .A1(n1047), .A2(G953), .ZN(n1132) );
NOR3_X1 U812 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G66) );
NOR2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U814 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR3_X1 U815 ( .A1(n1147), .A2(KEYINPUT56), .A3(KEYINPUT12), .ZN(n1146) );
AND2_X1 U816 ( .A1(n1147), .A2(KEYINPUT56), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1141) );
NOR2_X1 U818 ( .A1(KEYINPUT12), .A2(n1147), .ZN(n1148) );
OR2_X1 U819 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
XOR2_X1 U820 ( .A(KEYINPUT4), .B(n1152), .Z(n1151) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1153), .ZN(G63) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U823 ( .A1(n1156), .A2(n1150), .ZN(n1155) );
INV_X1 U824 ( .A(G478), .ZN(n1156) );
NOR2_X1 U825 ( .A1(n1140), .A2(n1157), .ZN(G60) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1160), .B(n1161), .Z(n1159) );
AND2_X1 U828 ( .A1(n1162), .A2(KEYINPUT62), .ZN(n1161) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1150), .ZN(n1160) );
NOR2_X1 U830 ( .A1(KEYINPUT62), .A2(n1162), .ZN(n1158) );
NAND3_X1 U831 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(G6) );
NAND2_X1 U832 ( .A1(G104), .A2(n1167), .ZN(n1166) );
NAND3_X1 U833 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
NAND2_X1 U834 ( .A1(KEYINPUT47), .A2(KEYINPUT44), .ZN(n1170) );
NAND2_X1 U835 ( .A1(KEYINPUT10), .A2(n1171), .ZN(n1169) );
NAND2_X1 U836 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
INV_X1 U837 ( .A(KEYINPUT10), .ZN(n1173) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1174), .ZN(n1172) );
NAND2_X1 U839 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND4_X1 U840 ( .A1(n1171), .A2(n1177), .A3(KEYINPUT47), .A4(n1175), .ZN(n1165) );
INV_X1 U841 ( .A(KEYINPUT44), .ZN(n1175) );
NAND2_X1 U842 ( .A1(KEYINPUT44), .A2(n1178), .ZN(n1164) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1179), .ZN(n1178) );
NAND2_X1 U844 ( .A1(n1177), .A2(n1176), .ZN(n1179) );
INV_X1 U845 ( .A(KEYINPUT47), .ZN(n1176) );
INV_X1 U846 ( .A(G104), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1140), .A2(n1180), .ZN(G57) );
XOR2_X1 U848 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U849 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U850 ( .A1(n1185), .A2(n1150), .ZN(n1184) );
INV_X1 U851 ( .A(G472), .ZN(n1185) );
NOR2_X1 U852 ( .A1(n1140), .A2(n1186), .ZN(G54) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U854 ( .A(n1189), .B(n1129), .Z(n1188) );
XOR2_X1 U855 ( .A(n1190), .B(n1191), .Z(n1187) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1150), .ZN(n1191) );
INV_X1 U857 ( .A(G469), .ZN(n1192) );
XNOR2_X1 U858 ( .A(KEYINPUT31), .B(KEYINPUT30), .ZN(n1190) );
NOR2_X1 U859 ( .A1(n1140), .A2(n1193), .ZN(G51) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U861 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U862 ( .A(n1198), .B(KEYINPUT52), .Z(n1197) );
NAND2_X1 U863 ( .A1(n1136), .A2(n1199), .ZN(n1198) );
NOR2_X1 U864 ( .A1(n1136), .A2(n1199), .ZN(n1196) );
NAND2_X1 U865 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
OR2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U867 ( .A1(n1101), .A2(n1150), .ZN(n1194) );
NAND2_X1 U868 ( .A1(G902), .A2(n1204), .ZN(n1150) );
NAND2_X1 U869 ( .A1(n1047), .A2(n1048), .ZN(n1204) );
INV_X1 U870 ( .A(n1131), .ZN(n1048) );
NAND4_X1 U871 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1131) );
NOR3_X1 U872 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
NOR3_X1 U873 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
XOR2_X1 U874 ( .A(n1215), .B(KEYINPUT28), .Z(n1213) );
NOR2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1209) );
NOR2_X1 U876 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NOR2_X1 U877 ( .A1(n1220), .A2(n1065), .ZN(n1219) );
NOR2_X1 U878 ( .A1(n1221), .A2(n1089), .ZN(n1218) );
NOR2_X1 U879 ( .A1(n1222), .A2(n1053), .ZN(n1221) );
NOR3_X1 U880 ( .A1(n1215), .A2(n1223), .A3(n1224), .ZN(n1222) );
AND2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1047) );
AND4_X1 U882 ( .A1(n1040), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1226) );
NAND3_X1 U883 ( .A1(n1054), .A2(n1230), .A3(n1231), .ZN(n1040) );
NOR4_X1 U884 ( .A1(n1232), .A2(n1233), .A3(n1171), .A4(n1234), .ZN(n1225) );
NOR3_X1 U885 ( .A1(n1220), .A2(n1235), .A3(n1067), .ZN(n1234) );
NOR3_X1 U886 ( .A1(n1060), .A2(n1235), .A3(n1214), .ZN(n1171) );
INV_X1 U887 ( .A(n1054), .ZN(n1060) );
NOR2_X1 U888 ( .A1(n1130), .A2(G952), .ZN(n1140) );
XOR2_X1 U889 ( .A(G146), .B(n1236), .Z(G48) );
AND2_X1 U890 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U891 ( .A(n1239), .B(n1240), .Z(G45) );
NAND4_X1 U892 ( .A1(n1241), .A2(n1069), .A3(n1242), .A4(n1243), .ZN(n1240) );
XOR2_X1 U893 ( .A(KEYINPUT6), .B(n1086), .Z(n1243) );
NOR2_X1 U894 ( .A1(n1223), .A2(n1224), .ZN(n1242) );
XOR2_X1 U895 ( .A(G140), .B(n1244), .Z(G42) );
NOR4_X1 U896 ( .A1(n1079), .A2(n1220), .A3(n1065), .A4(n1245), .ZN(n1244) );
XNOR2_X1 U897 ( .A(KEYINPUT39), .B(n1246), .ZN(n1245) );
INV_X1 U898 ( .A(n1085), .ZN(n1220) );
INV_X1 U899 ( .A(n1090), .ZN(n1079) );
NAND2_X1 U900 ( .A1(n1247), .A2(n1248), .ZN(G39) );
NAND2_X1 U901 ( .A1(n1210), .A2(n1249), .ZN(n1248) );
XOR2_X1 U902 ( .A(n1250), .B(KEYINPUT45), .Z(n1247) );
OR2_X1 U903 ( .A1(n1249), .A2(n1210), .ZN(n1250) );
NOR3_X1 U904 ( .A1(n1212), .A2(n1067), .A3(n1073), .ZN(n1210) );
INV_X1 U905 ( .A(G137), .ZN(n1249) );
NAND2_X1 U906 ( .A1(n1251), .A2(n1252), .ZN(G36) );
OR2_X1 U907 ( .A1(n1253), .A2(G134), .ZN(n1252) );
NAND2_X1 U908 ( .A1(G134), .A2(n1254), .ZN(n1251) );
NAND2_X1 U909 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
OR2_X1 U910 ( .A1(n1207), .A2(KEYINPUT63), .ZN(n1256) );
INV_X1 U911 ( .A(n1257), .ZN(n1207) );
NAND2_X1 U912 ( .A1(KEYINPUT63), .A2(n1253), .ZN(n1255) );
NAND2_X1 U913 ( .A1(KEYINPUT21), .A2(n1257), .ZN(n1253) );
NOR4_X1 U914 ( .A1(n1073), .A2(n1217), .A3(n1089), .A4(n1072), .ZN(n1257) );
XOR2_X1 U915 ( .A(G131), .B(n1258), .Z(G33) );
NOR3_X1 U916 ( .A1(n1065), .A2(n1259), .A3(n1217), .ZN(n1258) );
XOR2_X1 U917 ( .A(n1089), .B(KEYINPUT59), .Z(n1259) );
INV_X1 U918 ( .A(n1053), .ZN(n1065) );
NOR2_X1 U919 ( .A1(n1073), .A2(n1214), .ZN(n1053) );
OR2_X1 U920 ( .A1(n1070), .A2(n1108), .ZN(n1073) );
INV_X1 U921 ( .A(n1071), .ZN(n1108) );
XOR2_X1 U922 ( .A(n1205), .B(n1260), .Z(G30) );
NAND2_X1 U923 ( .A1(KEYINPUT54), .A2(G128), .ZN(n1260) );
NAND3_X1 U924 ( .A1(n1231), .A2(n1069), .A3(n1238), .ZN(n1205) );
INV_X1 U925 ( .A(n1212), .ZN(n1238) );
NAND3_X1 U926 ( .A1(n1261), .A2(n1262), .A3(n1241), .ZN(n1212) );
INV_X1 U927 ( .A(n1217), .ZN(n1241) );
NAND2_X1 U928 ( .A1(n1090), .A2(n1246), .ZN(n1217) );
XOR2_X1 U929 ( .A(G101), .B(n1233), .Z(G3) );
NOR3_X1 U930 ( .A1(n1089), .A2(n1235), .A3(n1067), .ZN(n1233) );
XOR2_X1 U931 ( .A(n1206), .B(n1263), .Z(G27) );
NAND2_X1 U932 ( .A1(KEYINPUT5), .A2(G125), .ZN(n1263) );
NAND4_X1 U933 ( .A1(n1237), .A2(n1085), .A3(n1055), .A4(n1246), .ZN(n1206) );
NAND2_X1 U934 ( .A1(n1061), .A2(n1264), .ZN(n1246) );
NAND3_X1 U935 ( .A1(G902), .A2(n1265), .A3(n1121), .ZN(n1264) );
NOR2_X1 U936 ( .A1(G900), .A2(n1130), .ZN(n1121) );
NOR2_X1 U937 ( .A1(n1214), .A2(n1215), .ZN(n1237) );
XOR2_X1 U938 ( .A(n1232), .B(n1266), .Z(G24) );
NOR2_X1 U939 ( .A1(KEYINPUT29), .A2(n1267), .ZN(n1266) );
AND4_X1 U940 ( .A1(n1268), .A2(n1054), .A3(n1269), .A4(n1270), .ZN(n1232) );
NOR2_X1 U941 ( .A1(n1099), .A2(n1262), .ZN(n1054) );
XNOR2_X1 U942 ( .A(G119), .B(n1229), .ZN(G21) );
NAND4_X1 U943 ( .A1(n1262), .A2(n1271), .A3(n1261), .A4(n1268), .ZN(n1229) );
XNOR2_X1 U944 ( .A(G116), .B(n1228), .ZN(G18) );
NAND3_X1 U945 ( .A1(n1268), .A2(n1231), .A3(n1086), .ZN(n1228) );
INV_X1 U946 ( .A(n1072), .ZN(n1231) );
NAND2_X1 U947 ( .A1(n1224), .A2(n1270), .ZN(n1072) );
NAND2_X1 U948 ( .A1(n1272), .A2(n1273), .ZN(G15) );
NAND2_X1 U949 ( .A1(G113), .A2(n1227), .ZN(n1273) );
XOR2_X1 U950 ( .A(KEYINPUT58), .B(n1274), .Z(n1272) );
NOR2_X1 U951 ( .A1(G113), .A2(n1227), .ZN(n1274) );
NAND3_X1 U952 ( .A1(n1086), .A2(n1268), .A3(n1275), .ZN(n1227) );
INV_X1 U953 ( .A(n1214), .ZN(n1275) );
NAND2_X1 U954 ( .A1(n1223), .A2(n1269), .ZN(n1214) );
AND2_X1 U955 ( .A1(n1276), .A2(n1055), .ZN(n1268) );
INV_X1 U956 ( .A(n1059), .ZN(n1055) );
INV_X1 U957 ( .A(n1089), .ZN(n1086) );
NAND2_X1 U958 ( .A1(n1261), .A2(n1277), .ZN(n1089) );
XNOR2_X1 U959 ( .A(n1099), .B(KEYINPUT20), .ZN(n1261) );
XOR2_X1 U960 ( .A(n1278), .B(n1279), .Z(G12) );
NAND3_X1 U961 ( .A1(n1230), .A2(n1280), .A3(n1271), .ZN(n1279) );
INV_X1 U962 ( .A(n1067), .ZN(n1271) );
NAND2_X1 U963 ( .A1(n1223), .A2(n1224), .ZN(n1067) );
INV_X1 U964 ( .A(n1269), .ZN(n1224) );
NAND2_X1 U965 ( .A1(n1094), .A2(n1281), .ZN(n1269) );
OR2_X1 U966 ( .A1(n1163), .A2(n1112), .ZN(n1281) );
NAND2_X1 U967 ( .A1(n1112), .A2(n1163), .ZN(n1094) );
INV_X1 U968 ( .A(G475), .ZN(n1163) );
AND2_X1 U969 ( .A1(n1162), .A2(n1282), .ZN(n1112) );
XNOR2_X1 U970 ( .A(n1283), .B(n1284), .ZN(n1162) );
XOR2_X1 U971 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U972 ( .A(n1287), .B(n1288), .ZN(n1286) );
NAND2_X1 U973 ( .A1(G214), .A2(n1289), .ZN(n1287) );
XOR2_X1 U974 ( .A(n1290), .B(n1291), .Z(n1283) );
XOR2_X1 U975 ( .A(G146), .B(G131), .Z(n1291) );
XOR2_X1 U976 ( .A(n1292), .B(G113), .Z(n1290) );
NAND2_X1 U977 ( .A1(n1293), .A2(KEYINPUT17), .ZN(n1292) );
XNOR2_X1 U978 ( .A(KEYINPUT27), .B(n1126), .ZN(n1293) );
XOR2_X1 U979 ( .A(G140), .B(G125), .Z(n1126) );
INV_X1 U980 ( .A(n1270), .ZN(n1223) );
NAND2_X1 U981 ( .A1(n1294), .A2(n1110), .ZN(n1270) );
NAND2_X1 U982 ( .A1(G478), .A2(n1295), .ZN(n1110) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1282), .ZN(n1295) );
INV_X1 U984 ( .A(n1154), .ZN(n1296) );
XNOR2_X1 U985 ( .A(n1109), .B(KEYINPUT23), .ZN(n1294) );
NOR3_X1 U986 ( .A1(G478), .A2(G902), .A3(n1154), .ZN(n1109) );
XOR2_X1 U987 ( .A(n1297), .B(n1298), .Z(n1154) );
XOR2_X1 U988 ( .A(n1285), .B(n1299), .Z(n1298) );
XNOR2_X1 U989 ( .A(n1300), .B(n1301), .ZN(n1299) );
NOR3_X1 U990 ( .A1(n1152), .A2(KEYINPUT51), .A3(n1302), .ZN(n1301) );
INV_X1 U991 ( .A(G217), .ZN(n1152) );
NOR2_X1 U992 ( .A1(KEYINPUT61), .A2(n1303), .ZN(n1300) );
XOR2_X1 U993 ( .A(KEYINPUT26), .B(G116), .Z(n1303) );
XOR2_X1 U994 ( .A(n1267), .B(G143), .Z(n1285) );
XNOR2_X1 U995 ( .A(G107), .B(n1304), .ZN(n1297) );
XOR2_X1 U996 ( .A(G134), .B(G128), .Z(n1304) );
XOR2_X1 U997 ( .A(KEYINPUT49), .B(n1085), .Z(n1280) );
NOR2_X1 U998 ( .A1(n1277), .A2(n1099), .ZN(n1085) );
XNOR2_X1 U999 ( .A(n1305), .B(G472), .ZN(n1099) );
NAND2_X1 U1000 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1001 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1002 ( .A(n1181), .B(KEYINPUT40), .Z(n1309) );
XOR2_X1 U1003 ( .A(n1310), .B(G101), .Z(n1181) );
NAND2_X1 U1004 ( .A1(G210), .A2(n1289), .ZN(n1310) );
NOR2_X1 U1005 ( .A1(G953), .A2(G237), .ZN(n1289) );
NAND2_X1 U1006 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
NAND2_X1 U1007 ( .A1(n1183), .A2(n1313), .ZN(n1312) );
INV_X1 U1008 ( .A(KEYINPUT2), .ZN(n1313) );
XOR2_X1 U1009 ( .A(n1314), .B(n1315), .Z(n1183) );
NAND3_X1 U1010 ( .A1(n1315), .A2(n1314), .A3(KEYINPUT2), .ZN(n1311) );
XOR2_X1 U1011 ( .A(n1316), .B(n1129), .Z(n1314) );
XNOR2_X1 U1012 ( .A(n1317), .B(n1318), .ZN(n1315) );
XOR2_X1 U1013 ( .A(G113), .B(n1319), .Z(n1318) );
NOR2_X1 U1014 ( .A1(G119), .A2(KEYINPUT9), .ZN(n1319) );
XOR2_X1 U1015 ( .A(n1320), .B(G116), .Z(n1317) );
XNOR2_X1 U1016 ( .A(KEYINPUT33), .B(KEYINPUT1), .ZN(n1320) );
XOR2_X1 U1017 ( .A(n1282), .B(KEYINPUT60), .Z(n1306) );
INV_X1 U1018 ( .A(n1262), .ZN(n1277) );
XOR2_X1 U1019 ( .A(n1321), .B(n1106), .Z(n1262) );
AND2_X1 U1020 ( .A1(G217), .A2(n1322), .ZN(n1106) );
NAND2_X1 U1021 ( .A1(KEYINPUT37), .A2(n1104), .ZN(n1321) );
NAND2_X1 U1022 ( .A1(n1149), .A2(n1282), .ZN(n1104) );
INV_X1 U1023 ( .A(n1143), .ZN(n1149) );
XOR2_X1 U1024 ( .A(n1323), .B(n1324), .Z(n1143) );
XOR2_X1 U1025 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1026 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1329), .ZN(n1327) );
INV_X1 U1028 ( .A(n1302), .ZN(n1329) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1130), .ZN(n1302) );
XOR2_X1 U1030 ( .A(n1330), .B(G119), .Z(n1325) );
NAND2_X1 U1031 ( .A1(KEYINPUT25), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1032 ( .A(KEYINPUT32), .B(G137), .Z(n1331) );
XOR2_X1 U1033 ( .A(n1332), .B(n1333), .Z(n1323) );
XOR2_X1 U1034 ( .A(G128), .B(G125), .Z(n1333) );
XOR2_X1 U1035 ( .A(KEYINPUT27), .B(n1334), .Z(n1332) );
INV_X1 U1036 ( .A(n1235), .ZN(n1230) );
NAND2_X1 U1037 ( .A1(n1276), .A2(n1090), .ZN(n1235) );
NAND2_X1 U1038 ( .A1(n1335), .A2(n1336), .ZN(n1090) );
OR2_X1 U1039 ( .A1(n1059), .A2(KEYINPUT15), .ZN(n1336) );
NAND2_X1 U1040 ( .A1(n1337), .A2(n1081), .ZN(n1059) );
INV_X1 U1041 ( .A(n1082), .ZN(n1337) );
NAND3_X1 U1042 ( .A1(n1082), .A2(n1081), .A3(KEYINPUT15), .ZN(n1335) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1322), .ZN(n1081) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1282), .ZN(n1322) );
XNOR2_X1 U1045 ( .A(n1338), .B(G469), .ZN(n1082) );
NAND2_X1 U1046 ( .A1(n1339), .A2(n1282), .ZN(n1338) );
XOR2_X1 U1047 ( .A(n1340), .B(n1341), .Z(n1339) );
INV_X1 U1048 ( .A(n1189), .ZN(n1341) );
XOR2_X1 U1049 ( .A(n1342), .B(n1343), .Z(n1189) );
XNOR2_X1 U1050 ( .A(n1328), .B(n1344), .ZN(n1343) );
XNOR2_X1 U1051 ( .A(n1128), .B(n1288), .ZN(n1344) );
XOR2_X1 U1052 ( .A(n1345), .B(n1346), .Z(n1128) );
NOR2_X1 U1053 ( .A1(G128), .A2(KEYINPUT13), .ZN(n1346) );
NAND2_X1 U1054 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
NAND2_X1 U1055 ( .A1(G143), .A2(n1334), .ZN(n1348) );
XOR2_X1 U1056 ( .A(n1349), .B(KEYINPUT7), .Z(n1347) );
NAND2_X1 U1057 ( .A1(G146), .A2(n1239), .ZN(n1349) );
XOR2_X1 U1058 ( .A(G140), .B(G110), .Z(n1328) );
XOR2_X1 U1059 ( .A(n1350), .B(n1351), .Z(n1342) );
XOR2_X1 U1060 ( .A(G101), .B(n1352), .Z(n1351) );
NOR2_X1 U1061 ( .A1(G953), .A2(n1120), .ZN(n1352) );
INV_X1 U1062 ( .A(G227), .ZN(n1120) );
XNOR2_X1 U1063 ( .A(G107), .B(KEYINPUT22), .ZN(n1350) );
NAND2_X1 U1064 ( .A1(KEYINPUT53), .A2(n1129), .ZN(n1340) );
XOR2_X1 U1065 ( .A(G131), .B(n1353), .Z(n1129) );
XOR2_X1 U1066 ( .A(G137), .B(G134), .Z(n1353) );
AND2_X1 U1067 ( .A1(n1069), .A2(n1354), .ZN(n1276) );
NAND2_X1 U1068 ( .A1(n1061), .A2(n1355), .ZN(n1354) );
NAND3_X1 U1069 ( .A1(G902), .A2(n1265), .A3(n1138), .ZN(n1355) );
NOR2_X1 U1070 ( .A1(n1130), .A2(G898), .ZN(n1138) );
NAND3_X1 U1071 ( .A1(n1265), .A2(n1130), .A3(G952), .ZN(n1061) );
NAND2_X1 U1072 ( .A1(G237), .A2(G234), .ZN(n1265) );
INV_X1 U1073 ( .A(n1215), .ZN(n1069) );
NAND2_X1 U1074 ( .A1(n1070), .A2(n1071), .ZN(n1215) );
NAND2_X1 U1075 ( .A1(G214), .A2(n1356), .ZN(n1071) );
XOR2_X1 U1076 ( .A(n1103), .B(n1101), .Z(n1070) );
NAND2_X1 U1077 ( .A1(G210), .A2(n1356), .ZN(n1101) );
NAND2_X1 U1078 ( .A1(n1282), .A2(n1357), .ZN(n1356) );
INV_X1 U1079 ( .A(G237), .ZN(n1357) );
NAND2_X1 U1080 ( .A1(n1358), .A2(n1282), .ZN(n1103) );
INV_X1 U1081 ( .A(G902), .ZN(n1282) );
XNOR2_X1 U1082 ( .A(n1359), .B(n1136), .ZN(n1358) );
XNOR2_X1 U1083 ( .A(n1360), .B(n1361), .ZN(n1136) );
XOR2_X1 U1084 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1085 ( .A(G113), .B(G107), .Z(n1363) );
XOR2_X1 U1086 ( .A(G119), .B(G116), .Z(n1362) );
XOR2_X1 U1087 ( .A(n1364), .B(n1365), .Z(n1360) );
NOR2_X1 U1088 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NOR2_X1 U1089 ( .A1(n1267), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1090 ( .A(KEYINPUT50), .B(G110), .Z(n1368) );
INV_X1 U1091 ( .A(G122), .ZN(n1267) );
NOR2_X1 U1092 ( .A1(G122), .A2(n1369), .ZN(n1366) );
XOR2_X1 U1093 ( .A(n1278), .B(KEYINPUT14), .Z(n1369) );
XNOR2_X1 U1094 ( .A(n1370), .B(n1371), .ZN(n1364) );
NAND2_X1 U1095 ( .A1(KEYINPUT24), .A2(n1372), .ZN(n1371) );
INV_X1 U1096 ( .A(G101), .ZN(n1372) );
NAND2_X1 U1097 ( .A1(KEYINPUT34), .A2(n1288), .ZN(n1370) );
XNOR2_X1 U1098 ( .A(G104), .B(KEYINPUT36), .ZN(n1288) );
NAND3_X1 U1099 ( .A1(n1373), .A2(n1374), .A3(n1200), .ZN(n1359) );
NAND2_X1 U1100 ( .A1(n1203), .A2(n1202), .ZN(n1200) );
OR3_X1 U1101 ( .A1(n1203), .A2(KEYINPUT3), .A3(n1202), .ZN(n1374) );
AND2_X1 U1102 ( .A1(G224), .A2(n1130), .ZN(n1203) );
INV_X1 U1103 ( .A(G953), .ZN(n1130) );
NAND2_X1 U1104 ( .A1(KEYINPUT3), .A2(n1202), .ZN(n1373) );
XOR2_X1 U1105 ( .A(n1316), .B(G125), .Z(n1202) );
NAND2_X1 U1106 ( .A1(n1375), .A2(n1376), .ZN(n1316) );
NAND2_X1 U1107 ( .A1(n1377), .A2(n1334), .ZN(n1376) );
INV_X1 U1108 ( .A(G146), .ZN(n1334) );
XOR2_X1 U1109 ( .A(KEYINPUT35), .B(n1378), .Z(n1377) );
NAND2_X1 U1110 ( .A1(n1379), .A2(G146), .ZN(n1375) );
XOR2_X1 U1111 ( .A(KEYINPUT46), .B(n1378), .Z(n1379) );
XOR2_X1 U1112 ( .A(n1380), .B(n1239), .Z(n1378) );
INV_X1 U1113 ( .A(G143), .ZN(n1239) );
NAND2_X1 U1114 ( .A1(KEYINPUT38), .A2(n1381), .ZN(n1380) );
INV_X1 U1115 ( .A(G128), .ZN(n1381) );
INV_X1 U1116 ( .A(G110), .ZN(n1278) );
endmodule


