//Key = 1011011100101001101011110000001001000110110011000110111111000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208;

XNOR2_X1 U673 ( .A(G107), .B(n916), .ZN(G9) );
NOR2_X1 U674 ( .A1(n917), .A2(n918), .ZN(G75) );
NOR4_X1 U675 ( .A1(G953), .A2(n919), .A3(n920), .A4(n921), .ZN(n918) );
NOR3_X1 U676 ( .A1(n922), .A2(n923), .A3(n924), .ZN(n920) );
NOR2_X1 U677 ( .A1(n925), .A2(n926), .ZN(n924) );
NOR3_X1 U678 ( .A1(n927), .A2(n928), .A3(n929), .ZN(n926) );
NOR2_X1 U679 ( .A1(n930), .A2(n931), .ZN(n928) );
NOR2_X1 U680 ( .A1(n932), .A2(n933), .ZN(n931) );
NOR3_X1 U681 ( .A1(n934), .A2(n935), .A3(n936), .ZN(n932) );
NOR2_X1 U682 ( .A1(n937), .A2(n938), .ZN(n936) );
NOR2_X1 U683 ( .A1(n939), .A2(n940), .ZN(n937) );
NOR2_X1 U684 ( .A1(n941), .A2(n942), .ZN(n939) );
XOR2_X1 U685 ( .A(n943), .B(KEYINPUT54), .Z(n941) );
NOR3_X1 U686 ( .A1(n944), .A2(n945), .A3(n946), .ZN(n935) );
NOR2_X1 U687 ( .A1(n947), .A2(n948), .ZN(n934) );
XOR2_X1 U688 ( .A(n945), .B(KEYINPUT8), .Z(n947) );
NOR3_X1 U689 ( .A1(n945), .A2(n949), .A3(n938), .ZN(n930) );
NOR2_X1 U690 ( .A1(n950), .A2(n951), .ZN(n949) );
XOR2_X1 U691 ( .A(KEYINPUT35), .B(n952), .Z(n951) );
NOR2_X1 U692 ( .A1(n953), .A2(n954), .ZN(n950) );
NOR4_X1 U693 ( .A1(n955), .A2(n933), .A3(n938), .A4(n945), .ZN(n925) );
INV_X1 U694 ( .A(n956), .ZN(n933) );
NOR2_X1 U695 ( .A1(n957), .A2(n958), .ZN(n955) );
NOR3_X1 U696 ( .A1(n919), .A2(G953), .A3(G952), .ZN(n917) );
AND4_X1 U697 ( .A1(n959), .A2(n960), .A3(n961), .A4(n962), .ZN(n919) );
NOR4_X1 U698 ( .A1(n963), .A2(n964), .A3(n965), .A4(n966), .ZN(n962) );
XOR2_X1 U699 ( .A(n967), .B(n968), .Z(n966) );
XOR2_X1 U700 ( .A(n969), .B(KEYINPUT52), .Z(n967) );
XOR2_X1 U701 ( .A(n970), .B(n971), .Z(n965) );
XOR2_X1 U702 ( .A(KEYINPUT45), .B(G478), .Z(n971) );
INV_X1 U703 ( .A(n944), .ZN(n964) );
INV_X1 U704 ( .A(n942), .ZN(n963) );
NOR2_X1 U705 ( .A1(n953), .A2(n972), .ZN(n961) );
XNOR2_X1 U706 ( .A(G475), .B(n973), .ZN(n972) );
XOR2_X1 U707 ( .A(n974), .B(n975), .Z(n960) );
XOR2_X1 U708 ( .A(n976), .B(KEYINPUT56), .Z(n975) );
XOR2_X1 U709 ( .A(KEYINPUT37), .B(n946), .Z(n959) );
NAND2_X1 U710 ( .A1(n977), .A2(n978), .ZN(G72) );
NAND2_X1 U711 ( .A1(n979), .A2(n980), .ZN(n978) );
XOR2_X1 U712 ( .A(n981), .B(KEYINPUT43), .Z(n977) );
OR2_X1 U713 ( .A1(n980), .A2(n979), .ZN(n981) );
NAND2_X1 U714 ( .A1(n982), .A2(n983), .ZN(n979) );
NAND2_X1 U715 ( .A1(n984), .A2(n985), .ZN(n983) );
XNOR2_X1 U716 ( .A(n986), .B(n987), .ZN(n984) );
NOR2_X1 U717 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND3_X1 U718 ( .A1(G900), .A2(n986), .A3(G953), .ZN(n982) );
XOR2_X1 U719 ( .A(n990), .B(n991), .Z(n986) );
XOR2_X1 U720 ( .A(n992), .B(KEYINPUT60), .Z(n990) );
NAND3_X1 U721 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NAND2_X1 U722 ( .A1(n996), .A2(n997), .ZN(n995) );
INV_X1 U723 ( .A(KEYINPUT16), .ZN(n997) );
NAND3_X1 U724 ( .A1(KEYINPUT16), .A2(n998), .A3(n999), .ZN(n994) );
OR2_X1 U725 ( .A1(n999), .A2(n998), .ZN(n993) );
NOR2_X1 U726 ( .A1(n1000), .A2(n996), .ZN(n998) );
INV_X1 U727 ( .A(KEYINPUT5), .ZN(n1000) );
XOR2_X1 U728 ( .A(n1001), .B(KEYINPUT6), .Z(n999) );
NAND2_X1 U729 ( .A1(n1002), .A2(n1003), .ZN(n980) );
NAND2_X1 U730 ( .A1(G900), .A2(G227), .ZN(n1003) );
INV_X1 U731 ( .A(n1004), .ZN(n1002) );
XOR2_X1 U732 ( .A(n1005), .B(n1006), .Z(G69) );
NOR2_X1 U733 ( .A1(n1007), .A2(n1004), .ZN(n1006) );
XOR2_X1 U734 ( .A(n985), .B(KEYINPUT32), .Z(n1004) );
NOR2_X1 U735 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U736 ( .A1(n1010), .A2(n1011), .ZN(n1005) );
NAND2_X1 U737 ( .A1(n1012), .A2(n985), .ZN(n1011) );
XOR2_X1 U738 ( .A(n1013), .B(n1014), .Z(n1012) );
NAND2_X1 U739 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND3_X1 U740 ( .A1(G898), .A2(n1014), .A3(G953), .ZN(n1010) );
NOR2_X1 U741 ( .A1(n1017), .A2(n1018), .ZN(G66) );
NOR3_X1 U742 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NOR2_X1 U743 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
AND3_X1 U744 ( .A1(n1023), .A2(G902), .A3(n1022), .ZN(n1020) );
NOR3_X1 U745 ( .A1(KEYINPUT1), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR2_X1 U746 ( .A1(n1017), .A2(n1026), .ZN(G63) );
XOR2_X1 U747 ( .A(n1027), .B(n1028), .Z(n1026) );
NAND3_X1 U748 ( .A1(G478), .A2(n921), .A3(n1029), .ZN(n1027) );
XOR2_X1 U749 ( .A(n1030), .B(KEYINPUT53), .Z(n1029) );
NOR2_X1 U750 ( .A1(n1017), .A2(n1031), .ZN(G60) );
XOR2_X1 U751 ( .A(n1032), .B(KEYINPUT57), .Z(n1031) );
NAND3_X1 U752 ( .A1(n1033), .A2(n1034), .A3(n973), .ZN(n1032) );
NAND2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
OR3_X1 U754 ( .A1(n1030), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U755 ( .A1(G475), .A2(n921), .ZN(n1036) );
XOR2_X1 U756 ( .A(G104), .B(n1037), .Z(G6) );
NOR2_X1 U757 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U758 ( .A1(n1017), .A2(n1040), .ZN(G57) );
XOR2_X1 U759 ( .A(n1041), .B(n1042), .Z(n1040) );
XOR2_X1 U760 ( .A(KEYINPUT44), .B(n1043), .Z(n1042) );
NOR2_X1 U761 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XOR2_X1 U762 ( .A(n1046), .B(n1047), .Z(n1045) );
NAND2_X1 U763 ( .A1(KEYINPUT12), .A2(n1048), .ZN(n1047) );
NAND3_X1 U764 ( .A1(G472), .A2(n921), .A3(G902), .ZN(n1046) );
NOR2_X1 U765 ( .A1(KEYINPUT12), .A2(n1048), .ZN(n1044) );
XNOR2_X1 U766 ( .A(n1049), .B(n1050), .ZN(n1048) );
XOR2_X1 U767 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U768 ( .A(n1053), .B(KEYINPUT40), .Z(n1049) );
NOR2_X1 U769 ( .A1(KEYINPUT59), .A2(n1054), .ZN(n1041) );
NOR2_X1 U770 ( .A1(n1017), .A2(n1055), .ZN(G54) );
XOR2_X1 U771 ( .A(n1056), .B(n1057), .Z(n1055) );
XNOR2_X1 U772 ( .A(n1058), .B(n1059), .ZN(n1057) );
XOR2_X1 U773 ( .A(n1060), .B(n1061), .Z(n1056) );
NOR2_X1 U774 ( .A1(KEYINPUT58), .A2(n1001), .ZN(n1061) );
NAND3_X1 U775 ( .A1(G902), .A2(G469), .A3(n1062), .ZN(n1060) );
XOR2_X1 U776 ( .A(n921), .B(KEYINPUT4), .Z(n1062) );
NOR2_X1 U777 ( .A1(n1017), .A2(n1063), .ZN(G51) );
XOR2_X1 U778 ( .A(n1064), .B(n1065), .Z(n1063) );
XNOR2_X1 U779 ( .A(n1066), .B(n1067), .ZN(n1065) );
NOR4_X1 U780 ( .A1(KEYINPUT62), .A2(n1024), .A3(n974), .A4(n1030), .ZN(n1067) );
INV_X1 U781 ( .A(n921), .ZN(n1024) );
NAND4_X1 U782 ( .A1(n1015), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n921) );
XNOR2_X1 U783 ( .A(KEYINPUT9), .B(n988), .ZN(n1070) );
NAND4_X1 U784 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n988) );
OR2_X1 U785 ( .A1(n1075), .A2(KEYINPUT48), .ZN(n1074) );
NAND3_X1 U786 ( .A1(n1076), .A2(n1077), .A3(KEYINPUT48), .ZN(n1073) );
NAND2_X1 U787 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND3_X1 U788 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1072) );
XOR2_X1 U789 ( .A(n945), .B(KEYINPUT38), .Z(n1082) );
NAND2_X1 U790 ( .A1(n940), .A2(n1083), .ZN(n1071) );
NAND2_X1 U791 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND3_X1 U792 ( .A1(n929), .A2(n927), .A3(n1086), .ZN(n1085) );
NAND2_X1 U793 ( .A1(n1081), .A2(n953), .ZN(n1084) );
INV_X1 U794 ( .A(n1087), .ZN(n1081) );
XNOR2_X1 U795 ( .A(KEYINPUT30), .B(n1016), .ZN(n1069) );
INV_X1 U796 ( .A(n989), .ZN(n1068) );
NAND4_X1 U797 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n989) );
AND4_X1 U798 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1015) );
AND4_X1 U799 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n916), .ZN(n1095) );
NAND4_X1 U800 ( .A1(n957), .A2(n956), .A3(n1099), .A4(n940), .ZN(n916) );
NOR2_X1 U801 ( .A1(n1100), .A2(n948), .ZN(n1099) );
NAND2_X1 U802 ( .A1(n940), .A2(n1101), .ZN(n1094) );
XNOR2_X1 U803 ( .A(KEYINPUT25), .B(n1039), .ZN(n1101) );
NAND4_X1 U804 ( .A1(n958), .A2(n956), .A3(n1102), .A4(n1103), .ZN(n1039) );
NAND2_X1 U805 ( .A1(KEYINPUT10), .A2(n1051), .ZN(n1066) );
NOR2_X1 U806 ( .A1(n985), .A2(G952), .ZN(n1017) );
XOR2_X1 U807 ( .A(G146), .B(n1104), .Z(G48) );
NOR4_X1 U808 ( .A1(KEYINPUT28), .A2(n1080), .A3(n1038), .A4(n1087), .ZN(n1104) );
XNOR2_X1 U809 ( .A(G143), .B(n1105), .ZN(G45) );
NAND4_X1 U810 ( .A1(n1106), .A2(n1086), .A3(n929), .A4(n927), .ZN(n1105) );
XOR2_X1 U811 ( .A(n1038), .B(KEYINPUT61), .Z(n1106) );
XOR2_X1 U812 ( .A(G140), .B(n1107), .Z(G42) );
NOR4_X1 U813 ( .A1(KEYINPUT13), .A2(n953), .A3(n945), .A4(n1087), .ZN(n1107) );
NAND3_X1 U814 ( .A1(n1108), .A2(n958), .A3(n1078), .ZN(n1087) );
NAND2_X1 U815 ( .A1(n1109), .A2(n1110), .ZN(G39) );
NAND2_X1 U816 ( .A1(G137), .A2(n1075), .ZN(n1110) );
XOR2_X1 U817 ( .A(n1111), .B(KEYINPUT27), .Z(n1109) );
NAND2_X1 U818 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
INV_X1 U819 ( .A(n1075), .ZN(n1113) );
NAND3_X1 U820 ( .A1(n1078), .A2(n1079), .A3(n1076), .ZN(n1075) );
XNOR2_X1 U821 ( .A(G137), .B(KEYINPUT31), .ZN(n1112) );
XNOR2_X1 U822 ( .A(G134), .B(n1088), .ZN(G36) );
NAND3_X1 U823 ( .A1(n1086), .A2(n957), .A3(n1076), .ZN(n1088) );
XNOR2_X1 U824 ( .A(G131), .B(n1089), .ZN(G33) );
NAND3_X1 U825 ( .A1(n1086), .A2(n958), .A3(n1076), .ZN(n1089) );
INV_X1 U826 ( .A(n945), .ZN(n1076) );
NAND2_X1 U827 ( .A1(n943), .A2(n942), .ZN(n945) );
AND2_X1 U828 ( .A1(n1078), .A2(n952), .ZN(n1086) );
XNOR2_X1 U829 ( .A(G128), .B(n1090), .ZN(G30) );
NAND3_X1 U830 ( .A1(n1108), .A2(n1078), .A3(n1114), .ZN(n1090) );
AND3_X1 U831 ( .A1(n957), .A2(n953), .A3(n940), .ZN(n1114) );
NOR2_X1 U832 ( .A1(n948), .A2(n1115), .ZN(n1078) );
XNOR2_X1 U833 ( .A(G101), .B(n1092), .ZN(G3) );
NAND2_X1 U834 ( .A1(n1116), .A2(n952), .ZN(n1092) );
XOR2_X1 U835 ( .A(n1117), .B(n1091), .Z(G27) );
NAND4_X1 U836 ( .A1(n1108), .A2(n1118), .A3(n958), .A4(n1119), .ZN(n1091) );
NOR3_X1 U837 ( .A1(n1038), .A2(n1115), .A3(n953), .ZN(n1119) );
AND2_X1 U838 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U839 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
INV_X1 U840 ( .A(G900), .ZN(n1123) );
INV_X1 U841 ( .A(n938), .ZN(n1118) );
XNOR2_X1 U842 ( .A(G122), .B(n1098), .ZN(G24) );
NAND4_X1 U843 ( .A1(n929), .A2(n1124), .A3(n956), .A4(n927), .ZN(n1098) );
NOR2_X1 U844 ( .A1(n1125), .A2(n953), .ZN(n956) );
INV_X1 U845 ( .A(n1080), .ZN(n953) );
XNOR2_X1 U846 ( .A(n1097), .B(n1126), .ZN(G21) );
XOR2_X1 U847 ( .A(KEYINPUT42), .B(G119), .Z(n1126) );
NAND2_X1 U848 ( .A1(n1079), .A2(n1124), .ZN(n1097) );
NOR4_X1 U849 ( .A1(n954), .A2(n927), .A3(n1080), .A4(n929), .ZN(n1079) );
INV_X1 U850 ( .A(n1108), .ZN(n954) );
XNOR2_X1 U851 ( .A(G116), .B(n1096), .ZN(G18) );
NAND3_X1 U852 ( .A1(n1124), .A2(n957), .A3(n952), .ZN(n1096) );
NOR2_X1 U853 ( .A1(n929), .A2(n1127), .ZN(n957) );
XNOR2_X1 U854 ( .A(G113), .B(n1016), .ZN(G15) );
NAND3_X1 U855 ( .A1(n952), .A2(n1124), .A3(n958), .ZN(n1016) );
AND2_X1 U856 ( .A1(n929), .A2(n1127), .ZN(n958) );
NOR3_X1 U857 ( .A1(n1038), .A2(n1100), .A3(n938), .ZN(n1124) );
NAND2_X1 U858 ( .A1(n1128), .A2(n944), .ZN(n938) );
NOR2_X1 U859 ( .A1(n1125), .A2(n1080), .ZN(n952) );
XNOR2_X1 U860 ( .A(n1093), .B(n1129), .ZN(G12) );
NOR2_X1 U861 ( .A1(KEYINPUT46), .A2(n1130), .ZN(n1129) );
INV_X1 U862 ( .A(G110), .ZN(n1130) );
NAND3_X1 U863 ( .A1(n1108), .A2(n1080), .A3(n1116), .ZN(n1093) );
AND4_X1 U864 ( .A1(n1127), .A2(n940), .A3(n1131), .A4(n1102), .ZN(n1116) );
INV_X1 U865 ( .A(n948), .ZN(n1102) );
NAND2_X1 U866 ( .A1(n946), .A2(n944), .ZN(n948) );
NAND2_X1 U867 ( .A1(G221), .A2(n1132), .ZN(n944) );
INV_X1 U868 ( .A(n1128), .ZN(n946) );
XOR2_X1 U869 ( .A(n1133), .B(G469), .Z(n1128) );
NAND2_X1 U870 ( .A1(n1134), .A2(n1030), .ZN(n1133) );
XNOR2_X1 U871 ( .A(n1001), .B(n1135), .ZN(n1134) );
XOR2_X1 U872 ( .A(n1136), .B(n1058), .Z(n1135) );
XOR2_X1 U873 ( .A(n1137), .B(n1138), .Z(n1058) );
XNOR2_X1 U874 ( .A(G107), .B(n1139), .ZN(n1138) );
NAND2_X1 U875 ( .A1(G227), .A2(n1140), .ZN(n1139) );
XOR2_X1 U876 ( .A(KEYINPUT50), .B(G953), .Z(n1140) );
XOR2_X1 U877 ( .A(n1053), .B(n1141), .Z(n1137) );
NAND2_X1 U878 ( .A1(KEYINPUT3), .A2(n1059), .ZN(n1136) );
XNOR2_X1 U879 ( .A(G110), .B(G140), .ZN(n1059) );
NOR2_X1 U880 ( .A1(n1100), .A2(n929), .ZN(n1131) );
XOR2_X1 U881 ( .A(n973), .B(n1142), .Z(n929) );
NOR2_X1 U882 ( .A1(G475), .A2(KEYINPUT47), .ZN(n1142) );
NAND2_X1 U883 ( .A1(n1035), .A2(n1030), .ZN(n973) );
XNOR2_X1 U884 ( .A(n1143), .B(n991), .ZN(n1035) );
XOR2_X1 U885 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U886 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U887 ( .A(G131), .B(G122), .Z(n1147) );
XOR2_X1 U888 ( .A(KEYINPUT26), .B(KEYINPUT20), .Z(n1146) );
XOR2_X1 U889 ( .A(n1148), .B(n1149), .Z(n1144) );
XOR2_X1 U890 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U891 ( .A(n1152), .B(G113), .Z(n1148) );
NAND2_X1 U892 ( .A1(G214), .A2(n1153), .ZN(n1152) );
INV_X1 U893 ( .A(n1103), .ZN(n1100) );
NAND2_X1 U894 ( .A1(n1120), .A2(n1154), .ZN(n1103) );
NAND2_X1 U895 ( .A1(n1122), .A2(n1009), .ZN(n1154) );
INV_X1 U896 ( .A(G898), .ZN(n1009) );
NOR3_X1 U897 ( .A1(n985), .A2(n923), .A3(n1030), .ZN(n1122) );
NAND3_X1 U898 ( .A1(n1155), .A2(n985), .A3(n1156), .ZN(n1120) );
XNOR2_X1 U899 ( .A(n923), .B(KEYINPUT17), .ZN(n1156) );
AND2_X1 U900 ( .A1(G237), .A2(G234), .ZN(n923) );
XOR2_X1 U901 ( .A(G952), .B(n922), .Z(n1155) );
INV_X1 U902 ( .A(KEYINPUT33), .ZN(n922) );
INV_X1 U903 ( .A(n1038), .ZN(n940) );
NAND2_X1 U904 ( .A1(n1157), .A2(n942), .ZN(n1038) );
NAND2_X1 U905 ( .A1(G214), .A2(n1158), .ZN(n942) );
INV_X1 U906 ( .A(n943), .ZN(n1157) );
XOR2_X1 U907 ( .A(n976), .B(n1159), .Z(n943) );
NOR2_X1 U908 ( .A1(KEYINPUT36), .A2(n974), .ZN(n1159) );
NAND2_X1 U909 ( .A1(G210), .A2(n1158), .ZN(n974) );
NAND2_X1 U910 ( .A1(n1160), .A2(n1030), .ZN(n1158) );
XOR2_X1 U911 ( .A(KEYINPUT0), .B(G237), .Z(n1160) );
NAND2_X1 U912 ( .A1(n1161), .A2(n1030), .ZN(n976) );
XNOR2_X1 U913 ( .A(n1064), .B(n1051), .ZN(n1161) );
XOR2_X1 U914 ( .A(n1014), .B(n1162), .Z(n1064) );
XOR2_X1 U915 ( .A(G125), .B(n1163), .Z(n1162) );
NOR2_X1 U916 ( .A1(G953), .A2(n1008), .ZN(n1163) );
INV_X1 U917 ( .A(G224), .ZN(n1008) );
XNOR2_X1 U918 ( .A(n1164), .B(n1165), .ZN(n1014) );
XNOR2_X1 U919 ( .A(n1141), .B(n1166), .ZN(n1165) );
XNOR2_X1 U920 ( .A(KEYINPUT63), .B(n1167), .ZN(n1166) );
NOR2_X1 U921 ( .A1(KEYINPUT34), .A2(n1168), .ZN(n1167) );
XOR2_X1 U922 ( .A(G101), .B(n1150), .Z(n1141) );
XOR2_X1 U923 ( .A(G104), .B(KEYINPUT11), .Z(n1150) );
XOR2_X1 U924 ( .A(n1169), .B(n1170), .Z(n1164) );
INV_X1 U925 ( .A(n927), .ZN(n1127) );
NAND2_X1 U926 ( .A1(n1171), .A2(n1172), .ZN(n927) );
NAND2_X1 U927 ( .A1(KEYINPUT14), .A2(n1173), .ZN(n1172) );
XOR2_X1 U928 ( .A(n970), .B(n1174), .Z(n1171) );
NOR2_X1 U929 ( .A1(KEYINPUT14), .A2(n1173), .ZN(n1174) );
XOR2_X1 U930 ( .A(KEYINPUT41), .B(G478), .Z(n1173) );
NAND2_X1 U931 ( .A1(n1175), .A2(n1030), .ZN(n970) );
XOR2_X1 U932 ( .A(KEYINPUT22), .B(n1176), .Z(n1175) );
INV_X1 U933 ( .A(n1028), .ZN(n1176) );
XOR2_X1 U934 ( .A(n1177), .B(n1178), .Z(n1028) );
XNOR2_X1 U935 ( .A(G134), .B(n1179), .ZN(n1178) );
NAND2_X1 U936 ( .A1(KEYINPUT21), .A2(n1180), .ZN(n1179) );
XOR2_X1 U937 ( .A(G143), .B(G128), .Z(n1180) );
XOR2_X1 U938 ( .A(n1169), .B(n1181), .Z(n1177) );
NOR2_X1 U939 ( .A1(n1182), .A2(KEYINPUT29), .ZN(n1181) );
NOR2_X1 U940 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U941 ( .A(KEYINPUT55), .B(G217), .Z(n1184) );
XNOR2_X1 U942 ( .A(G107), .B(n1185), .ZN(n1169) );
XOR2_X1 U943 ( .A(G122), .B(G116), .Z(n1185) );
XOR2_X1 U944 ( .A(n1186), .B(G472), .Z(n1080) );
NAND2_X1 U945 ( .A1(n1187), .A2(n1030), .ZN(n1186) );
XOR2_X1 U946 ( .A(n1188), .B(n1189), .Z(n1187) );
XNOR2_X1 U947 ( .A(n1054), .B(n1052), .ZN(n1189) );
XOR2_X1 U948 ( .A(n1190), .B(n1168), .Z(n1052) );
XNOR2_X1 U949 ( .A(G113), .B(KEYINPUT2), .ZN(n1168) );
NAND2_X1 U950 ( .A1(KEYINPUT18), .A2(n1191), .ZN(n1190) );
XOR2_X1 U951 ( .A(G119), .B(G116), .Z(n1191) );
XOR2_X1 U952 ( .A(n1192), .B(G101), .Z(n1054) );
NAND2_X1 U953 ( .A1(G210), .A2(n1153), .ZN(n1192) );
NOR2_X1 U954 ( .A1(G953), .A2(G237), .ZN(n1153) );
XOR2_X1 U955 ( .A(n1193), .B(KEYINPUT51), .Z(n1188) );
NAND2_X1 U956 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U957 ( .A1(n1053), .A2(n1051), .ZN(n1195) );
XOR2_X1 U958 ( .A(n1196), .B(KEYINPUT39), .Z(n1194) );
OR2_X1 U959 ( .A1(n1051), .A2(n1053), .ZN(n1196) );
XNOR2_X1 U960 ( .A(n996), .B(KEYINPUT49), .ZN(n1053) );
XOR2_X1 U961 ( .A(G131), .B(n1197), .Z(n996) );
XOR2_X1 U962 ( .A(G137), .B(G134), .Z(n1197) );
XNOR2_X1 U963 ( .A(n1001), .B(KEYINPUT19), .ZN(n1051) );
XNOR2_X1 U964 ( .A(G128), .B(n1151), .ZN(n1001) );
XOR2_X1 U965 ( .A(G143), .B(G146), .Z(n1151) );
XOR2_X1 U966 ( .A(n1125), .B(KEYINPUT24), .Z(n1108) );
NAND2_X1 U967 ( .A1(n1198), .A2(n1199), .ZN(n1125) );
NAND2_X1 U968 ( .A1(n968), .A2(n969), .ZN(n1199) );
XOR2_X1 U969 ( .A(KEYINPUT23), .B(n1200), .Z(n1198) );
NOR2_X1 U970 ( .A1(n968), .A2(n969), .ZN(n1200) );
INV_X1 U971 ( .A(n1019), .ZN(n969) );
NOR2_X1 U972 ( .A1(n1023), .A2(G902), .ZN(n1019) );
XOR2_X1 U973 ( .A(n1201), .B(n1202), .Z(n1023) );
XOR2_X1 U974 ( .A(n1203), .B(n991), .Z(n1202) );
XOR2_X1 U975 ( .A(n1117), .B(G140), .Z(n991) );
INV_X1 U976 ( .A(G125), .ZN(n1117) );
NAND2_X1 U977 ( .A1(KEYINPUT7), .A2(n1204), .ZN(n1203) );
XOR2_X1 U978 ( .A(G128), .B(n1170), .Z(n1204) );
XOR2_X1 U979 ( .A(G110), .B(G119), .Z(n1170) );
XOR2_X1 U980 ( .A(n1205), .B(n1206), .Z(n1201) );
XOR2_X1 U981 ( .A(G146), .B(G137), .Z(n1206) );
NAND2_X1 U982 ( .A1(G221), .A2(n1207), .ZN(n1205) );
INV_X1 U983 ( .A(n1183), .ZN(n1207) );
NAND2_X1 U984 ( .A1(G234), .A2(n985), .ZN(n1183) );
INV_X1 U985 ( .A(G953), .ZN(n985) );
INV_X1 U986 ( .A(n1025), .ZN(n968) );
NAND2_X1 U987 ( .A1(G217), .A2(n1132), .ZN(n1025) );
NAND2_X1 U988 ( .A1(n1208), .A2(n1030), .ZN(n1132) );
INV_X1 U989 ( .A(G902), .ZN(n1030) );
XNOR2_X1 U990 ( .A(G234), .B(KEYINPUT15), .ZN(n1208) );
endmodule


