//Key = 0000000000000001000000000000001000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000
module c5315 ( G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, 
        G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, 
        G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, 
        G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, 
        G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, 
        G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, 
        G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, 
        G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, 
        G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, 
        G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, 
        G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, 
        G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, 
        G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, 
        G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, 
        G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, 
        KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, 
        KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, 
        KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, 
        KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, 
        KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, 
        KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, 
        KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, 
        KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, 
        KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, 
        KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, 
        KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65, 
        KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71, 
        KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77, 
        KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83, 
        KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89, 
        KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95, 
        KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100, 
        KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105, 
        KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110, 
        KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115, 
        KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120, 
        KEYINPUT121, KEYINPUT122, KEYINPUT123, G144, G298, G973, G594, G599, 
        G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, 
        G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, 
        G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, 
        G707, G715, G598_enc, G610_enc, G588_enc, G615_enc, G626_enc, G632_enc,  G1002, G1004, 
        G591, G618, G621, G629, G822, G838, G861, G623, G722,         
        G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575_enc,         
        G585_enc, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,  G642, G664, 
        G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,         
        G828, G830, G854_enc, G863, G865, G867, G869, G712, G727, G732, G737,  
        G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688,  
        G843, G882, G767, G807, G658, G690 );
  input G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
         G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
         G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
         G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
         G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136,
         G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164,
         G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197,
         G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234,
         G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273,
         G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315,
         G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358,
         G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422,
         G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545,
         G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694,
         G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724,
         G4087, G4088, G4089, G4090, G4091, G4092, G4115, KEYINPUT0, KEYINPUT1,
         KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
         KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
         KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
         KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
         KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
         KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33,
         KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
         KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
         KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
         KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
         KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
         KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63,
         KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
         KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73,
         KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78,
         KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
         KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
         KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
         KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
         KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
         KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
         KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
         KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
         KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123;
         
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
         G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926,
         G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939,
         G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598_enc,
         G610_enc, G588_enc, G615_enc, G626_enc, G632_enc, G1002, G1004, G591, 
         G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836,         
         G859, G871, G873, G875, G877, G998, G1000, G575_enc, G585_enc, G661, 
         G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667,
          G670, G676, G696, G699, G702, G818, G813, G824, G826, G828,         
          G830, G854_enc, G863, G865, G867, G869, G712, G727, G732, G737, G742, 
          G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, 
          G882, G767, G807, G658, G690;
  wire   n3379, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486;

  NOR3_X2 U2403 ( .A1(n3647), .A2(G1689), .A3(n3744), .ZN(n3687) );
  NOR3_X2 U2404 ( .A1(n3647), .A2(G1691), .A3(n3619), .ZN(n3596) );
  NOR3_X2 U2405 ( .A1(n3747), .A2(n3647), .A3(n3744), .ZN(n3688) );
  NOR2_X2 U2406 ( .A1(n3395), .A2(G4091), .ZN(n3680) );
  NOR3_X2 U2407 ( .A1(n3623), .A2(n3647), .A3(n3619), .ZN(n3597) );
  NOR2_X2 U2408 ( .A1(G4091), .A2(G4092), .ZN(n3396) );
  BUF_X1 U2409 ( .A(G293), .Z(G298) );
  BUF_X1 U2410 ( .A(G3173), .Z(G973) );
  BUF_X1 U2411 ( .A(G594), .Z(G604) );
  BUF_X1 U2412 ( .A(G594), .Z(G603) );
  BUF_X1 U2413 ( .A(G137), .Z(G926) );
  BUF_X1 U2414 ( .A(G141), .Z(G923) );
  BUF_X1 U2415 ( .A(G141), .Z(G144) );
  BUF_X1 U2416 ( .A(G549), .Z(G892) );
  INV_X1 U2417 ( .A(G1), .ZN(n3379) );
  INV_X1 U2418 ( .A(n3379), .ZN(G939) );
  INV_X1 U2419 ( .A(n3379), .ZN(G921) );
  INV_X1 U2420 ( .A(n3379), .ZN(G949) );
  INV_X1 U2421 ( .A(n3379), .ZN(G993) );
  INV_X1 U2422 ( .A(n3379), .ZN(G978) );
  BUF_X1 U2423 ( .A(G299), .Z(G889) );
  BUF_X1 U2424 ( .A(G299), .Z(G887) );
  BUF_X1 U2425 ( .A(G717), .Z(G704) );
  BUF_X1 U2426 ( .A(G606), .Z(G602) );
  NAND3_X1 U2427 ( .A1(n3389), .A2(n3390), .A3(n3391), .ZN(G882) );
  NAND2_X1 U2428 ( .A1(G4092), .A2(G118), .ZN(n3391) );
  NAND2_X1 U2429 ( .A1(G4091), .A2(n3392), .ZN(n3390) );
  NAND3_X1 U2430 ( .A1(n3393), .A2(n3394), .A3(n3395), .ZN(n3392) );
  NAND2_X1 U2431 ( .A1(n3396), .A2(n3397), .ZN(n3389) );
  INV_X1 U2432 ( .A(n3398), .ZN(G865) );
  INV_X1 U2433 ( .A(n3399), .ZN(G861) );
  NAND4_X1 U2434 ( .A1(n3400), .A2(n3401), .A3(n3402), .A4(n3403), .ZN(G859) );
  NAND2_X1 U2435 ( .A1(n3404), .A2(n3399), .ZN(n3403) );
  NAND2_X1 U2436 ( .A1(n3405), .A2(n3406), .ZN(n3402) );
  NAND2_X1 U2437 ( .A1(G11), .A2(n3407), .ZN(n3401) );
  NAND2_X1 U2438 ( .A1(G61), .A2(n3408), .ZN(n3400) );
  OR2_X1 U2439 ( .A1(n3409), .A2(KEYINPUT6), .ZN(G854_enc) );
  NOR3_X1 U2440 ( .A1(n3410), .A2(G848), .A3(n3411), .ZN(n3409) );
  NOR2_X1 U2441 ( .A1(KEYINPUT68), .A2(n3412), .ZN(n3411) );
  NOR3_X1 U2442 ( .A1(n3413), .A2(G1000), .A3(G1002), .ZN(n3412) );
  OR3_X1 U2443 ( .A1(G998), .A2(G850), .A3(G1004), .ZN(n3413) );
  XNOR2_X1 U2444 ( .A(n3414), .B(n3415), .ZN(G998) );
  XOR2_X1 U2445 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR2_X1 U2446 ( .A(n3418), .B(n3419), .Z(n3417) );
  NAND2_X1 U2447 ( .A1(n3420), .A2(n3421), .ZN(n3419) );
  NAND2_X1 U2448 ( .A1(n3422), .A2(n3423), .ZN(n3421) );
  XNOR2_X1 U2449 ( .A(n3424), .B(G369), .ZN(n3422) );
  NAND2_X1 U2450 ( .A1(n3425), .A2(G332), .ZN(n3420) );
  XNOR2_X1 U2451 ( .A(n3424), .B(G372), .ZN(n3425) );
  XNOR2_X1 U2452 ( .A(n3426), .B(n3427), .ZN(n3416) );
  XOR2_X1 U2453 ( .A(n3428), .B(n3429), .Z(n3414) );
  XOR2_X1 U2454 ( .A(n3430), .B(n3431), .Z(n3429) );
  XNOR2_X1 U2455 ( .A(n3432), .B(n3433), .ZN(n3428) );
  NOR2_X1 U2456 ( .A1(n3434), .A2(KEYINPUT77), .ZN(n3410) );
  NOR3_X1 U2457 ( .A1(G847), .A2(G851), .A3(G849), .ZN(n3434) );
  INV_X1 U2458 ( .A(G559), .ZN(G851) );
  INV_X1 U2459 ( .A(G245), .ZN(G848) );
  NAND2_X1 U2460 ( .A1(G556), .A2(G386), .ZN(G847) );
  NAND2_X1 U2461 ( .A1(n3435), .A2(G27), .ZN(G845) );
  INV_X1 U2462 ( .A(G2824), .ZN(n3435) );
  NAND3_X1 U2463 ( .A1(n3436), .A2(n3437), .A3(n3438), .ZN(G843) );
  NAND2_X1 U2464 ( .A1(G120), .A2(G4092), .ZN(n3438) );
  NAND2_X1 U2465 ( .A1(G4091), .A2(n3439), .ZN(n3437) );
  NAND3_X1 U2466 ( .A1(n3440), .A2(n3441), .A3(n3395), .ZN(n3439) );
  NAND2_X1 U2467 ( .A1(n3396), .A2(n3442), .ZN(n3436) );
  INV_X1 U2468 ( .A(n3443), .ZN(G826) );
  INV_X1 U2469 ( .A(n3406), .ZN(G822) );
  NAND2_X1 U2470 ( .A1(G83), .A2(n3444), .ZN(G820) );
  AND3_X1 U2471 ( .A1(n3445), .A2(n3446), .A3(n3447), .ZN(G818) );
  NAND2_X1 U2472 ( .A1(G4115), .A2(G135), .ZN(n3447) );
  NAND2_X1 U2473 ( .A1(n3448), .A2(n3449), .ZN(n3446) );
  INV_X1 U2474 ( .A(G3724), .ZN(n3449) );
  NAND2_X1 U2475 ( .A1(n3450), .A2(n3451), .ZN(n3448) );
  OR2_X1 U2476 ( .A1(n3452), .A2(G123), .ZN(n3451) );
  OR2_X1 U2477 ( .A1(n3453), .A2(G3717), .ZN(n3450) );
  NAND2_X1 U2478 ( .A1(G3724), .A2(n3454), .ZN(n3445) );
  NAND2_X1 U2479 ( .A1(n3455), .A2(n3456), .ZN(n3454) );
  NAND2_X1 U2480 ( .A1(G3717), .A2(G623), .ZN(n3456) );
  NAND2_X1 U2481 ( .A1(n3457), .A2(n3452), .ZN(n3455) );
  INV_X1 U2482 ( .A(G3717), .ZN(n3452) );
  XOR2_X1 U2483 ( .A(n3458), .B(G132), .Z(n3457) );
  NOR2_X1 U2484 ( .A1(G3173), .A2(n3459), .ZN(G815) );
  INV_X1 U2485 ( .A(G136), .ZN(n3459) );
  XNOR2_X1 U2486 ( .A(G132), .B(n3460), .ZN(G813) );
  AND2_X1 U2487 ( .A1(G141), .A2(G145), .ZN(G810) );
  NAND4_X1 U2488 ( .A1(n3461), .A2(n3462), .A3(n3463), .A4(n3464), .ZN(G807) );
  NAND2_X1 U2489 ( .A1(n3404), .A2(n3465), .ZN(n3464) );
  NAND2_X1 U2490 ( .A1(n3405), .A2(n3466), .ZN(n3463) );
  NAND2_X1 U2491 ( .A1(G14), .A2(n3407), .ZN(n3462) );
  NAND2_X1 U2492 ( .A1(G64), .A2(n3408), .ZN(n3461) );
  NAND4_X1 U2493 ( .A1(n3467), .A2(n3468), .A3(n3469), .A4(n3470), .ZN(G802) );
  NAND2_X1 U2494 ( .A1(n3405), .A2(n3471), .ZN(n3470) );
  NOR2_X1 U2495 ( .A1(KEYINPUT108), .A2(n3472), .ZN(n3469) );
  NOR2_X1 U2496 ( .A1(G877), .A2(n3473), .ZN(n3472) );
  NAND2_X1 U2497 ( .A1(G67), .A2(n3407), .ZN(n3468) );
  NAND2_X1 U2498 ( .A1(G70), .A2(n3408), .ZN(n3467) );
  NAND4_X1 U2499 ( .A1(n3474), .A2(n3475), .A3(n3476), .A4(n3477), .ZN(G797) );
  NAND2_X1 U2500 ( .A1(n3405), .A2(n3478), .ZN(n3477) );
  NOR2_X1 U2501 ( .A1(KEYINPUT116), .A2(n3479), .ZN(n3476) );
  NOR2_X1 U2502 ( .A1(G875), .A2(n3473), .ZN(n3479) );
  NAND2_X1 U2503 ( .A1(G73), .A2(n3407), .ZN(n3475) );
  NAND2_X1 U2504 ( .A1(G17), .A2(n3408), .ZN(n3474) );
  NAND3_X1 U2505 ( .A1(n3480), .A2(n3481), .A3(n3482), .ZN(G792) );
  NOR3_X1 U2506 ( .A1(n3483), .A2(KEYINPUT120), .A3(n3484), .ZN(n3482) );
  NOR2_X1 U2507 ( .A1(G873), .A2(n3473), .ZN(n3484) );
  NOR2_X1 U2508 ( .A1(G834), .A2(n3485), .ZN(n3483) );
  INV_X1 U2509 ( .A(n3405), .ZN(n3485) );
  NAND2_X1 U2510 ( .A1(G76), .A2(n3407), .ZN(n3481) );
  NAND2_X1 U2511 ( .A1(G20), .A2(n3408), .ZN(n3480) );
  NAND4_X1 U2512 ( .A1(n3486), .A2(n3487), .A3(n3488), .A4(n3489), .ZN(G787) );
  NAND2_X1 U2513 ( .A1(n3404), .A2(n3490), .ZN(n3489) );
  NAND2_X1 U2514 ( .A1(n3405), .A2(n3491), .ZN(n3488) );
  NAND2_X1 U2515 ( .A1(G43), .A2(n3407), .ZN(n3487) );
  NAND2_X1 U2516 ( .A1(G37), .A2(n3408), .ZN(n3486) );
  NAND4_X1 U2517 ( .A1(n3492), .A2(n3493), .A3(n3494), .A4(n3495), .ZN(G782) );
  NAND2_X1 U2518 ( .A1(n3405), .A2(n3496), .ZN(n3495) );
  NOR2_X1 U2519 ( .A1(KEYINPUT110), .A2(n3497), .ZN(n3494) );
  NOR2_X1 U2520 ( .A1(G869), .A2(n3473), .ZN(n3497) );
  NAND2_X1 U2521 ( .A1(G91), .A2(n3407), .ZN(n3493) );
  NAND2_X1 U2522 ( .A1(G40), .A2(n3408), .ZN(n3492) );
  NAND4_X1 U2523 ( .A1(n3498), .A2(n3499), .A3(n3500), .A4(n3501), .ZN(G777) );
  NOR3_X1 U2524 ( .A1(n3502), .A2(KEYINPUT98), .A3(KEYINPUT102), .ZN(n3501) );
  NOR2_X1 U2525 ( .A1(G867), .A2(n3473), .ZN(n3502) );
  INV_X1 U2526 ( .A(n3503), .ZN(G867) );
  NAND2_X1 U2527 ( .A1(G103), .A2(n3408), .ZN(n3500) );
  NAND2_X1 U2528 ( .A1(n3405), .A2(n3504), .ZN(n3499) );
  NAND2_X1 U2529 ( .A1(G100), .A2(n3407), .ZN(n3498) );
  NAND4_X1 U2530 ( .A1(n3505), .A2(n3506), .A3(n3507), .A4(n3508), .ZN(G772) );
  NAND2_X1 U2531 ( .A1(n3404), .A2(n3398), .ZN(n3508) );
  NAND2_X1 U2532 ( .A1(n3405), .A2(n3443), .ZN(n3507) );
  NAND2_X1 U2533 ( .A1(G46), .A2(n3407), .ZN(n3506) );
  NAND2_X1 U2534 ( .A1(G49), .A2(n3408), .ZN(n3505) );
  NAND4_X1 U2535 ( .A1(n3509), .A2(n3510), .A3(n3511), .A4(n3512), .ZN(G767) );
  NAND2_X1 U2536 ( .A1(n3513), .A2(n3466), .ZN(n3512) );
  NAND2_X1 U2537 ( .A1(n3514), .A2(G14), .ZN(n3511) );
  NAND2_X1 U2538 ( .A1(n3515), .A2(n3465), .ZN(n3510) );
  NAND2_X1 U2539 ( .A1(n3516), .A2(G64), .ZN(n3509) );
  NAND3_X1 U2540 ( .A1(n3517), .A2(n3518), .A3(n3519), .ZN(G762) );
  NOR3_X1 U2541 ( .A1(n3520), .A2(KEYINPUT107), .A3(n3521), .ZN(n3519) );
  NOR2_X1 U2542 ( .A1(G838), .A2(n3522), .ZN(n3521) );
  AND2_X1 U2543 ( .A1(G67), .A2(n3514), .ZN(n3520) );
  NAND2_X1 U2544 ( .A1(n3515), .A2(n3523), .ZN(n3518) );
  NAND2_X1 U2545 ( .A1(n3516), .A2(G70), .ZN(n3517) );
  NAND4_X1 U2546 ( .A1(n3524), .A2(n3525), .A3(n3526), .A4(n3527), .ZN(G757) );
  NAND2_X1 U2547 ( .A1(n3514), .A2(G73), .ZN(n3527) );
  NOR2_X1 U2548 ( .A1(KEYINPUT115), .A2(n3528), .ZN(n3526) );
  NOR2_X1 U2549 ( .A1(G836), .A2(n3522), .ZN(n3528) );
  NAND2_X1 U2550 ( .A1(n3515), .A2(n3529), .ZN(n3525) );
  NAND2_X1 U2551 ( .A1(n3516), .A2(G17), .ZN(n3524) );
  NAND3_X1 U2552 ( .A1(n3530), .A2(n3531), .A3(n3532), .ZN(G752) );
  NOR3_X1 U2553 ( .A1(n3533), .A2(KEYINPUT119), .A3(n3534), .ZN(n3532) );
  NOR2_X1 U2554 ( .A1(G834), .A2(n3522), .ZN(n3534) );
  AND2_X1 U2555 ( .A1(G76), .A2(n3514), .ZN(n3533) );
  NAND2_X1 U2556 ( .A1(n3515), .A2(n3535), .ZN(n3531) );
  NAND2_X1 U2557 ( .A1(n3516), .A2(G20), .ZN(n3530) );
  NAND4_X1 U2558 ( .A1(n3536), .A2(n3537), .A3(n3538), .A4(n3539), .ZN(G747) );
  NAND2_X1 U2559 ( .A1(n3514), .A2(G43), .ZN(n3539) );
  NOR2_X1 U2560 ( .A1(KEYINPUT123), .A2(n3540), .ZN(n3538) );
  NOR2_X1 U2561 ( .A1(G832), .A2(n3522), .ZN(n3540) );
  NAND2_X1 U2562 ( .A1(n3515), .A2(n3490), .ZN(n3537) );
  NAND2_X1 U2563 ( .A1(n3516), .A2(G37), .ZN(n3536) );
  NAND4_X1 U2564 ( .A1(n3541), .A2(n3542), .A3(n3543), .A4(n3544), .ZN(G742) );
  NAND2_X1 U2565 ( .A1(n3514), .A2(G91), .ZN(n3544) );
  NOR2_X1 U2566 ( .A1(KEYINPUT109), .A2(n3545), .ZN(n3543) );
  NOR2_X1 U2567 ( .A1(G830), .A2(n3522), .ZN(n3545) );
  NAND2_X1 U2568 ( .A1(n3515), .A2(n3546), .ZN(n3542) );
  NAND2_X1 U2569 ( .A1(n3516), .A2(G40), .ZN(n3541) );
  NAND4_X1 U2570 ( .A1(n3547), .A2(n3548), .A3(n3549), .A4(n3550), .ZN(G737) );
  NOR3_X1 U2571 ( .A1(n3551), .A2(KEYINPUT97), .A3(KEYINPUT101), .ZN(n3550) );
  NOR2_X1 U2572 ( .A1(G828), .A2(n3522), .ZN(n3551) );
  NAND2_X1 U2573 ( .A1(n3516), .A2(G103), .ZN(n3549) );
  NAND2_X1 U2574 ( .A1(n3514), .A2(G100), .ZN(n3548) );
  NAND2_X1 U2575 ( .A1(n3515), .A2(n3503), .ZN(n3547) );
  NAND4_X1 U2576 ( .A1(n3552), .A2(n3553), .A3(n3554), .A4(n3555), .ZN(G732) );
  NAND2_X1 U2577 ( .A1(n3513), .A2(n3443), .ZN(n3555) );
  NAND2_X1 U2578 ( .A1(n3514), .A2(G46), .ZN(n3554) );
  NAND2_X1 U2579 ( .A1(n3515), .A2(n3398), .ZN(n3553) );
  NAND2_X1 U2580 ( .A1(n3516), .A2(G49), .ZN(n3552) );
  NAND4_X1 U2581 ( .A1(n3556), .A2(n3557), .A3(n3558), .A4(n3559), .ZN(G727) );
  NAND2_X1 U2582 ( .A1(G109), .A2(n3514), .ZN(n3559) );
  NOR2_X1 U2583 ( .A1(KEYINPUT91), .A2(n3560), .ZN(n3558) );
  NOR2_X1 U2584 ( .A1(G824), .A2(n3522), .ZN(n3560) );
  INV_X1 U2585 ( .A(n3513), .ZN(n3522) );
  NAND2_X1 U2586 ( .A1(n3515), .A2(n3561), .ZN(n3557) );
  NAND2_X1 U2587 ( .A1(G106), .A2(n3516), .ZN(n3556) );
  NAND4_X1 U2588 ( .A1(n3562), .A2(n3563), .A3(n3564), .A4(n3565), .ZN(G722) );
  NAND2_X1 U2589 ( .A1(n3513), .A2(n3406), .ZN(n3565) );
  NOR2_X1 U2590 ( .A1(G4087), .A2(G4088), .ZN(n3513) );
  NAND2_X1 U2591 ( .A1(n3514), .A2(G11), .ZN(n3564) );
  NOR2_X1 U2592 ( .A1(n3566), .A2(G4088), .ZN(n3514) );
  NAND2_X1 U2593 ( .A1(n3515), .A2(n3399), .ZN(n3563) );
  NOR2_X1 U2594 ( .A1(n3567), .A2(G4087), .ZN(n3515) );
  NAND2_X1 U2595 ( .A1(n3516), .A2(G61), .ZN(n3562) );
  NOR2_X1 U2596 ( .A1(n3567), .A2(n3566), .ZN(n3516) );
  INV_X1 U2597 ( .A(G4087), .ZN(n3566) );
  INV_X1 U2598 ( .A(G4088), .ZN(n3567) );
  OR3_X1 U2599 ( .A1(n3568), .A2(n3569), .A3(G809), .ZN(G717) );
  NOR2_X1 U2600 ( .A1(G88), .A2(G2358), .ZN(n3569) );
  NOR2_X1 U2601 ( .A1(G34), .A2(n3570), .ZN(n3568) );
  NOR2_X1 U2602 ( .A1(n3571), .A2(n3572), .ZN(G715) );
  NOR3_X1 U2603 ( .A1(n3573), .A2(KEYINPUT87), .A3(KEYINPUT86), .ZN(n3571) );
  NAND3_X1 U2604 ( .A1(n3574), .A2(n3575), .A3(n3444), .ZN(n3573) );
  NAND2_X1 U2605 ( .A1(G82), .A2(n3570), .ZN(n3575) );
  NAND2_X1 U2606 ( .A1(G80), .A2(G2358), .ZN(n3574) );
  NAND4_X1 U2607 ( .A1(n3576), .A2(n3577), .A3(n3578), .A4(n3579), .ZN(G712) );
  NAND2_X1 U2608 ( .A1(n3405), .A2(n3580), .ZN(n3579) );
  NOR2_X1 U2609 ( .A1(G4089), .A2(G4090), .ZN(n3405) );
  NOR2_X1 U2610 ( .A1(KEYINPUT94), .A2(n3581), .ZN(n3578) );
  NOR2_X1 U2611 ( .A1(G863), .A2(n3473), .ZN(n3581) );
  INV_X1 U2612 ( .A(n3404), .ZN(n3473) );
  NOR2_X1 U2613 ( .A1(n3582), .A2(G4090), .ZN(n3404) );
  NAND2_X1 U2614 ( .A1(G109), .A2(n3407), .ZN(n3577) );
  NOR2_X1 U2615 ( .A1(n3583), .A2(G4089), .ZN(n3407) );
  NAND2_X1 U2616 ( .A1(G106), .A2(n3408), .ZN(n3576) );
  NOR2_X1 U2617 ( .A1(n3583), .A2(n3582), .ZN(n3408) );
  INV_X1 U2618 ( .A(G4089), .ZN(n3582) );
  INV_X1 U2619 ( .A(G4090), .ZN(n3583) );
  NOR2_X1 U2620 ( .A1(n3584), .A2(n3572), .ZN(G707) );
  NOR3_X1 U2621 ( .A1(n3585), .A2(KEYINPUT85), .A3(KEYINPUT84), .ZN(n3584) );
  NAND3_X1 U2622 ( .A1(n3586), .A2(n3587), .A3(n3444), .ZN(n3585) );
  NAND2_X1 U2623 ( .A1(G79), .A2(n3570), .ZN(n3587) );
  NAND2_X1 U2624 ( .A1(G23), .A2(G2358), .ZN(n3586) );
  NAND3_X1 U2625 ( .A1(n3588), .A2(n3589), .A3(n3590), .ZN(G702) );
  NOR3_X1 U2626 ( .A1(n3591), .A2(n3592), .A3(n3593), .ZN(n3590) );
  NOR2_X1 U2627 ( .A1(G873), .A2(n3594), .ZN(n3593) );
  NOR2_X1 U2628 ( .A1(G834), .A2(n3595), .ZN(n3592) );
  AND2_X1 U2629 ( .A1(n3596), .A2(G149), .ZN(n3591) );
  NAND2_X1 U2630 ( .A1(G146), .A2(n3597), .ZN(n3589) );
  NAND2_X1 U2631 ( .A1(KEYINPUT118), .A2(G137), .ZN(n3588) );
  NAND4_X1 U2632 ( .A1(n3598), .A2(n3599), .A3(n3600), .A4(n3601), .ZN(G699) );
  NAND2_X1 U2633 ( .A1(G155), .A2(n3596), .ZN(n3601) );
  NOR2_X1 U2634 ( .A1(n3602), .A2(n3603), .ZN(n3600) );
  NOR2_X1 U2635 ( .A1(G875), .A2(n3594), .ZN(n3603) );
  NOR2_X1 U2636 ( .A1(G836), .A2(n3595), .ZN(n3602) );
  NAND2_X1 U2637 ( .A1(G152), .A2(n3597), .ZN(n3599) );
  NAND2_X1 U2638 ( .A1(KEYINPUT114), .A2(G137), .ZN(n3598) );
  NAND4_X1 U2639 ( .A1(n3604), .A2(n3605), .A3(n3606), .A4(n3607), .ZN(G696) );
  NAND2_X1 U2640 ( .A1(G188), .A2(n3596), .ZN(n3607) );
  NOR2_X1 U2641 ( .A1(n3608), .A2(n3609), .ZN(n3606) );
  NOR2_X1 U2642 ( .A1(G877), .A2(n3594), .ZN(n3609) );
  NOR2_X1 U2643 ( .A1(G838), .A2(n3595), .ZN(n3608) );
  NAND2_X1 U2644 ( .A1(G158), .A2(n3597), .ZN(n3605) );
  NAND2_X1 U2645 ( .A1(KEYINPUT106), .A2(G137), .ZN(n3604) );
  NAND4_X1 U2646 ( .A1(n3610), .A2(n3611), .A3(n3612), .A4(n3613), .ZN(G693) );
  NAND2_X1 U2647 ( .A1(n3614), .A2(n3406), .ZN(n3613) );
  NAND2_X1 U2648 ( .A1(n3615), .A2(n3399), .ZN(n3612) );
  NAND2_X1 U2649 ( .A1(G182), .A2(n3596), .ZN(n3611) );
  NAND2_X1 U2650 ( .A1(G185), .A2(n3597), .ZN(n3610) );
  NAND3_X1 U2651 ( .A1(n3616), .A2(n3617), .A3(G137), .ZN(G690) );
  NAND2_X1 U2652 ( .A1(n3618), .A2(n3619), .ZN(n3617) );
  NAND2_X1 U2653 ( .A1(n3620), .A2(n3621), .ZN(n3618) );
  NAND2_X1 U2654 ( .A1(n3622), .A2(n3623), .ZN(n3621) );
  NAND2_X1 U2655 ( .A1(n3624), .A2(G1691), .ZN(n3620) );
  NAND2_X1 U2656 ( .A1(n3625), .A2(G1694), .ZN(n3616) );
  NAND2_X1 U2657 ( .A1(n3626), .A2(n3627), .ZN(n3625) );
  NAND2_X1 U2658 ( .A1(G1691), .A2(n3628), .ZN(n3627) );
  NAND2_X1 U2659 ( .A1(n3623), .A2(n3629), .ZN(n3626) );
  NAND4_X1 U2660 ( .A1(n3630), .A2(n3631), .A3(n3632), .A4(n3633), .ZN(G688) );
  NAND2_X1 U2661 ( .A1(G191), .A2(n3596), .ZN(n3633) );
  NOR2_X1 U2662 ( .A1(n3634), .A2(n3635), .ZN(n3632) );
  NOR2_X1 U2663 ( .A1(G863), .A2(n3594), .ZN(n3635) );
  NOR2_X1 U2664 ( .A1(G824), .A2(n3595), .ZN(n3634) );
  NAND2_X1 U2665 ( .A1(G161), .A2(n3597), .ZN(n3631) );
  NAND2_X1 U2666 ( .A1(KEYINPUT93), .A2(G137), .ZN(n3630) );
  NAND4_X1 U2667 ( .A1(n3636), .A2(n3637), .A3(n3638), .A4(n3639), .ZN(G685) );
  NAND2_X1 U2668 ( .A1(n3614), .A2(n3443), .ZN(n3639) );
  NAND2_X1 U2669 ( .A1(n3615), .A2(n3398), .ZN(n3638) );
  NAND2_X1 U2670 ( .A1(G194), .A2(n3596), .ZN(n3637) );
  NAND2_X1 U2671 ( .A1(G164), .A2(n3597), .ZN(n3636) );
  NAND4_X1 U2672 ( .A1(n3640), .A2(n3641), .A3(n3642), .A4(n3643), .ZN(G682) );
  NAND2_X1 U2673 ( .A1(n3615), .A2(n3503), .ZN(n3643) );
  NOR2_X1 U2674 ( .A1(n3644), .A2(n3645), .ZN(n3642) );
  NOR2_X1 U2675 ( .A1(G828), .A2(n3595), .ZN(n3645) );
  NOR2_X1 U2676 ( .A1(n3646), .A2(n3647), .ZN(n3644) );
  NOR2_X1 U2677 ( .A1(KEYINPUT100), .A2(KEYINPUT104), .ZN(n3646) );
  NAND2_X1 U2678 ( .A1(G197), .A2(n3596), .ZN(n3641) );
  NAND2_X1 U2679 ( .A1(G167), .A2(n3597), .ZN(n3640) );
  NAND4_X1 U2680 ( .A1(n3648), .A2(n3649), .A3(n3650), .A4(n3651), .ZN(G679) );
  NAND2_X1 U2681 ( .A1(G203), .A2(n3596), .ZN(n3651) );
  NOR2_X1 U2682 ( .A1(n3652), .A2(n3653), .ZN(n3650) );
  NOR2_X1 U2683 ( .A1(G869), .A2(n3594), .ZN(n3653) );
  NOR2_X1 U2684 ( .A1(G830), .A2(n3595), .ZN(n3652) );
  NAND2_X1 U2685 ( .A1(G173), .A2(n3597), .ZN(n3649) );
  NAND2_X1 U2686 ( .A1(KEYINPUT112), .A2(G137), .ZN(n3648) );
  NAND4_X1 U2687 ( .A1(n3654), .A2(n3655), .A3(n3656), .A4(n3657), .ZN(G676) );
  NAND2_X1 U2688 ( .A1(G200), .A2(n3596), .ZN(n3657) );
  NOR2_X1 U2689 ( .A1(n3658), .A2(n3659), .ZN(n3656) );
  NOR2_X1 U2690 ( .A1(G871), .A2(n3594), .ZN(n3659) );
  INV_X1 U2691 ( .A(n3615), .ZN(n3594) );
  NOR3_X1 U2692 ( .A1(n3647), .A2(G1694), .A3(n3623), .ZN(n3615) );
  NOR2_X1 U2693 ( .A1(G832), .A2(n3595), .ZN(n3658) );
  INV_X1 U2694 ( .A(n3614), .ZN(n3595) );
  NOR3_X1 U2695 ( .A1(G1691), .A2(G1694), .A3(n3647), .ZN(n3614) );
  NAND2_X1 U2696 ( .A1(G170), .A2(n3597), .ZN(n3655) );
  INV_X1 U2697 ( .A(G1694), .ZN(n3619) );
  INV_X1 U2698 ( .A(G1691), .ZN(n3623) );
  NAND2_X1 U2699 ( .A1(KEYINPUT122), .A2(G137), .ZN(n3654) );
  NOR2_X1 U2700 ( .A1(n3660), .A2(n3572), .ZN(G673) );
  NOR3_X1 U2701 ( .A1(n3661), .A2(KEYINPUT83), .A3(KEYINPUT82), .ZN(n3660) );
  NAND3_X1 U2702 ( .A1(n3662), .A2(n3663), .A3(n3444), .ZN(n3661) );
  NAND2_X1 U2703 ( .A1(G26), .A2(n3570), .ZN(n3663) );
  NAND2_X1 U2704 ( .A1(G81), .A2(G2358), .ZN(n3662) );
  NAND3_X1 U2705 ( .A1(n3664), .A2(n3665), .A3(n3666), .ZN(G670) );
  NOR3_X1 U2706 ( .A1(n3667), .A2(n3668), .A3(n3669), .ZN(n3666) );
  NOR2_X1 U2707 ( .A1(G834), .A2(n3670), .ZN(n3669) );
  AND3_X1 U2708 ( .A1(n3671), .A2(n3672), .A3(n3673), .ZN(G834) );
  NAND2_X1 U2709 ( .A1(n3674), .A2(n3675), .ZN(n3673) );
  NAND3_X1 U2710 ( .A1(n3676), .A2(n3677), .A3(n3396), .ZN(n3672) );
  NAND2_X1 U2711 ( .A1(G514), .A2(n3678), .ZN(n3677) );
  NAND2_X1 U2712 ( .A1(G3546), .A2(n3679), .ZN(n3676) );
  NAND2_X1 U2713 ( .A1(G130), .A2(n3680), .ZN(n3671) );
  NOR2_X1 U2714 ( .A1(G873), .A2(n3681), .ZN(n3668) );
  INV_X1 U2715 ( .A(n3535), .ZN(G873) );
  NAND3_X1 U2716 ( .A1(n3682), .A2(n3683), .A3(n3684), .ZN(n3535) );
  NAND2_X1 U2717 ( .A1(G128), .A2(n3680), .ZN(n3684) );
  NAND2_X1 U2718 ( .A1(n3685), .A2(n3675), .ZN(n3683) );
  NAND2_X1 U2719 ( .A1(n3686), .A2(n3396), .ZN(n3682) );
  AND2_X1 U2720 ( .A1(G149), .A2(n3687), .ZN(n3667) );
  NAND2_X1 U2721 ( .A1(n3688), .A2(G146), .ZN(n3665) );
  NAND2_X1 U2722 ( .A1(KEYINPUT117), .A2(G137), .ZN(n3664) );
  NAND4_X1 U2723 ( .A1(n3689), .A2(n3690), .A3(n3691), .A4(n3692), .ZN(G667) );
  NAND2_X1 U2724 ( .A1(n3687), .A2(G155), .ZN(n3692) );
  NOR2_X1 U2725 ( .A1(n3693), .A2(n3694), .ZN(n3691) );
  NOR2_X1 U2726 ( .A1(G836), .A2(n3670), .ZN(n3694) );
  INV_X1 U2727 ( .A(n3478), .ZN(G836) );
  NAND3_X1 U2728 ( .A1(n3695), .A2(n3696), .A3(n3697), .ZN(n3478) );
  NAND2_X1 U2729 ( .A1(G119), .A2(n3680), .ZN(n3697) );
  NAND3_X1 U2730 ( .A1(n3698), .A2(n3699), .A3(n3396), .ZN(n3696) );
  NAND2_X1 U2731 ( .A1(n3700), .A2(n3675), .ZN(n3695) );
  NOR2_X1 U2732 ( .A1(G875), .A2(n3681), .ZN(n3693) );
  INV_X1 U2733 ( .A(n3529), .ZN(G875) );
  NAND3_X1 U2734 ( .A1(n3701), .A2(n3702), .A3(n3703), .ZN(n3529) );
  NAND2_X1 U2735 ( .A1(G127), .A2(n3680), .ZN(n3703) );
  NAND2_X1 U2736 ( .A1(n3704), .A2(n3675), .ZN(n3702) );
  NAND2_X1 U2737 ( .A1(n3705), .A2(n3396), .ZN(n3701) );
  NAND2_X1 U2738 ( .A1(n3688), .A2(G152), .ZN(n3690) );
  NAND2_X1 U2739 ( .A1(KEYINPUT113), .A2(G137), .ZN(n3689) );
  NAND4_X1 U2740 ( .A1(n3706), .A2(n3707), .A3(n3708), .A4(n3709), .ZN(G664) );
  NAND2_X1 U2741 ( .A1(n3687), .A2(G188), .ZN(n3709) );
  NOR2_X1 U2742 ( .A1(n3710), .A2(n3711), .ZN(n3708) );
  NOR2_X1 U2743 ( .A1(G838), .A2(n3670), .ZN(n3711) );
  INV_X1 U2744 ( .A(n3471), .ZN(G838) );
  NAND3_X1 U2745 ( .A1(n3712), .A2(n3713), .A3(n3714), .ZN(n3471) );
  NAND2_X1 U2746 ( .A1(G129), .A2(n3680), .ZN(n3714) );
  NAND3_X1 U2747 ( .A1(n3715), .A2(n3716), .A3(n3396), .ZN(n3713) );
  NAND2_X1 U2748 ( .A1(n3717), .A2(n3675), .ZN(n3712) );
  XNOR2_X1 U2749 ( .A(n3718), .B(n3719), .ZN(n3717) );
  NOR2_X1 U2750 ( .A1(G877), .A2(n3681), .ZN(n3710) );
  INV_X1 U2751 ( .A(n3523), .ZN(G877) );
  NAND3_X1 U2752 ( .A1(n3720), .A2(n3721), .A3(n3722), .ZN(n3523) );
  NAND2_X1 U2753 ( .A1(n3675), .A2(n3723), .ZN(n3722) );
  NAND2_X1 U2754 ( .A1(n3724), .A2(n3396), .ZN(n3721) );
  NAND2_X1 U2755 ( .A1(G126), .A2(n3680), .ZN(n3720) );
  NAND2_X1 U2756 ( .A1(n3688), .A2(G158), .ZN(n3707) );
  NAND2_X1 U2757 ( .A1(KEYINPUT105), .A2(G137), .ZN(n3706) );
  NAND4_X1 U2758 ( .A1(n3725), .A2(n3726), .A3(n3727), .A4(n3728), .ZN(G661) );
  NAND2_X1 U2759 ( .A1(n3729), .A2(n3406), .ZN(n3728) );
  NAND3_X1 U2760 ( .A1(n3730), .A2(n3731), .A3(n3732), .ZN(n3406) );
  NAND2_X1 U2761 ( .A1(G131), .A2(n3680), .ZN(n3732) );
  NAND2_X1 U2762 ( .A1(n3675), .A2(n3733), .ZN(n3731) );
  NAND2_X1 U2763 ( .A1(n3396), .A2(n3734), .ZN(n3730) );
  NAND2_X1 U2764 ( .A1(n3735), .A2(n3399), .ZN(n3727) );
  NAND3_X1 U2765 ( .A1(n3736), .A2(n3737), .A3(n3738), .ZN(n3399) );
  NAND2_X1 U2766 ( .A1(G117), .A2(n3680), .ZN(n3738) );
  NAND2_X1 U2767 ( .A1(n3675), .A2(n3739), .ZN(n3737) );
  NAND2_X1 U2768 ( .A1(n3740), .A2(n3396), .ZN(n3736) );
  NAND2_X1 U2769 ( .A1(n3687), .A2(G182), .ZN(n3726) );
  NAND2_X1 U2770 ( .A1(n3688), .A2(G185), .ZN(n3725) );
  NAND3_X1 U2771 ( .A1(n3741), .A2(n3742), .A3(G137), .ZN(G658) );
  NAND2_X1 U2772 ( .A1(n3743), .A2(n3744), .ZN(n3742) );
  NAND2_X1 U2773 ( .A1(n3745), .A2(n3746), .ZN(n3743) );
  NAND2_X1 U2774 ( .A1(n3622), .A2(n3747), .ZN(n3746) );
  INV_X1 U2775 ( .A(n3466), .ZN(n3622) );
  NAND3_X1 U2776 ( .A1(n3748), .A2(n3749), .A3(n3750), .ZN(n3466) );
  NAND2_X1 U2777 ( .A1(G94), .A2(G4092), .ZN(n3750) );
  NAND3_X1 U2778 ( .A1(n3440), .A2(n3441), .A3(n3675), .ZN(n3749) );
  NAND2_X1 U2779 ( .A1(n3751), .A2(n3752), .ZN(n3441) );
  INV_X1 U2780 ( .A(G2174), .ZN(n3752) );
  XOR2_X1 U2781 ( .A(n3753), .B(n3754), .Z(n3751) );
  XNOR2_X1 U2782 ( .A(n3755), .B(n3756), .ZN(n3754) );
  XOR2_X1 U2783 ( .A(n3757), .B(n3758), .Z(n3753) );
  NOR3_X1 U2784 ( .A1(n3759), .A2(KEYINPUT66), .A3(KEYINPUT43), .ZN(n3758) );
  NAND2_X1 U2785 ( .A1(n3760), .A2(G2174), .ZN(n3440) );
  XOR2_X1 U2786 ( .A(n3761), .B(n3762), .Z(n3760) );
  XNOR2_X1 U2787 ( .A(n3424), .B(n3763), .ZN(n3762) );
  NAND2_X1 U2788 ( .A1(n3764), .A2(n3765), .ZN(n3763) );
  NAND3_X1 U2789 ( .A1(n3766), .A2(n3767), .A3(n3768), .ZN(n3765) );
  OR2_X1 U2790 ( .A1(n3766), .A2(n3768), .ZN(n3764) );
  XOR2_X1 U2791 ( .A(n3757), .B(n3769), .Z(n3761) );
  NOR4_X1 U2792 ( .A1(n3770), .A2(KEYINPUT42), .A3(KEYINPUT67), .A4(KEYINPUT65), .ZN(n3769) );
  NAND3_X1 U2793 ( .A1(n3771), .A2(n3772), .A3(n3773), .ZN(n3770) );
  NAND2_X1 U2794 ( .A1(n3774), .A2(n3775), .ZN(n3773) );
  NAND2_X1 U2795 ( .A1(n3776), .A2(n3766), .ZN(n3771) );
  NAND2_X1 U2796 ( .A1(n3777), .A2(n3778), .ZN(n3766) );
  XOR2_X1 U2797 ( .A(n3779), .B(n3780), .Z(n3757) );
  XNOR2_X1 U2798 ( .A(n3781), .B(n3782), .ZN(n3780) );
  INV_X1 U2799 ( .A(n3783), .ZN(n3782) );
  NAND3_X1 U2800 ( .A1(n3784), .A2(n3785), .A3(n3786), .ZN(n3781) );
  NAND2_X1 U2801 ( .A1(n3787), .A2(n3788), .ZN(n3786) );
  XNOR2_X1 U2802 ( .A(n3718), .B(n3789), .ZN(n3787) );
  NAND3_X1 U2803 ( .A1(n3775), .A2(n3767), .A3(n3718), .ZN(n3785) );
  NAND2_X1 U2804 ( .A1(n3776), .A2(n3777), .ZN(n3784) );
  NAND2_X1 U2805 ( .A1(n3790), .A2(n3791), .ZN(n3779) );
  NAND2_X1 U2806 ( .A1(n3792), .A2(n3793), .ZN(n3791) );
  XOR2_X1 U2807 ( .A(n3794), .B(n3427), .Z(n3792) );
  XOR2_X1 U2808 ( .A(n3795), .B(n3796), .Z(n3794) );
  NOR3_X1 U2809 ( .A1(n3797), .A2(n3798), .A3(n3799), .ZN(n3796) );
  NOR2_X1 U2810 ( .A1(KEYINPUT73), .A2(n3800), .ZN(n3799) );
  NAND3_X1 U2811 ( .A1(n3801), .A2(n3802), .A3(n3803), .ZN(n3795) );
  NAND3_X1 U2812 ( .A1(n3804), .A2(n3805), .A3(n3806), .ZN(n3803) );
  NAND2_X1 U2813 ( .A1(n3807), .A2(n3808), .ZN(n3790) );
  INV_X1 U2814 ( .A(n3793), .ZN(n3808) );
  NAND2_X1 U2815 ( .A1(n3809), .A2(n3810), .ZN(n3793) );
  NAND2_X1 U2816 ( .A1(G2174), .A2(n3811), .ZN(n3810) );
  NAND2_X1 U2817 ( .A1(KEYINPUT30), .A2(n3812), .ZN(n3811) );
  XNOR2_X1 U2818 ( .A(n3813), .B(n3427), .ZN(n3807) );
  XOR2_X1 U2819 ( .A(n3458), .B(n3800), .Z(n3427) );
  NAND3_X1 U2820 ( .A1(n3814), .A2(n3815), .A3(n3816), .ZN(n3813) );
  NAND2_X1 U2821 ( .A1(n3817), .A2(n3806), .ZN(n3816) );
  XNOR2_X1 U2822 ( .A(n3818), .B(n3804), .ZN(n3817) );
  OR3_X1 U2823 ( .A1(n3806), .A2(n3819), .A3(n3818), .ZN(n3815) );
  NAND2_X1 U2824 ( .A1(n3798), .A2(n3818), .ZN(n3814) );
  NAND3_X1 U2825 ( .A1(n3820), .A2(n3821), .A3(n3822), .ZN(n3818) );
  NAND2_X1 U2826 ( .A1(n3823), .A2(n3824), .ZN(n3822) );
  INV_X1 U2827 ( .A(KEYINPUT90), .ZN(n3824) );
  NAND2_X1 U2828 ( .A1(n3825), .A2(n3826), .ZN(n3823) );
  NAND2_X1 U2829 ( .A1(n3827), .A2(n3828), .ZN(n3821) );
  NAND2_X1 U2830 ( .A1(n3825), .A2(n3829), .ZN(n3828) );
  NAND2_X1 U2831 ( .A1(KEYINPUT90), .A2(n3826), .ZN(n3829) );
  INV_X1 U2832 ( .A(n3797), .ZN(n3825) );
  OR3_X1 U2833 ( .A1(n3797), .A2(n3826), .A3(n3827), .ZN(n3820) );
  NOR2_X1 U2834 ( .A1(KEYINPUT74), .A2(n3800), .ZN(n3826) );
  NAND2_X1 U2835 ( .A1(n3830), .A2(n3396), .ZN(n3748) );
  INV_X1 U2836 ( .A(n3442), .ZN(n3830) );
  XNOR2_X1 U2837 ( .A(n3831), .B(n3832), .ZN(n3442) );
  XOR2_X1 U2838 ( .A(n3833), .B(n3834), .Z(n3832) );
  XOR2_X1 U2839 ( .A(n3835), .B(n3836), .Z(n3834) );
  NAND2_X1 U2840 ( .A1(n3837), .A2(n3838), .ZN(n3835) );
  NAND2_X1 U2841 ( .A1(n3839), .A2(n3679), .ZN(n3838) );
  XNOR2_X1 U2842 ( .A(G242), .B(n3840), .ZN(n3839) );
  NAND2_X1 U2843 ( .A1(n3841), .A2(G514), .ZN(n3837) );
  XNOR2_X1 U2844 ( .A(n3840), .B(n3842), .ZN(n3841) );
  NAND2_X1 U2845 ( .A1(n3843), .A2(n3844), .ZN(n3840) );
  NAND2_X1 U2846 ( .A1(n3845), .A2(n3846), .ZN(n3844) );
  NAND2_X1 U2847 ( .A1(n3847), .A2(n3848), .ZN(n3845) );
  NAND2_X1 U2848 ( .A1(n3849), .A2(n3850), .ZN(n3848) );
  NAND2_X1 U2849 ( .A1(G351), .A2(n3851), .ZN(n3847) );
  NAND2_X1 U2850 ( .A1(n3852), .A2(G534), .ZN(n3843) );
  NAND2_X1 U2851 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  NAND2_X1 U2852 ( .A1(G251), .A2(n3850), .ZN(n3854) );
  NAND2_X1 U2853 ( .A1(G351), .A2(G248), .ZN(n3853) );
  XOR2_X1 U2854 ( .A(n3855), .B(n3856), .Z(n3833) );
  XOR2_X1 U2855 ( .A(n3857), .B(n3858), .Z(n3831) );
  XOR2_X1 U2856 ( .A(n3859), .B(n3453), .Z(n3858) );
  NAND2_X1 U2857 ( .A1(n3860), .A2(n3861), .ZN(n3859) );
  NAND2_X1 U2858 ( .A1(n3862), .A2(n3863), .ZN(n3861) );
  NAND2_X1 U2859 ( .A1(n3864), .A2(n3865), .ZN(n3862) );
  NAND2_X1 U2860 ( .A1(n3849), .A2(n3866), .ZN(n3865) );
  NAND2_X1 U2861 ( .A1(G324), .A2(n3851), .ZN(n3864) );
  NAND2_X1 U2862 ( .A1(n3867), .A2(G503), .ZN(n3860) );
  NAND2_X1 U2863 ( .A1(n3868), .A2(n3869), .ZN(n3867) );
  NAND2_X1 U2864 ( .A1(G251), .A2(n3866), .ZN(n3869) );
  NAND2_X1 U2865 ( .A1(G324), .A2(G248), .ZN(n3868) );
  XNOR2_X1 U2866 ( .A(n3870), .B(n3734), .ZN(n3857) );
  NAND2_X1 U2867 ( .A1(n3871), .A2(n3872), .ZN(n3870) );
  NAND2_X1 U2868 ( .A1(n3873), .A2(n3874), .ZN(n3872) );
  NAND2_X1 U2869 ( .A1(n3875), .A2(n3876), .ZN(n3873) );
  NAND2_X1 U2870 ( .A1(n3849), .A2(n3877), .ZN(n3876) );
  NAND2_X1 U2871 ( .A1(G341), .A2(n3851), .ZN(n3875) );
  NAND2_X1 U2872 ( .A1(n3878), .A2(G523), .ZN(n3871) );
  NAND2_X1 U2873 ( .A1(n3879), .A2(n3880), .ZN(n3878) );
  NAND2_X1 U2874 ( .A1(G251), .A2(n3877), .ZN(n3880) );
  NAND2_X1 U2875 ( .A1(G341), .A2(G248), .ZN(n3879) );
  NAND2_X1 U2876 ( .A1(n3624), .A2(G1689), .ZN(n3745) );
  INV_X1 U2877 ( .A(n3465), .ZN(n3624) );
  NAND3_X1 U2878 ( .A1(n3881), .A2(n3882), .A3(n3883), .ZN(n3465) );
  NAND2_X1 U2879 ( .A1(G97), .A2(G4092), .ZN(n3883) );
  NAND3_X1 U2880 ( .A1(n3393), .A2(n3394), .A3(n3675), .ZN(n3882) );
  NAND2_X1 U2881 ( .A1(n3884), .A2(n3885), .ZN(n3394) );
  INV_X1 U2882 ( .A(G1497), .ZN(n3885) );
  XNOR2_X1 U2883 ( .A(n3886), .B(n3887), .ZN(n3884) );
  XOR2_X1 U2884 ( .A(n3888), .B(n3889), .Z(n3887) );
  NOR4_X1 U2885 ( .A1(KEYINPUT60), .A2(n3890), .A3(n3891), .A4(n3892), .ZN(n3888) );
  XNOR2_X1 U2886 ( .A(n3893), .B(n3894), .ZN(n3886) );
  XNOR2_X1 U2887 ( .A(n3895), .B(n3896), .ZN(n3894) );
  NOR4_X1 U2888 ( .A1(KEYINPUT58), .A2(KEYINPUT27), .A3(n3897), .A4(n3898),  .ZN(n3896) );
  NOR2_X1 U2889 ( .A1(n3899), .A2(n3900), .ZN(n3897) );
  NOR2_X1 U2890 ( .A1(n3891), .A2(n3892), .ZN(n3899) );
  NOR3_X1 U2891 ( .A1(n3895), .A2(n3901), .A3(n3902), .ZN(n3892) );
  NOR2_X1 U2892 ( .A1(n3903), .A2(n3902), .ZN(n3891) );
  NAND2_X1 U2893 ( .A1(n3904), .A2(G1497), .ZN(n3393) );
  XOR2_X1 U2894 ( .A(n3905), .B(n3906), .Z(n3904) );
  XNOR2_X1 U2895 ( .A(n3907), .B(n3889), .ZN(n3906) );
  XNOR2_X1 U2896 ( .A(n3908), .B(n3909), .ZN(n3889) );
  XOR2_X1 U2897 ( .A(n3910), .B(n3911), .Z(n3909) );
  XNOR2_X1 U2898 ( .A(n3902), .B(n3912), .ZN(n3911) );
  NOR4_X1 U2899 ( .A1(n3913), .A2(n3914), .A3(KEYINPUT95), .A4(KEYINPUT88),  .ZN(n3912) );
  NOR2_X1 U2900 ( .A1(n3915), .A2(n3916), .ZN(n3914) );
  XOR2_X1 U2901 ( .A(n3917), .B(n3918), .Z(n3915) );
  XNOR2_X1 U2902 ( .A(n3919), .B(n3920), .ZN(n3918) );
  NAND2_X1 U2903 ( .A1(n3921), .A2(n3922), .ZN(n3917) );
  NAND2_X1 U2904 ( .A1(n3923), .A2(n3924), .ZN(n3922) );
  NAND2_X1 U2905 ( .A1(n3925), .A2(n3926), .ZN(n3923) );
  NAND4_X1 U2906 ( .A1(n3927), .A2(n3926), .A3(n3928), .A4(n3929), .ZN(n3921) );
  INV_X1 U2907 ( .A(n3924), .ZN(n3929) );
  NAND2_X1 U2908 ( .A1(n3930), .A2(KEYINPUT89), .ZN(n3924) );
  XOR2_X1 U2909 ( .A(n3931), .B(n3932), .Z(n3930) );
  NAND2_X1 U2910 ( .A1(n3933), .A2(n3934), .ZN(n3928) );
  INV_X1 U2911 ( .A(KEYINPUT55), .ZN(n3926) );
  NOR2_X1 U2912 ( .A1(n3935), .A2(n3936), .ZN(n3913) );
  XOR2_X1 U2913 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR2_X1 U2914 ( .A(n3939), .B(n3940), .Z(n3938) );
  NOR2_X1 U2915 ( .A1(KEYINPUT54), .A2(n3941), .ZN(n3940) );
  NAND2_X1 U2916 ( .A1(n3942), .A2(n3943), .ZN(n3939) );
  NAND2_X1 U2917 ( .A1(n3932), .A2(n3944), .ZN(n3943) );
  OR3_X1 U2918 ( .A1(n3932), .A2(n3945), .A3(n3944), .ZN(n3942) );
  XOR2_X1 U2919 ( .A(n3920), .B(n3946), .Z(n3937) );
  NAND3_X1 U2920 ( .A1(n3947), .A2(n3948), .A3(n3949), .ZN(n3920) );
  NAND2_X1 U2921 ( .A1(n3950), .A2(n3951), .ZN(n3948) );
  INV_X1 U2922 ( .A(n3952), .ZN(n3951) );
  XNOR2_X1 U2923 ( .A(n3934), .B(n3953), .ZN(n3950) );
  NAND3_X1 U2924 ( .A1(n3953), .A2(n3954), .A3(n3952), .ZN(n3947) );
  INV_X1 U2925 ( .A(n3916), .ZN(n3935) );
  NAND2_X1 U2926 ( .A1(n3955), .A2(n3956), .ZN(n3916) );
  NAND2_X1 U2927 ( .A1(G1497), .A2(n3957), .ZN(n3956) );
  NAND2_X1 U2928 ( .A1(KEYINPUT15), .A2(n3958), .ZN(n3957) );
  NOR2_X1 U2929 ( .A1(n3959), .A2(n3960), .ZN(n3910) );
  AND2_X1 U2930 ( .A1(n3961), .A2(n3901), .ZN(n3959) );
  XNOR2_X1 U2931 ( .A(n3962), .B(n3963), .ZN(n3908) );
  NAND3_X1 U2932 ( .A1(n3964), .A2(n3965), .A3(n3966), .ZN(n3907) );
  NOR3_X1 U2933 ( .A1(KEYINPUT26), .A2(KEYINPUT57), .A3(KEYINPUT40), .ZN(n3966) );
  NAND2_X1 U2934 ( .A1(n3960), .A2(n3967), .ZN(n3965) );
  INV_X1 U2935 ( .A(n3968), .ZN(n3964) );
  NAND2_X1 U2936 ( .A1(n3969), .A2(n3970), .ZN(n3905) );
  NAND2_X1 U2937 ( .A1(n3971), .A2(n3972), .ZN(n3970) );
  NAND2_X1 U2938 ( .A1(n3973), .A2(n3903), .ZN(n3972) );
  NAND2_X1 U2939 ( .A1(n3974), .A2(n3975), .ZN(n3973) );
  NAND2_X1 U2940 ( .A1(n3961), .A2(n3895), .ZN(n3975) );
  OR3_X1 U2941 ( .A1(n3976), .A2(n3960), .A3(n3971), .ZN(n3969) );
  XNOR2_X1 U2942 ( .A(n3977), .B(n3978), .ZN(n3971) );
  NOR3_X1 U2943 ( .A1(n3979), .A2(KEYINPUT59), .A3(n3890), .ZN(n3978) );
  NOR2_X1 U2944 ( .A1(n3980), .A2(n3902), .ZN(n3979) );
  NOR2_X1 U2945 ( .A1(n3960), .A2(n3976), .ZN(n3980) );
  NAND2_X1 U2946 ( .A1(n3396), .A2(n3981), .ZN(n3881) );
  INV_X1 U2947 ( .A(n3397), .ZN(n3981) );
  XOR2_X1 U2948 ( .A(n3982), .B(n3983), .Z(n3397) );
  XOR2_X1 U2949 ( .A(n3984), .B(n3985), .Z(n3983) );
  XOR2_X1 U2950 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR2_X1 U2951 ( .A(n3988), .B(n3989), .Z(n3987) );
  NAND2_X1 U2952 ( .A1(n3990), .A2(n3991), .ZN(n3989) );
  NAND2_X1 U2953 ( .A1(n3992), .A2(n3993), .ZN(n3991) );
  NAND2_X1 U2954 ( .A1(n3994), .A2(n3995), .ZN(n3992) );
  NAND2_X1 U2955 ( .A1(G234), .A2(n3851), .ZN(n3995) );
  NAND2_X1 U2956 ( .A1(n3996), .A2(n3849), .ZN(n3994) );
  NAND2_X1 U2957 ( .A1(n3997), .A2(G435), .ZN(n3990) );
  NAND2_X1 U2958 ( .A1(n3998), .A2(n3999), .ZN(n3997) );
  NAND2_X1 U2959 ( .A1(G251), .A2(n3996), .ZN(n3999) );
  NAND2_X1 U2960 ( .A1(G234), .A2(G248), .ZN(n3998) );
  NAND2_X1 U2961 ( .A1(n4000), .A2(n4001), .ZN(n3988) );
  NAND2_X1 U2962 ( .A1(n4002), .A2(n4003), .ZN(n4001) );
  NAND2_X1 U2963 ( .A1(n4004), .A2(n4005), .ZN(n4002) );
  NAND2_X1 U2964 ( .A1(n3849), .A2(n4006), .ZN(n4005) );
  NAND2_X1 U2965 ( .A1(G273), .A2(n3851), .ZN(n4004) );
  NAND2_X1 U2966 ( .A1(n4007), .A2(G411), .ZN(n4000) );
  NAND2_X1 U2967 ( .A1(n4008), .A2(n4009), .ZN(n4007) );
  NAND2_X1 U2968 ( .A1(G251), .A2(n4006), .ZN(n4009) );
  NAND2_X1 U2969 ( .A1(G273), .A2(G248), .ZN(n4008) );
  XOR2_X1 U2970 ( .A(n4010), .B(n4011), .Z(n3986) );
  NAND2_X1 U2971 ( .A1(n4012), .A2(n4013), .ZN(n4011) );
  NAND2_X1 U2972 ( .A1(n4014), .A2(n4015), .ZN(n4013) );
  NAND2_X1 U2973 ( .A1(n4016), .A2(n4017), .ZN(n4014) );
  NAND2_X1 U2974 ( .A1(G226), .A2(n3851), .ZN(n4017) );
  NAND2_X1 U2975 ( .A1(n4018), .A2(n3849), .ZN(n4016) );
  NAND2_X1 U2976 ( .A1(n4019), .A2(G422), .ZN(n4012) );
  NAND2_X1 U2977 ( .A1(n4020), .A2(n4021), .ZN(n4019) );
  NAND2_X1 U2978 ( .A1(G251), .A2(n4018), .ZN(n4021) );
  NAND2_X1 U2979 ( .A1(G226), .A2(G248), .ZN(n4020) );
  NAND2_X1 U2980 ( .A1(n4022), .A2(n4023), .ZN(n4010) );
  NAND2_X1 U2981 ( .A1(n4024), .A2(n4025), .ZN(n4023) );
  NAND2_X1 U2982 ( .A1(n4026), .A2(n4027), .ZN(n4024) );
  NAND2_X1 U2983 ( .A1(n3849), .A2(n4028), .ZN(n4027) );
  NAND2_X1 U2984 ( .A1(G265), .A2(n3851), .ZN(n4026) );
  NAND2_X1 U2985 ( .A1(n4029), .A2(G400), .ZN(n4022) );
  NAND2_X1 U2986 ( .A1(n4030), .A2(n4031), .ZN(n4029) );
  NAND2_X1 U2987 ( .A1(G251), .A2(n4028), .ZN(n4031) );
  NAND2_X1 U2988 ( .A1(G265), .A2(G248), .ZN(n4030) );
  XOR2_X1 U2989 ( .A(n4032), .B(n4033), .Z(n3984) );
  XOR2_X1 U2990 ( .A(n4034), .B(n4035), .Z(n4033) );
  NAND2_X1 U2991 ( .A1(n4036), .A2(n4037), .ZN(n4035) );
  NAND2_X1 U2992 ( .A1(n4038), .A2(n4039), .ZN(n4037) );
  NAND2_X1 U2993 ( .A1(n4040), .A2(n4041), .ZN(n4038) );
  NAND2_X1 U2994 ( .A1(n3849), .A2(n4042), .ZN(n4041) );
  NAND2_X1 U2995 ( .A1(G281), .A2(n3851), .ZN(n4040) );
  NAND2_X1 U2996 ( .A1(n4043), .A2(G374), .ZN(n4036) );
  NAND2_X1 U2997 ( .A1(n4044), .A2(n4045), .ZN(n4043) );
  NAND2_X1 U2998 ( .A1(G251), .A2(n4042), .ZN(n4045) );
  NAND2_X1 U2999 ( .A1(G281), .A2(G248), .ZN(n4044) );
  NAND2_X1 U3000 ( .A1(n4046), .A2(n4047), .ZN(n4034) );
  NAND2_X1 U3001 ( .A1(n4048), .A2(n4049), .ZN(n4047) );
  NAND2_X1 U3002 ( .A1(n4050), .A2(n4051), .ZN(n4048) );
  NAND2_X1 U3003 ( .A1(n3849), .A2(n4052), .ZN(n4051) );
  NAND2_X1 U3004 ( .A1(G257), .A2(n3851), .ZN(n4050) );
  NAND2_X1 U3005 ( .A1(n4053), .A2(G389), .ZN(n4046) );
  NAND2_X1 U3006 ( .A1(n4054), .A2(n4055), .ZN(n4053) );
  NAND2_X1 U3007 ( .A1(G251), .A2(n4052), .ZN(n4055) );
  NAND2_X1 U3008 ( .A1(G257), .A2(G248), .ZN(n4054) );
  XOR2_X1 U3009 ( .A(n4056), .B(n4057), .Z(n4032) );
  NAND2_X1 U3010 ( .A1(n4058), .A2(n4059), .ZN(n4057) );
  NAND2_X1 U3011 ( .A1(n4060), .A2(n4061), .ZN(n4059) );
  NAND2_X1 U3012 ( .A1(n4062), .A2(n4063), .ZN(n4060) );
  NAND2_X1 U3013 ( .A1(G218), .A2(n3851), .ZN(n4063) );
  NAND2_X1 U3014 ( .A1(n4064), .A2(n3849), .ZN(n4062) );
  NAND2_X1 U3015 ( .A1(n4065), .A2(G468), .ZN(n4058) );
  NAND2_X1 U3016 ( .A1(n4066), .A2(n4067), .ZN(n4065) );
  NAND2_X1 U3017 ( .A1(G251), .A2(n4064), .ZN(n4067) );
  NAND2_X1 U3018 ( .A1(G218), .A2(G248), .ZN(n4066) );
  NAND2_X1 U3019 ( .A1(n4068), .A2(n4069), .ZN(n4056) );
  NAND2_X1 U3020 ( .A1(n4070), .A2(n4071), .ZN(n4069) );
  NAND2_X1 U3021 ( .A1(n4072), .A2(n4073), .ZN(n4070) );
  NAND2_X1 U3022 ( .A1(G210), .A2(n3851), .ZN(n4073) );
  NAND2_X1 U3023 ( .A1(n4074), .A2(n3849), .ZN(n4072) );
  NAND2_X1 U3024 ( .A1(n4075), .A2(G457), .ZN(n4068) );
  NAND2_X1 U3025 ( .A1(n4076), .A2(n4077), .ZN(n4075) );
  NAND2_X1 U3026 ( .A1(G251), .A2(n4074), .ZN(n4077) );
  NAND2_X1 U3027 ( .A1(G210), .A2(G248), .ZN(n4076) );
  NAND2_X1 U3028 ( .A1(n4078), .A2(G1690), .ZN(n3741) );
  NAND2_X1 U3029 ( .A1(n4079), .A2(n4080), .ZN(n4078) );
  NAND2_X1 U3030 ( .A1(G1689), .A2(n3628), .ZN(n4080) );
  INV_X1 U3031 ( .A(G179), .ZN(n3628) );
  NAND2_X1 U3032 ( .A1(n3747), .A2(n3629), .ZN(n4079) );
  INV_X1 U3033 ( .A(G176), .ZN(n3629) );
  NAND2_X1 U3034 ( .A1(G140), .A2(n3444), .ZN(G656) );
  NAND4_X1 U3035 ( .A1(n4081), .A2(n4082), .A3(n4083), .A4(n4084), .ZN(G654) );
  NAND2_X1 U3036 ( .A1(n3687), .A2(G191), .ZN(n4084) );
  NOR2_X1 U3037 ( .A1(n4085), .A2(n4086), .ZN(n4083) );
  NOR2_X1 U3038 ( .A1(G824), .A2(n3670), .ZN(n4086) );
  INV_X1 U3039 ( .A(n3580), .ZN(G824) );
  NAND3_X1 U3040 ( .A1(n4087), .A2(n4088), .A3(n4089), .ZN(n3580) );
  NAND2_X1 U3041 ( .A1(n3675), .A2(n4090), .ZN(n4089) );
  NAND2_X1 U3042 ( .A1(n3396), .A2(n3453), .ZN(n4088) );
  NAND2_X1 U3043 ( .A1(G123), .A2(n3680), .ZN(n4087) );
  NOR2_X1 U3044 ( .A1(G863), .A2(n3681), .ZN(n4085) );
  INV_X1 U3045 ( .A(n3561), .ZN(G863) );
  NAND3_X1 U3046 ( .A1(n4091), .A2(n4092), .A3(n4093), .ZN(n3561) );
  NAND2_X1 U3047 ( .A1(n4094), .A2(n3675), .ZN(n4093) );
  NAND2_X1 U3048 ( .A1(n3396), .A2(n3982), .ZN(n4092) );
  NAND2_X1 U3049 ( .A1(G115), .A2(n3680), .ZN(n4091) );
  NAND2_X1 U3050 ( .A1(n3688), .A2(G161), .ZN(n4082) );
  NAND2_X1 U3051 ( .A1(KEYINPUT92), .A2(G137), .ZN(n4081) );
  NAND4_X1 U3052 ( .A1(n4095), .A2(n4096), .A3(n4097), .A4(n4098), .ZN(G651) );
  NAND2_X1 U3053 ( .A1(n3729), .A2(n3443), .ZN(n4098) );
  NAND3_X1 U3054 ( .A1(n4099), .A2(n4100), .A3(n4101), .ZN(n3443) );
  NAND2_X1 U3055 ( .A1(n3675), .A2(n4102), .ZN(n4101) );
  NAND2_X1 U3056 ( .A1(n3396), .A2(n3856), .ZN(n4100) );
  NAND2_X1 U3057 ( .A1(G121), .A2(n3680), .ZN(n4099) );
  NAND2_X1 U3058 ( .A1(n3735), .A2(n3398), .ZN(n4097) );
  NAND3_X1 U3059 ( .A1(n4103), .A2(n4104), .A3(n4105), .ZN(n3398) );
  NAND2_X1 U3060 ( .A1(n4106), .A2(n3675), .ZN(n4105) );
  NAND2_X1 U3061 ( .A1(n4107), .A2(n3396), .ZN(n4104) );
  NAND2_X1 U3062 ( .A1(G114), .A2(n3680), .ZN(n4103) );
  NAND2_X1 U3063 ( .A1(n3687), .A2(G194), .ZN(n4096) );
  NAND2_X1 U3064 ( .A1(n3688), .A2(G164), .ZN(n4095) );
  NAND4_X1 U3065 ( .A1(n4108), .A2(n4109), .A3(n4110), .A4(n4111), .ZN(G648) );
  NAND2_X1 U3066 ( .A1(n3735), .A2(n3503), .ZN(n4111) );
  NAND3_X1 U3067 ( .A1(n4112), .A2(n4113), .A3(n4114), .ZN(n3503) );
  NAND2_X1 U3068 ( .A1(n4115), .A2(n3675), .ZN(n4114) );
  NAND2_X1 U3069 ( .A1(n4116), .A2(n3396), .ZN(n4113) );
  NAND2_X1 U3070 ( .A1(G53), .A2(n3680), .ZN(n4112) );
  NOR2_X1 U3071 ( .A1(n4117), .A2(n4118), .ZN(n4110) );
  NOR2_X1 U3072 ( .A1(G828), .A2(n3670), .ZN(n4118) );
  INV_X1 U3073 ( .A(n3504), .ZN(G828) );
  NAND3_X1 U3074 ( .A1(n4119), .A2(n4120), .A3(n4121), .ZN(n3504) );
  NAND2_X1 U3075 ( .A1(n3675), .A2(n4122), .ZN(n4121) );
  NAND2_X1 U3076 ( .A1(n3836), .A2(n3396), .ZN(n4120) );
  NAND2_X1 U3077 ( .A1(G116), .A2(n3680), .ZN(n4119) );
  NOR2_X1 U3078 ( .A1(n4123), .A2(n3647), .ZN(n4117) );
  NOR2_X1 U3079 ( .A1(KEYINPUT103), .A2(KEYINPUT99), .ZN(n4123) );
  NAND2_X1 U3080 ( .A1(n3687), .A2(G197), .ZN(n4109) );
  NAND2_X1 U3081 ( .A1(n3688), .A2(G167), .ZN(n4108) );
  NAND4_X1 U3082 ( .A1(n4124), .A2(n4125), .A3(n4126), .A4(n4127), .ZN(G645) );
  NAND2_X1 U3083 ( .A1(n3687), .A2(G203), .ZN(n4127) );
  NOR2_X1 U3084 ( .A1(n4128), .A2(n4129), .ZN(n4126) );
  NOR2_X1 U3085 ( .A1(G869), .A2(n3681), .ZN(n4129) );
  INV_X1 U3086 ( .A(n3546), .ZN(G869) );
  NAND3_X1 U3087 ( .A1(n4130), .A2(n4131), .A3(n4132), .ZN(n3546) );
  NAND2_X1 U3088 ( .A1(G113), .A2(n3680), .ZN(n4132) );
  NAND2_X1 U3089 ( .A1(n4133), .A2(n3675), .ZN(n4131) );
  NAND2_X1 U3090 ( .A1(n4134), .A2(n3396), .ZN(n4130) );
  NOR2_X1 U3091 ( .A1(G830), .A2(n3670), .ZN(n4128) );
  INV_X1 U3092 ( .A(n3496), .ZN(G830) );
  NAND3_X1 U3093 ( .A1(n4135), .A2(n4136), .A3(n4137), .ZN(n3496) );
  NAND2_X1 U3094 ( .A1(G112), .A2(n3680), .ZN(n4137) );
  NAND2_X1 U3095 ( .A1(n4138), .A2(n3675), .ZN(n4136) );
  XNOR2_X1 U3096 ( .A(n3819), .B(n4139), .ZN(n4138) );
  INV_X1 U3097 ( .A(n3804), .ZN(n3819) );
  NAND2_X1 U3098 ( .A1(n3855), .A2(n3396), .ZN(n4135) );
  NAND2_X1 U3099 ( .A1(n3688), .A2(G173), .ZN(n4125) );
  NAND2_X1 U3100 ( .A1(KEYINPUT111), .A2(G137), .ZN(n4124) );
  NAND4_X1 U3101 ( .A1(n4140), .A2(n4141), .A3(n4142), .A4(n4143), .ZN(G642) );
  NAND2_X1 U3102 ( .A1(n3687), .A2(G200), .ZN(n4143) );
  NOR2_X1 U3103 ( .A1(n4144), .A2(n4145), .ZN(n4142) );
  NOR2_X1 U3104 ( .A1(G871), .A2(n3681), .ZN(n4145) );
  INV_X1 U3105 ( .A(n3735), .ZN(n3681) );
  NOR3_X1 U3106 ( .A1(n3647), .A2(G1690), .A3(n3747), .ZN(n3735) );
  INV_X1 U3107 ( .A(n3490), .ZN(G871) );
  NAND3_X1 U3108 ( .A1(n4146), .A2(n4147), .A3(n4148), .ZN(n3490) );
  NAND2_X1 U3109 ( .A1(G122), .A2(n3680), .ZN(n4148) );
  NAND2_X1 U3110 ( .A1(n4149), .A2(n3675), .ZN(n4147) );
  NAND2_X1 U3111 ( .A1(n4150), .A2(n3396), .ZN(n4146) );
  NOR2_X1 U3112 ( .A1(G832), .A2(n3670), .ZN(n4144) );
  INV_X1 U3113 ( .A(n3729), .ZN(n3670) );
  NOR3_X1 U3114 ( .A1(G1689), .A2(G1690), .A3(n3647), .ZN(n3729) );
  INV_X1 U3115 ( .A(n3491), .ZN(G832) );
  NAND3_X1 U3116 ( .A1(n4151), .A2(n4152), .A3(n4153), .ZN(n3491) );
  NAND2_X1 U3117 ( .A1(G52), .A2(n3680), .ZN(n4153) );
  NAND2_X1 U3118 ( .A1(n4154), .A2(n3675), .ZN(n4152) );
  AND2_X1 U3119 ( .A1(G4091), .A2(n3395), .ZN(n3675) );
  INV_X1 U3120 ( .A(G4092), .ZN(n3395) );
  NAND2_X1 U3121 ( .A1(n4155), .A2(n3396), .ZN(n4151) );
  NAND2_X1 U3122 ( .A1(n3688), .A2(G170), .ZN(n4141) );
  INV_X1 U3123 ( .A(G1690), .ZN(n3744) );
  INV_X1 U3124 ( .A(G137), .ZN(n3647) );
  INV_X1 U3125 ( .A(G1689), .ZN(n3747) );
  NAND2_X1 U3126 ( .A1(KEYINPUT121), .A2(G137), .ZN(n4140) );
  NOR2_X1 U3127 ( .A1(n4156), .A2(n3572), .ZN(G639) );
  INV_X1 U3128 ( .A(G141), .ZN(n3572) );
  NOR3_X1 U3129 ( .A1(n4157), .A2(KEYINPUT81), .A3(KEYINPUT80), .ZN(n4156) );
  NAND3_X1 U3130 ( .A1(n4158), .A2(n4159), .A3(n3444), .ZN(n4157) );
  INV_X1 U3131 ( .A(G809), .ZN(n3444) );
  NAND2_X1 U3132 ( .A1(G24), .A2(n3570), .ZN(n4159) );
  NAND2_X1 U3133 ( .A1(G25), .A2(G2358), .ZN(n4158) );
  OR3_X1 U3134 ( .A1(n4160), .A2(n4161), .A3(G809), .ZN(G636) );
  NAND2_X1 U3135 ( .A1(G31), .A2(G27), .ZN(G809) );
  NOR2_X1 U3136 ( .A1(G86), .A2(G2358), .ZN(n4161) );
  NOR2_X1 U3137 ( .A1(G87), .A2(n3570), .ZN(n4160) );
  INV_X1 U3138 ( .A(G2358), .ZN(n3570) );
  AND2_X1 U3139 ( .A1(G1), .A2(G373), .ZN(G634) );
  OR2_X1 U3140 ( .A1(n4162), .A2(KEYINPUT1), .ZN(G632_enc) );
  NOR2_X1 U3141 ( .A1(n4163), .A2(n4164), .ZN(n4162) );
  NAND3_X1 U3142 ( .A1(n4165), .A2(n4166), .A3(n4167), .ZN(G629) );
  NOR3_X1 U3143 ( .A1(KEYINPUT34), .A2(KEYINPUT79), .A3(KEYINPUT37), .ZN(n4167) );
  NAND2_X1 U3144 ( .A1(n4168), .A2(n4169), .ZN(n4166) );
  INV_X1 U3145 ( .A(n3809), .ZN(n4169) );
  NOR4_X1 U3146 ( .A1(KEYINPUT19), .A2(n4170), .A3(KEYINPUT64), .A4(KEYINPUT29), .ZN(n3809) );
  OR2_X1 U3147 ( .A1(n4171), .A2(KEYINPUT76), .ZN(n4168) );
  OR2_X1 U3148 ( .A1(n4172), .A2(KEYINPUT5), .ZN(G626_enc) );
  NOR2_X1 U3149 ( .A1(n3812), .A2(n4173), .ZN(n4172) );
  NOR2_X1 U3150 ( .A1(n4171), .A2(KEYINPUT76), .ZN(n4173) );
  NOR2_X1 U3151 ( .A1(n4174), .A2(KEYINPUT32), .ZN(n3812) );
  NAND3_X1 U3152 ( .A1(n4175), .A2(n4176), .A3(n4177), .ZN(G621) );
  NOR3_X1 U3153 ( .A1(KEYINPUT14), .A2(KEYINPUT48), .A3(KEYINPUT22), .ZN(n4177) );
  NAND2_X1 U3154 ( .A1(n4178), .A2(n4179), .ZN(n4176) );
  INV_X1 U3155 ( .A(n4163), .ZN(n4178) );
  NOR2_X1 U3156 ( .A1(n4180), .A2(KEYINPUT38), .ZN(n4163) );
  NAND3_X1 U3157 ( .A1(n4165), .A2(n4181), .A3(n4182), .ZN(G618) );
  NOR3_X1 U3158 ( .A1(KEYINPUT33), .A2(KEYINPUT78), .A3(KEYINPUT36), .ZN(n4182) );
  NAND2_X1 U3159 ( .A1(n4183), .A2(n4184), .ZN(n4181) );
  INV_X1 U3160 ( .A(n4185), .ZN(n4183) );
  NOR3_X1 U3161 ( .A1(n3458), .A2(n3800), .A3(n3797), .ZN(n4165) );
  OR2_X1 U3162 ( .A1(n4186), .A2(KEYINPUT4), .ZN(G615_enc) );
  NOR2_X1 U3163 ( .A1(n4185), .A2(n4187), .ZN(n4186) );
  NOR2_X1 U3164 ( .A1(n4171), .A2(KEYINPUT75), .ZN(n4185) );
  NOR3_X1 U3165 ( .A1(n3458), .A2(n3800), .A3(n3802), .ZN(n4171) );
  INV_X1 U3166 ( .A(G358), .ZN(G612) );
  INV_X1 U3167 ( .A(G338), .ZN(G611) );
  OR2_X1 U3168 ( .A1(n4188), .A2(KEYINPUT3), .ZN(G610_enc) );
  NOR3_X1 U3169 ( .A1(n3982), .A2(n4189), .A3(n4190), .ZN(n4188) );
  NOR2_X1 U3170 ( .A1(n4191), .A2(KEYINPUT45), .ZN(n4190) );
  NOR4_X1 U3171 ( .A1(n3724), .A2(n3705), .A3(n3686), .A4(n3740), .ZN(n4191) );
  AND2_X1 U3172 ( .A1(n4192), .A2(n4193), .ZN(n3740) );
  NAND2_X1 U3173 ( .A1(n4194), .A2(n4039), .ZN(n4193) );
  NAND2_X1 U3174 ( .A1(n4195), .A2(n4196), .ZN(n4194) );
  NAND2_X1 U3175 ( .A1(G3548), .A2(n4042), .ZN(n4196) );
  NAND2_X1 U3176 ( .A1(G281), .A2(G3546), .ZN(n4195) );
  NAND2_X1 U3177 ( .A1(n4197), .A2(G374), .ZN(n4192) );
  NAND2_X1 U3178 ( .A1(n4198), .A2(n4199), .ZN(n4197) );
  NAND2_X1 U3179 ( .A1(G281), .A2(n3678), .ZN(n4199) );
  NAND2_X1 U3180 ( .A1(n4042), .A2(n4200), .ZN(n4198) );
  INV_X1 U3181 ( .A(G281), .ZN(n4042) );
  AND2_X1 U3182 ( .A1(n4201), .A2(n4202), .ZN(n3686) );
  NAND2_X1 U3183 ( .A1(n4203), .A2(n4049), .ZN(n4202) );
  INV_X1 U3184 ( .A(G389), .ZN(n4049) );
  NAND2_X1 U3185 ( .A1(n4204), .A2(n4205), .ZN(n4203) );
  NAND2_X1 U3186 ( .A1(G3548), .A2(n4052), .ZN(n4205) );
  NAND2_X1 U3187 ( .A1(G257), .A2(G3546), .ZN(n4204) );
  NAND2_X1 U3188 ( .A1(n4206), .A2(G389), .ZN(n4201) );
  NAND2_X1 U3189 ( .A1(n4207), .A2(n4208), .ZN(n4206) );
  NAND2_X1 U3190 ( .A1(G257), .A2(n3678), .ZN(n4208) );
  NAND2_X1 U3191 ( .A1(n4052), .A2(n4200), .ZN(n4207) );
  AND2_X1 U3192 ( .A1(n4209), .A2(n4210), .ZN(n3705) );
  NAND2_X1 U3193 ( .A1(n4211), .A2(n4025), .ZN(n4210) );
  NAND2_X1 U3194 ( .A1(n4212), .A2(n4213), .ZN(n4211) );
  NAND2_X1 U3195 ( .A1(G3548), .A2(n4028), .ZN(n4213) );
  NAND2_X1 U3196 ( .A1(G3546), .A2(G265), .ZN(n4212) );
  NAND2_X1 U3197 ( .A1(n4214), .A2(G400), .ZN(n4209) );
  NAND2_X1 U3198 ( .A1(n4215), .A2(n4216), .ZN(n4214) );
  NAND2_X1 U3199 ( .A1(G265), .A2(n3678), .ZN(n4216) );
  NAND2_X1 U3200 ( .A1(n4028), .A2(n4200), .ZN(n4215) );
  AND2_X1 U3201 ( .A1(n4217), .A2(n4218), .ZN(n3724) );
  NAND2_X1 U3202 ( .A1(n4219), .A2(n4003), .ZN(n4218) );
  NAND2_X1 U3203 ( .A1(n4220), .A2(n4221), .ZN(n4219) );
  NAND2_X1 U3204 ( .A1(G3548), .A2(n4006), .ZN(n4221) );
  NAND2_X1 U3205 ( .A1(G3546), .A2(G273), .ZN(n4220) );
  NAND2_X1 U3206 ( .A1(n4222), .A2(G411), .ZN(n4217) );
  NAND2_X1 U3207 ( .A1(n4223), .A2(n4224), .ZN(n4222) );
  NAND2_X1 U3208 ( .A1(G273), .A2(n3678), .ZN(n4224) );
  NAND2_X1 U3209 ( .A1(n4006), .A2(n4200), .ZN(n4223) );
  NOR2_X1 U3210 ( .A1(KEYINPUT44), .A2(n4225), .ZN(n4189) );
  NOR4_X1 U3211 ( .A1(n4150), .A2(n4134), .A3(n4116), .A4(n4107), .ZN(n4225) );
  AND2_X1 U3212 ( .A1(n4226), .A2(n4227), .ZN(n4107) );
  NAND2_X1 U3213 ( .A1(n4228), .A2(n4071), .ZN(n4227) );
  NAND2_X1 U3214 ( .A1(n4229), .A2(n4230), .ZN(n4228) );
  NAND2_X1 U3215 ( .A1(G3548), .A2(n4074), .ZN(n4230) );
  NAND2_X1 U3216 ( .A1(G3546), .A2(G210), .ZN(n4229) );
  NAND2_X1 U3217 ( .A1(n4231), .A2(G457), .ZN(n4226) );
  NAND2_X1 U3218 ( .A1(n4232), .A2(n4233), .ZN(n4231) );
  NAND2_X1 U3219 ( .A1(G210), .A2(n3678), .ZN(n4233) );
  NAND2_X1 U3220 ( .A1(n4074), .A2(n4200), .ZN(n4232) );
  AND2_X1 U3221 ( .A1(n4234), .A2(n4235), .ZN(n4116) );
  NAND2_X1 U3222 ( .A1(n4236), .A2(n4061), .ZN(n4235) );
  NAND2_X1 U3223 ( .A1(n4237), .A2(n4238), .ZN(n4236) );
  NAND2_X1 U3224 ( .A1(G3548), .A2(n4064), .ZN(n4238) );
  NAND2_X1 U3225 ( .A1(G3546), .A2(G218), .ZN(n4237) );
  NAND2_X1 U3226 ( .A1(n4239), .A2(G468), .ZN(n4234) );
  NAND2_X1 U3227 ( .A1(n4240), .A2(n4241), .ZN(n4239) );
  NAND2_X1 U3228 ( .A1(G218), .A2(n3678), .ZN(n4241) );
  NAND2_X1 U3229 ( .A1(n4064), .A2(n4200), .ZN(n4240) );
  AND2_X1 U3230 ( .A1(n4242), .A2(n4243), .ZN(n4134) );
  NAND2_X1 U3231 ( .A1(n4244), .A2(n4015), .ZN(n4243) );
  INV_X1 U3232 ( .A(G422), .ZN(n4015) );
  NAND2_X1 U3233 ( .A1(n4245), .A2(n4246), .ZN(n4244) );
  NAND2_X1 U3234 ( .A1(G3548), .A2(n4018), .ZN(n4246) );
  NAND2_X1 U3235 ( .A1(G226), .A2(G3546), .ZN(n4245) );
  NAND2_X1 U3236 ( .A1(n4247), .A2(G422), .ZN(n4242) );
  NAND2_X1 U3237 ( .A1(n4248), .A2(n4249), .ZN(n4247) );
  NAND2_X1 U3238 ( .A1(G226), .A2(n3678), .ZN(n4249) );
  NAND2_X1 U3239 ( .A1(n4018), .A2(n4200), .ZN(n4248) );
  AND2_X1 U3240 ( .A1(n4250), .A2(n4251), .ZN(n4150) );
  NAND2_X1 U3241 ( .A1(n4252), .A2(n3993), .ZN(n4251) );
  NAND2_X1 U3242 ( .A1(n4253), .A2(n4254), .ZN(n4252) );
  NAND2_X1 U3243 ( .A1(G3548), .A2(n3996), .ZN(n4254) );
  NAND2_X1 U3244 ( .A1(G234), .A2(G3546), .ZN(n4253) );
  NAND2_X1 U3245 ( .A1(n4255), .A2(G435), .ZN(n4250) );
  NAND2_X1 U3246 ( .A1(n4256), .A2(n4257), .ZN(n4255) );
  NAND2_X1 U3247 ( .A1(G234), .A2(n3678), .ZN(n4257) );
  NAND2_X1 U3248 ( .A1(n3996), .A2(n4200), .ZN(n4256) );
  INV_X1 U3249 ( .A(G234), .ZN(n3996) );
  AND2_X1 U3250 ( .A1(n4258), .A2(n4259), .ZN(n3982) );
  NAND2_X1 U3251 ( .A1(n4260), .A2(n4261), .ZN(n4259) );
  INV_X1 U3252 ( .A(G446), .ZN(n4261) );
  NAND2_X1 U3253 ( .A1(n4262), .A2(n4263), .ZN(n4260) );
  NAND2_X1 U3254 ( .A1(G206), .A2(n3851), .ZN(n4263) );
  NAND2_X1 U3255 ( .A1(n4264), .A2(n3849), .ZN(n4262) );
  NAND2_X1 U3256 ( .A1(n4265), .A2(G446), .ZN(n4258) );
  NAND2_X1 U3257 ( .A1(n4266), .A2(n4267), .ZN(n4265) );
  NAND2_X1 U3258 ( .A1(G251), .A2(n4264), .ZN(n4267) );
  INV_X1 U3259 ( .A(G206), .ZN(n4264) );
  NAND2_X1 U3260 ( .A1(G206), .A2(G248), .ZN(n4266) );
  INV_X1 U3261 ( .A(G549), .ZN(G606) );
  INV_X1 U3262 ( .A(G545), .ZN(G594) );
  NOR2_X1 U3263 ( .A1(G850), .A2(G849), .ZN(G601) );
  INV_X1 U3264 ( .A(G552), .ZN(G849) );
  INV_X1 U3265 ( .A(G562), .ZN(G850) );
  INV_X1 U3266 ( .A(G366), .ZN(G600) );
  OR2_X1 U3267 ( .A1(n4268), .A2(KEYINPUT2), .ZN(G598_enc) );
  NOR3_X1 U3268 ( .A1(n3734), .A2(n4269), .A3(n4270), .ZN(n4268) );
  NOR2_X1 U3269 ( .A1(n4271), .A2(KEYINPUT69), .ZN(n4270) );
  NOR4_X1 U3270 ( .A1(n3855), .A2(n3836), .A3(n3453), .A4(n3856), .ZN(n4271) );
  NAND2_X1 U3271 ( .A1(n4272), .A2(n4273), .ZN(n3856) );
  OR2_X1 U3272 ( .A1(G251), .A2(G302), .ZN(n4273) );
  NAND2_X1 U3273 ( .A1(G302), .A2(n3842), .ZN(n4272) );
  NAND2_X1 U3274 ( .A1(n4274), .A2(n4275), .ZN(n3453) );
  OR2_X1 U3275 ( .A1(n3849), .A2(G293), .ZN(n4275) );
  NAND2_X1 U3276 ( .A1(G293), .A2(G242), .ZN(n4274) );
  AND2_X1 U3277 ( .A1(n4276), .A2(n4277), .ZN(n3836) );
  NAND2_X1 U3278 ( .A1(n4278), .A2(n4279), .ZN(n4277) );
  INV_X1 U3279 ( .A(G479), .ZN(n4279) );
  NAND2_X1 U3280 ( .A1(n4280), .A2(n4281), .ZN(n4278) );
  NAND2_X1 U3281 ( .A1(n3849), .A2(n4282), .ZN(n4281) );
  NAND2_X1 U3282 ( .A1(G308), .A2(n3851), .ZN(n4280) );
  NAND2_X1 U3283 ( .A1(n4283), .A2(G479), .ZN(n4276) );
  NAND2_X1 U3284 ( .A1(n4284), .A2(n4285), .ZN(n4283) );
  NAND2_X1 U3285 ( .A1(G251), .A2(n4282), .ZN(n4285) );
  INV_X1 U3286 ( .A(G308), .ZN(n4282) );
  NAND2_X1 U3287 ( .A1(G308), .A2(G248), .ZN(n4284) );
  AND2_X1 U3288 ( .A1(n4286), .A2(n4287), .ZN(n3855) );
  NAND2_X1 U3289 ( .A1(n4288), .A2(n4289), .ZN(n4287) );
  NAND2_X1 U3290 ( .A1(n4290), .A2(n4291), .ZN(n4288) );
  NAND2_X1 U3291 ( .A1(n3849), .A2(n4292), .ZN(n4291) );
  INV_X1 U3292 ( .A(G254), .ZN(n3849) );
  NAND2_X1 U3293 ( .A1(G316), .A2(n3851), .ZN(n4290) );
  INV_X1 U3294 ( .A(G242), .ZN(n3851) );
  NAND2_X1 U3295 ( .A1(n4293), .A2(G490), .ZN(n4286) );
  NAND2_X1 U3296 ( .A1(n4294), .A2(n4295), .ZN(n4293) );
  NAND2_X1 U3297 ( .A1(G251), .A2(n4292), .ZN(n4295) );
  NAND2_X1 U3298 ( .A1(G316), .A2(G248), .ZN(n4294) );
  NOR2_X1 U3299 ( .A1(KEYINPUT61), .A2(n4296), .ZN(n4269) );
  NOR4_X1 U3300 ( .A1(n4297), .A2(n4155), .A3(n4298), .A4(n4299), .ZN(n4296) );
  NOR2_X1 U3301 ( .A1(G514), .A2(G3546), .ZN(n4299) );
  NOR2_X1 U3302 ( .A1(n3679), .A2(n3678), .ZN(n4298) );
  AND2_X1 U3303 ( .A1(n4300), .A2(n4301), .ZN(n4155) );
  NAND2_X1 U3304 ( .A1(n4302), .A2(n3863), .ZN(n4301) );
  INV_X1 U3305 ( .A(G503), .ZN(n3863) );
  NAND2_X1 U3306 ( .A1(n4303), .A2(n4304), .ZN(n4302) );
  NAND2_X1 U3307 ( .A1(G3548), .A2(n3866), .ZN(n4304) );
  NAND2_X1 U3308 ( .A1(G324), .A2(G3546), .ZN(n4303) );
  NAND2_X1 U3309 ( .A1(n4305), .A2(G503), .ZN(n4300) );
  NAND2_X1 U3310 ( .A1(n4306), .A2(n4307), .ZN(n4305) );
  NAND2_X1 U3311 ( .A1(G324), .A2(n3678), .ZN(n4307) );
  INV_X1 U3312 ( .A(G3552), .ZN(n3678) );
  NAND2_X1 U3313 ( .A1(n3866), .A2(n4200), .ZN(n4306) );
  INV_X1 U3314 ( .A(G3550), .ZN(n4200) );
  INV_X1 U3315 ( .A(G324), .ZN(n3866) );
  NAND2_X1 U3316 ( .A1(n4308), .A2(n4309), .ZN(n4297) );
  NAND2_X1 U3317 ( .A1(n3698), .A2(n3699), .ZN(n4309) );
  NAND3_X1 U3318 ( .A1(n4310), .A2(n4311), .A3(G523), .ZN(n3699) );
  NAND2_X1 U3319 ( .A1(G3550), .A2(n3877), .ZN(n4311) );
  NAND2_X1 U3320 ( .A1(G3552), .A2(G341), .ZN(n4310) );
  NAND3_X1 U3321 ( .A1(n4312), .A2(n4313), .A3(n3874), .ZN(n3698) );
  NAND2_X1 U3322 ( .A1(G341), .A2(n4314), .ZN(n4313) );
  NAND2_X1 U3323 ( .A1(n3877), .A2(n4315), .ZN(n4312) );
  NAND2_X1 U3324 ( .A1(n3715), .A2(n3716), .ZN(n4308) );
  NAND3_X1 U3325 ( .A1(n4316), .A2(n4317), .A3(n3846), .ZN(n3716) );
  INV_X1 U3326 ( .A(G534), .ZN(n3846) );
  NAND2_X1 U3327 ( .A1(G351), .A2(n4314), .ZN(n4317) );
  INV_X1 U3328 ( .A(G3546), .ZN(n4314) );
  NAND2_X1 U3329 ( .A1(n3850), .A2(n4315), .ZN(n4316) );
  INV_X1 U3330 ( .A(G3548), .ZN(n4315) );
  NAND3_X1 U3331 ( .A1(n4318), .A2(n4319), .A3(G534), .ZN(n3715) );
  NAND2_X1 U3332 ( .A1(G3550), .A2(n3850), .ZN(n4319) );
  NAND2_X1 U3333 ( .A1(G351), .A2(G3552), .ZN(n4318) );
  NAND2_X1 U3334 ( .A1(n4320), .A2(n4321), .ZN(n3734) );
  OR2_X1 U3335 ( .A1(G251), .A2(G361), .ZN(n4321) );
  NAND2_X1 U3336 ( .A1(G361), .A2(n3842), .ZN(n4320) );
  INV_X1 U3337 ( .A(G248), .ZN(n3842) );
  INV_X1 U3338 ( .A(G299), .ZN(G593) );
  NAND3_X1 U3339 ( .A1(n4175), .A2(n4322), .A3(n4323), .ZN(G591) );
  NOR3_X1 U3340 ( .A1(KEYINPUT13), .A2(KEYINPUT47), .A3(KEYINPUT21), .ZN(n4323) );
  NAND2_X1 U3341 ( .A1(n4324), .A2(n4325), .ZN(n4322) );
  INV_X1 U3342 ( .A(n3955), .ZN(n4325) );
  NOR4_X1 U3343 ( .A1(KEYINPUT11), .A2(n4326), .A3(KEYINPUT56), .A4(KEYINPUT25), .ZN(n3955) );
  OR2_X1 U3344 ( .A1(n4180), .A2(KEYINPUT39), .ZN(n4324) );
  AND2_X1 U3345 ( .A1(n4327), .A2(n4328), .ZN(n4175) );
  NAND2_X1 U3346 ( .A1(n3952), .A2(n4329), .ZN(n4328) );
  NAND2_X1 U3347 ( .A1(G446), .A2(n4330), .ZN(n4327) );
  OR2_X1 U3348 ( .A1(n4331), .A2(KEYINPUT0), .ZN(G588_enc) );
  NOR2_X1 U3349 ( .A1(n3958), .A2(n4332), .ZN(n4331) );
  NOR2_X1 U3350 ( .A1(n4180), .A2(KEYINPUT39), .ZN(n4332) );
  NOR2_X1 U3351 ( .A1(n3949), .A2(n3944), .ZN(n4180) );
  NAND3_X1 U3352 ( .A1(n3952), .A2(n3945), .A3(n3934), .ZN(n3949) );
  NOR2_X1 U3353 ( .A1(n4333), .A2(KEYINPUT17), .ZN(n3958) );
  OR2_X1 U3354 ( .A1(n4334), .A2(KEYINPUT7), .ZN(G585_enc) );
  NOR4_X1 U3355 ( .A1(n4335), .A2(n4336), .A3(n3777), .A4(n3804), .ZN(n4334) );
  OR3_X1 U3356 ( .A1(n3674), .A2(n3700), .A3(n4154), .ZN(n4336) );
  XOR2_X1 U3357 ( .A(n4337), .B(n3783), .Z(n4154) );
  NAND3_X1 U3358 ( .A1(n4338), .A2(n3772), .A3(n4339), .ZN(n4337) );
  NOR3_X1 U3359 ( .A1(KEYINPUT35), .A2(KEYINPUT63), .A3(KEYINPUT41), .ZN(n4339) );
  NAND2_X1 U3360 ( .A1(n3775), .A2(n4340), .ZN(n4338) );
  AND2_X1 U3361 ( .A1(n4341), .A2(n4342), .ZN(n3700) );
  OR2_X1 U3362 ( .A1(n4343), .A2(n3789), .ZN(n4342) );
  XOR2_X1 U3363 ( .A(n3788), .B(n4344), .Z(n3674) );
  NOR2_X1 U3364 ( .A1(KEYINPUT70), .A2(n4340), .ZN(n4344) );
  NAND2_X1 U3365 ( .A1(n3768), .A2(n4341), .ZN(n4340) );
  NAND2_X1 U3366 ( .A1(n3789), .A2(n4343), .ZN(n4341) );
  NAND2_X1 U3367 ( .A1(n3755), .A2(n4345), .ZN(n4343) );
  NAND2_X1 U3368 ( .A1(n3718), .A2(G54), .ZN(n4345) );
  INV_X1 U3369 ( .A(n4346), .ZN(n3755) );
  OR4_X1 U3370 ( .A1(n3733), .A2(n4122), .A3(n4090), .A4(n4102), .ZN(n4335) );
  XOR2_X1 U3371 ( .A(n3800), .B(n4347), .Z(n4102) );
  NOR2_X1 U3372 ( .A1(n4348), .A2(n3797), .ZN(n4347) );
  NOR2_X1 U3373 ( .A1(n4139), .A2(n3802), .ZN(n4348) );
  INV_X1 U3374 ( .A(n3798), .ZN(n3802) );
  INV_X1 U3375 ( .A(G623), .ZN(n4090) );
  XNOR2_X1 U3376 ( .A(n3458), .B(n3460), .ZN(G623) );
  NOR3_X1 U3377 ( .A1(n4349), .A2(n4350), .A3(n3800), .ZN(n3460) );
  NAND2_X1 U3378 ( .A1(n4351), .A2(n4352), .ZN(n3800) );
  NAND2_X1 U3379 ( .A1(G302), .A2(n3423), .ZN(n4352) );
  NAND2_X1 U3380 ( .A1(G307), .A2(G332), .ZN(n4351) );
  NOR2_X1 U3381 ( .A1(n4353), .A2(n4354), .ZN(n4350) );
  NOR2_X1 U3382 ( .A1(KEYINPUT72), .A2(n3797), .ZN(n4353) );
  NOR2_X1 U3383 ( .A1(n4139), .A2(n4355), .ZN(n4349) );
  NOR3_X1 U3384 ( .A1(n3797), .A2(KEYINPUT71), .A3(n3798), .ZN(n4355) );
  NOR2_X1 U3385 ( .A1(n3804), .A2(n3806), .ZN(n3798) );
  NAND2_X1 U3386 ( .A1(n4356), .A2(n3805), .ZN(n3804) );
  NAND2_X1 U3387 ( .A1(n4357), .A2(n4358), .ZN(n3797) );
  NAND2_X1 U3388 ( .A1(n3827), .A2(n4359), .ZN(n4358) );
  NAND2_X1 U3389 ( .A1(G479), .A2(n3431), .ZN(n4357) );
  NAND2_X1 U3390 ( .A1(n4360), .A2(n4361), .ZN(n3458) );
  NAND2_X1 U3391 ( .A1(G293), .A2(n3423), .ZN(n4361) );
  NAND2_X1 U3392 ( .A1(G332), .A2(G299), .ZN(n4360) );
  NAND3_X1 U3393 ( .A1(n4362), .A2(n4363), .A3(n3801), .ZN(n4122) );
  OR2_X1 U3394 ( .A1(n3805), .A2(n3806), .ZN(n3801) );
  NAND3_X1 U3395 ( .A1(n4139), .A2(n4356), .A3(n4359), .ZN(n4363) );
  NAND2_X1 U3396 ( .A1(n3806), .A2(n4364), .ZN(n4362) );
  NAND2_X1 U3397 ( .A1(n4356), .A2(n4365), .ZN(n4364) );
  NAND2_X1 U3398 ( .A1(n3805), .A2(n4354), .ZN(n4365) );
  INV_X1 U3399 ( .A(n4139), .ZN(n4354) );
  NOR3_X1 U3400 ( .A1(KEYINPUT12), .A2(n4366), .A3(n4184), .ZN(n4139) );
  OR4_X1 U3401 ( .A1(KEYINPUT18), .A2(n4170), .A3(KEYINPUT62), .A4(KEYINPUT28),  .ZN(n4184) );
  NAND2_X1 U3402 ( .A1(n4367), .A2(n4368), .ZN(n4170) );
  NAND2_X1 U3403 ( .A1(n3783), .A2(n3759), .ZN(n4368) );
  NAND2_X1 U3404 ( .A1(n3772), .A2(n4369), .ZN(n3759) );
  NAND2_X1 U3405 ( .A1(n3775), .A2(n3756), .ZN(n4369) );
  NAND2_X1 U3406 ( .A1(n3768), .A2(n4370), .ZN(n3756) );
  NAND2_X1 U3407 ( .A1(n3789), .A2(n4346), .ZN(n4370) );
  NAND2_X1 U3408 ( .A1(n3778), .A2(n4371), .ZN(n4346) );
  NAND2_X1 U3409 ( .A1(n3718), .A2(n4372), .ZN(n4371) );
  INV_X1 U3410 ( .A(n3767), .ZN(n3789) );
  INV_X1 U3411 ( .A(n3788), .ZN(n3775) );
  NAND2_X1 U3412 ( .A1(G503), .A2(n3430), .ZN(n4367) );
  NOR2_X1 U3413 ( .A1(n4187), .A2(n4373), .ZN(n4366) );
  NOR2_X1 U3414 ( .A1(n4174), .A2(KEYINPUT31), .ZN(n4187) );
  AND4_X1 U3415 ( .A1(n3718), .A2(n3776), .A3(n3783), .A4(n3424), .ZN(n4174) );
  XOR2_X1 U3416 ( .A(G503), .B(n3430), .Z(n3783) );
  NAND2_X1 U3417 ( .A1(n4374), .A2(n4375), .ZN(n3430) );
  NAND2_X1 U3418 ( .A1(G324), .A2(n3423), .ZN(n4375) );
  NAND2_X1 U3419 ( .A1(G331), .A2(G332), .ZN(n4374) );
  NOR2_X1 U3420 ( .A1(n3788), .A2(n3767), .ZN(n3776) );
  NAND2_X1 U3421 ( .A1(n3768), .A2(n4376), .ZN(n3767) );
  NAND2_X1 U3422 ( .A1(n3432), .A2(n3874), .ZN(n4376) );
  INV_X1 U3423 ( .A(n3774), .ZN(n3768) );
  NOR2_X1 U3424 ( .A1(n3874), .A2(n3432), .ZN(n3774) );
  NAND2_X1 U3425 ( .A1(n4377), .A2(n4378), .ZN(n3432) );
  NAND2_X1 U3426 ( .A1(G332), .A2(G599), .ZN(n4378) );
  INV_X1 U3427 ( .A(G348), .ZN(G599) );
  NAND2_X1 U3428 ( .A1(n3423), .A2(n3877), .ZN(n4377) );
  INV_X1 U3429 ( .A(G523), .ZN(n3874) );
  NAND2_X1 U3430 ( .A1(n4379), .A2(n3772), .ZN(n3788) );
  NAND2_X1 U3431 ( .A1(G514), .A2(n3426), .ZN(n3772) );
  INV_X1 U3432 ( .A(n4380), .ZN(n3426) );
  NAND2_X1 U3433 ( .A1(n4380), .A2(n3679), .ZN(n4379) );
  INV_X1 U3434 ( .A(G514), .ZN(n3679) );
  NOR2_X1 U3435 ( .A1(n3423), .A2(G338), .ZN(n4380) );
  INV_X1 U3436 ( .A(n3777), .ZN(n3718) );
  NAND2_X1 U3437 ( .A1(n3778), .A2(n4381), .ZN(n3777) );
  OR2_X1 U3438 ( .A1(n3418), .A2(G534), .ZN(n4381) );
  NAND2_X1 U3439 ( .A1(G534), .A2(n3418), .ZN(n3778) );
  NAND2_X1 U3440 ( .A1(n4382), .A2(n4383), .ZN(n3418) );
  NAND2_X1 U3441 ( .A1(G351), .A2(n3423), .ZN(n4383) );
  NAND2_X1 U3442 ( .A1(G332), .A2(G358), .ZN(n4382) );
  NAND2_X1 U3443 ( .A1(n4384), .A2(n4289), .ZN(n3805) );
  INV_X1 U3444 ( .A(n3827), .ZN(n4356) );
  NOR2_X1 U3445 ( .A1(n4289), .A2(n4384), .ZN(n3827) );
  INV_X1 U3446 ( .A(n3433), .ZN(n4384) );
  NAND2_X1 U3447 ( .A1(n4385), .A2(n4386), .ZN(n3433) );
  NAND2_X1 U3448 ( .A1(G316), .A2(n3423), .ZN(n4386) );
  NAND2_X1 U3449 ( .A1(G323), .A2(G332), .ZN(n4385) );
  INV_X1 U3450 ( .A(G490), .ZN(n4289) );
  INV_X1 U3451 ( .A(n4359), .ZN(n3806) );
  XOR2_X1 U3452 ( .A(G479), .B(n3431), .Z(n4359) );
  NAND2_X1 U3453 ( .A1(n4387), .A2(n4388), .ZN(n3431) );
  NAND2_X1 U3454 ( .A1(G308), .A2(n3423), .ZN(n4388) );
  NAND2_X1 U3455 ( .A1(G315), .A2(G332), .ZN(n4387) );
  OR2_X1 U3456 ( .A1(n3719), .A2(n4389), .ZN(n3733) );
  NOR2_X1 U3457 ( .A1(n4373), .A2(n3424), .ZN(n4389) );
  INV_X1 U3458 ( .A(n4372), .ZN(n3424) );
  INV_X1 U3459 ( .A(G54), .ZN(n4373) );
  NOR2_X1 U3460 ( .A1(n4372), .A2(G54), .ZN(n3719) );
  NAND2_X1 U3461 ( .A1(n4390), .A2(n4391), .ZN(n4372) );
  NAND2_X1 U3462 ( .A1(G361), .A2(n3423), .ZN(n4391) );
  INV_X1 U3463 ( .A(G332), .ZN(n3423) );
  NAND2_X1 U3464 ( .A1(G332), .A2(G366), .ZN(n4390) );
  OR2_X1 U3465 ( .A1(n4392), .A2(KEYINPUT8), .ZN(G575_enc) );
  NOR4_X1 U3466 ( .A1(n4393), .A2(n4394), .A3(n4133), .A4(n4149), .ZN(n4392) );
  XOR2_X1 U3467 ( .A(n4395), .B(n3962), .Z(n4149) );
  NAND3_X1 U3468 ( .A1(n4396), .A2(n4397), .A3(n4398), .ZN(n4395) );
  NOR3_X1 U3469 ( .A1(KEYINPUT20), .A2(KEYINPUT52), .A3(KEYINPUT24), .ZN(n4398) );
  NAND2_X1 U3470 ( .A1(n4399), .A2(n3963), .ZN(n4397) );
  XNOR2_X1 U3471 ( .A(n3919), .B(n4400), .ZN(n4133) );
  OR3_X1 U3472 ( .A1(n3704), .A2(n3723), .A3(n3685), .ZN(n4394) );
  XOR2_X1 U3473 ( .A(n3900), .B(n4401), .Z(n3685) );
  NOR4_X1 U3474 ( .A1(KEYINPUT53), .A2(KEYINPUT46), .A3(n3890), .A4(n4399),  .ZN(n4401) );
  AND2_X1 U3475 ( .A1(n4402), .A2(n4403), .ZN(n4399) );
  XOR2_X1 U3476 ( .A(n3901), .B(n4404), .Z(n3723) );
  NOR2_X1 U3477 ( .A1(n4405), .A2(n4406), .ZN(n4404) );
  NOR2_X1 U3478 ( .A1(n3961), .A2(n4407), .ZN(n4405) );
  XOR2_X1 U3479 ( .A(n4403), .B(n4402), .Z(n3704) );
  NAND2_X1 U3480 ( .A1(n3893), .A2(n4408), .ZN(n4403) );
  NAND2_X1 U3481 ( .A1(G4), .A2(n3960), .ZN(n4408) );
  INV_X1 U3482 ( .A(n3976), .ZN(n3893) );
  OR4_X1 U3483 ( .A1(n3739), .A2(n4094), .A3(n4106), .A4(n4115), .ZN(n4393) );
  XOR2_X1 U3484 ( .A(n3953), .B(n4409), .Z(n4115) );
  NOR2_X1 U3485 ( .A1(n4410), .A2(n3931), .ZN(n4409) );
  NOR2_X1 U3486 ( .A1(n3946), .A2(n4400), .ZN(n4410) );
  XOR2_X1 U3487 ( .A(n3954), .B(n4411), .Z(n4106) );
  NOR2_X1 U3488 ( .A1(n4412), .A2(n3932), .ZN(n4411) );
  NOR3_X1 U3489 ( .A1(n3944), .A2(n4400), .A3(n3953), .ZN(n4412) );
  INV_X1 U3490 ( .A(n3919), .ZN(n3944) );
  XOR2_X1 U3491 ( .A(n3952), .B(n4413), .Z(n4094) );
  NOR2_X1 U3492 ( .A1(n4414), .A2(n4415), .ZN(n4413) );
  NOR3_X1 U3493 ( .A1(n4416), .A2(KEYINPUT50), .A3(n4329), .ZN(n4415) );
  INV_X1 U3494 ( .A(n4400), .ZN(n4416) );
  NOR3_X1 U3495 ( .A1(n4400), .A2(KEYINPUT49), .A3(n3941), .ZN(n4414) );
  NAND2_X1 U3496 ( .A1(n3925), .A2(n4417), .ZN(n3941) );
  NAND3_X1 U3497 ( .A1(n3934), .A2(n3945), .A3(n3919), .ZN(n4417) );
  NOR2_X1 U3498 ( .A1(n3946), .A2(n3931), .ZN(n3919) );
  NOR2_X1 U3499 ( .A1(n4418), .A2(G422), .ZN(n3946) );
  INV_X1 U3500 ( .A(n4329), .ZN(n3925) );
  NAND2_X1 U3501 ( .A1(n3927), .A2(n4419), .ZN(n4329) );
  NAND2_X1 U3502 ( .A1(n3934), .A2(n3932), .ZN(n4419) );
  NAND2_X1 U3503 ( .A1(n4420), .A2(n4421), .ZN(n3932) );
  NAND2_X1 U3504 ( .A1(n3931), .A2(n3945), .ZN(n4421) );
  INV_X1 U3505 ( .A(n3953), .ZN(n3945) );
  NAND2_X1 U3506 ( .A1(n4420), .A2(n4422), .ZN(n3953) );
  NAND2_X1 U3507 ( .A1(n4423), .A2(n4061), .ZN(n4422) );
  AND2_X1 U3508 ( .A1(G422), .A2(n4418), .ZN(n3931) );
  INV_X1 U3509 ( .A(n3933), .ZN(n4420) );
  NOR2_X1 U3510 ( .A1(n4061), .A2(n4423), .ZN(n3933) );
  INV_X1 U3511 ( .A(G468), .ZN(n4061) );
  INV_X1 U3512 ( .A(n3954), .ZN(n3934) );
  NAND2_X1 U3513 ( .A1(n3927), .A2(n4424), .ZN(n3954) );
  NAND2_X1 U3514 ( .A1(n4425), .A2(n4071), .ZN(n4424) );
  OR2_X1 U3515 ( .A1(n4071), .A2(n4425), .ZN(n3927) );
  INV_X1 U3516 ( .A(G457), .ZN(n4071) );
  NOR3_X1 U3517 ( .A1(KEYINPUT9), .A2(n4426), .A3(n4179), .ZN(n4400) );
  OR4_X1 U3518 ( .A1(KEYINPUT10), .A2(n4326), .A3(KEYINPUT51), .A4(KEYINPUT23),  .ZN(n4179) );
  NAND2_X1 U3519 ( .A1(n4427), .A2(n4428), .ZN(n4326) );
  NAND2_X1 U3520 ( .A1(n3962), .A2(n3968), .ZN(n4428) );
  NAND2_X1 U3521 ( .A1(n4396), .A2(n4429), .ZN(n3968) );
  NAND2_X1 U3522 ( .A1(n3967), .A2(n3976), .ZN(n4429) );
  NAND2_X1 U3523 ( .A1(n3903), .A2(n4430), .ZN(n3976) );
  NAND2_X1 U3524 ( .A1(n4406), .A2(n3974), .ZN(n4430) );
  INV_X1 U3525 ( .A(n3901), .ZN(n3974) );
  INV_X1 U3526 ( .A(n3898), .ZN(n4396) );
  NAND2_X1 U3527 ( .A1(n4431), .A2(n4432), .ZN(n3898) );
  NAND2_X1 U3528 ( .A1(n3890), .A2(n3963), .ZN(n4432) );
  NAND2_X1 U3529 ( .A1(G389), .A2(n4433), .ZN(n4431) );
  NAND2_X1 U3530 ( .A1(G435), .A2(n4434), .ZN(n4427) );
  NOR2_X1 U3531 ( .A1(n4164), .A2(n4407), .ZN(n4426) );
  NOR2_X1 U3532 ( .A1(n4333), .A2(KEYINPUT16), .ZN(n4164) );
  AND3_X1 U3533 ( .A1(n3962), .A2(n3967), .A3(n3960), .ZN(n4333) );
  NOR2_X1 U3534 ( .A1(n3961), .A2(n3901), .ZN(n3960) );
  NAND2_X1 U3535 ( .A1(n3903), .A2(n4435), .ZN(n3901) );
  NAND2_X1 U3536 ( .A1(n4436), .A2(n4003), .ZN(n4435) );
  OR2_X1 U3537 ( .A1(n4003), .A2(n4436), .ZN(n3903) );
  INV_X1 U3538 ( .A(G411), .ZN(n4003) );
  NOR2_X1 U3539 ( .A1(n3902), .A2(n3900), .ZN(n3967) );
  INV_X1 U3540 ( .A(n3963), .ZN(n3900) );
  XOR2_X1 U3541 ( .A(G389), .B(n4433), .Z(n3963) );
  INV_X1 U3542 ( .A(n4402), .ZN(n3902) );
  NOR2_X1 U3543 ( .A1(n4437), .A2(n3890), .ZN(n4402) );
  NOR2_X1 U3544 ( .A1(n4025), .A2(n4438), .ZN(n3890) );
  AND2_X1 U3545 ( .A1(n4438), .A2(n4025), .ZN(n4437) );
  INV_X1 U3546 ( .A(G400), .ZN(n4025) );
  XNOR2_X1 U3547 ( .A(n3993), .B(n4434), .ZN(n3962) );
  INV_X1 U3548 ( .A(G435), .ZN(n3993) );
  XOR2_X1 U3549 ( .A(G446), .B(n4330), .Z(n3952) );
  XOR2_X1 U3550 ( .A(n3961), .B(n4407), .Z(n3739) );
  INV_X1 U3551 ( .A(G4), .ZN(n4407) );
  NAND2_X1 U3552 ( .A1(n3977), .A2(n3895), .ZN(n3961) );
  INV_X1 U3553 ( .A(n4406), .ZN(n3895) );
  NOR2_X1 U3554 ( .A1(n4039), .A2(n4439), .ZN(n4406) );
  NAND2_X1 U3555 ( .A1(n4439), .A2(n4039), .ZN(n3977) );
  INV_X1 U3556 ( .A(G374), .ZN(n4039) );
  XNOR2_X1 U3557 ( .A(n4440), .B(n4441), .ZN(G1004) );
  XNOR2_X1 U3558 ( .A(n4006), .B(G265), .ZN(n4441) );
  XOR2_X1 U3559 ( .A(n4442), .B(n4443), .Z(n4440) );
  XOR2_X1 U3560 ( .A(n4444), .B(n4445), .Z(n4443) );
  XNOR2_X1 U3561 ( .A(n4074), .B(G206), .ZN(n4445) );
  XNOR2_X1 U3562 ( .A(n4018), .B(G218), .ZN(n4444) );
  INV_X1 U3563 ( .A(G226), .ZN(n4018) );
  XOR2_X1 U3564 ( .A(n4446), .B(n4447), .Z(n4442) );
  XNOR2_X1 U3565 ( .A(n4052), .B(G234), .ZN(n4447) );
  INV_X1 U3566 ( .A(G257), .ZN(n4052) );
  XNOR2_X1 U3567 ( .A(G289), .B(G281), .ZN(n4446) );
  XOR2_X1 U3568 ( .A(n4448), .B(G369), .Z(G1002) );
  XOR2_X1 U3569 ( .A(n4449), .B(n4450), .Z(n4448) );
  XOR2_X1 U3570 ( .A(n4451), .B(n4452), .Z(n4450) );
  XNOR2_X1 U3571 ( .A(n3877), .B(G324), .ZN(n4452) );
  INV_X1 U3572 ( .A(G341), .ZN(n3877) );
  XNOR2_X1 U3573 ( .A(G361), .B(n3850), .ZN(n4451) );
  INV_X1 U3574 ( .A(G351), .ZN(n3850) );
  XOR2_X1 U3575 ( .A(n4453), .B(n4454), .Z(n4449) );
  XNOR2_X1 U3576 ( .A(n4292), .B(G308), .ZN(n4454) );
  INV_X1 U3577 ( .A(G316), .ZN(n4292) );
  XNOR2_X1 U3578 ( .A(G293), .B(G302), .ZN(n4453) );
  XOR2_X1 U3579 ( .A(n4455), .B(n4456), .Z(G1000) );
  XNOR2_X1 U3580 ( .A(n4439), .B(n4457), .ZN(n4456) );
  XOR2_X1 U3581 ( .A(n4436), .B(n4458), .Z(n4457) );
  NOR2_X1 U3582 ( .A1(KEYINPUT96), .A2(n4459), .ZN(n4458) );
  XOR2_X1 U3583 ( .A(n4460), .B(n4461), .Z(n4459) );
  XOR2_X1 U3584 ( .A(n4418), .B(n4462), .Z(n4461) );
  NAND2_X1 U3585 ( .A1(n4463), .A2(n4464), .ZN(n4462) );
  NAND2_X1 U3586 ( .A1(n4465), .A2(n4466), .ZN(n4464) );
  XOR2_X1 U3587 ( .A(G289), .B(n4467), .Z(n4465) );
  NAND2_X1 U3588 ( .A1(n4468), .A2(G335), .ZN(n4463) );
  XOR2_X1 U3589 ( .A(G292), .B(n4467), .Z(n4468) );
  XOR2_X1 U3590 ( .A(n4330), .B(n4434), .Z(n4467) );
  NAND2_X1 U3591 ( .A1(n4469), .A2(n4470), .ZN(n4434) );
  NAND2_X1 U3592 ( .A1(G234), .A2(n4466), .ZN(n4470) );
  NAND2_X1 U3593 ( .A1(G241), .A2(G335), .ZN(n4469) );
  NAND2_X1 U3594 ( .A1(n4471), .A2(n4472), .ZN(n4330) );
  NAND2_X1 U3595 ( .A1(G206), .A2(n4466), .ZN(n4472) );
  NAND2_X1 U3596 ( .A1(G209), .A2(G335), .ZN(n4471) );
  NAND2_X1 U3597 ( .A1(n4473), .A2(n4474), .ZN(n4418) );
  NAND2_X1 U3598 ( .A1(G226), .A2(n4466), .ZN(n4474) );
  NAND2_X1 U3599 ( .A1(G233), .A2(G335), .ZN(n4473) );
  XOR2_X1 U3600 ( .A(n4425), .B(n4423), .Z(n4460) );
  NAND2_X1 U3601 ( .A1(n4475), .A2(n4476), .ZN(n4423) );
  OR2_X1 U3602 ( .A1(G225), .A2(n4466), .ZN(n4476) );
  NAND2_X1 U3603 ( .A1(n4064), .A2(n4466), .ZN(n4475) );
  INV_X1 U3604 ( .A(G218), .ZN(n4064) );
  NAND2_X1 U3605 ( .A1(n4477), .A2(n4478), .ZN(n4425) );
  OR2_X1 U3606 ( .A1(G217), .A2(n4466), .ZN(n4478) );
  NAND2_X1 U3607 ( .A1(n4074), .A2(n4466), .ZN(n4477) );
  INV_X1 U3608 ( .A(G210), .ZN(n4074) );
  NAND2_X1 U3609 ( .A1(n4479), .A2(n4480), .ZN(n4436) );
  OR2_X1 U3610 ( .A1(G280), .A2(n4466), .ZN(n4480) );
  NAND2_X1 U3611 ( .A1(n4006), .A2(n4466), .ZN(n4479) );
  INV_X1 U3612 ( .A(G273), .ZN(n4006) );
  AND2_X1 U3613 ( .A1(n4481), .A2(n4482), .ZN(n4439) );
  NAND2_X1 U3614 ( .A1(G281), .A2(n4466), .ZN(n4482) );
  NAND2_X1 U3615 ( .A1(G288), .A2(G335), .ZN(n4481) );
  XNOR2_X1 U3616 ( .A(n4438), .B(n4433), .ZN(n4455) );
  NAND2_X1 U3617 ( .A1(n4483), .A2(n4484), .ZN(n4433) );
  NAND2_X1 U3618 ( .A1(G257), .A2(n4466), .ZN(n4484) );
  NAND2_X1 U3619 ( .A1(G264), .A2(G335), .ZN(n4483) );
  NAND2_X1 U3620 ( .A1(n4485), .A2(n4486), .ZN(n4438) );
  OR2_X1 U3621 ( .A1(G272), .A2(n4466), .ZN(n4486) );
  NAND2_X1 U3622 ( .A1(n4028), .A2(n4466), .ZN(n4485) );
  INV_X1 U3623 ( .A(G335), .ZN(n4466) );
  INV_X1 U3624 ( .A(G265), .ZN(n4028) );
endmodule

