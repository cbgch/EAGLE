//Key = 1010000000010110000111010111001110110011111111100011100011101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U752 ( .A(n1044), .B(n1045), .Z(G9) );
NAND2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U755 ( .A1(G953), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1049) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR4_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1057) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
XOR2_X1 U761 ( .A(n1065), .B(KEYINPUT53), .Z(n1063) );
NOR3_X1 U762 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1070), .A2(n1059), .ZN(n1069) );
NOR2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1060), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1046), .ZN(n1077) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1081), .ZN(n1068) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1058), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1060), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
XOR2_X1 U776 ( .A(n1088), .B(KEYINPUT41), .Z(n1086) );
AND2_X1 U777 ( .A1(n1089), .A2(n1058), .ZN(n1076) );
NAND2_X1 U778 ( .A1(n1090), .A2(n1080), .ZN(n1089) );
INV_X1 U779 ( .A(KEYINPUT57), .ZN(n1080) );
NOR3_X1 U780 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1050) );
NOR3_X1 U782 ( .A1(n1095), .A2(n1096), .A3(n1066), .ZN(n1094) );
INV_X1 U783 ( .A(n1064), .ZN(n1066) );
NAND3_X1 U784 ( .A1(n1097), .A2(n1098), .A3(n1087), .ZN(n1095) );
NOR3_X1 U785 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1093) );
XOR2_X1 U786 ( .A(n1102), .B(n1103), .Z(n1101) );
XNOR2_X1 U787 ( .A(n1104), .B(KEYINPUT39), .ZN(n1102) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1107), .B(G469), .Z(n1092) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1091) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(G72) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1113), .ZN(n1117) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND3_X1 U797 ( .A1(G900), .A2(n1120), .A3(G953), .ZN(n1116) );
XOR2_X1 U798 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(n1121) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U801 ( .A1(n1127), .A2(n1113), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1125) );
NAND2_X1 U804 ( .A1(n1132), .A2(n1113), .ZN(n1131) );
XOR2_X1 U805 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
XOR2_X1 U807 ( .A(KEYINPUT24), .B(n1137), .Z(n1136) );
NAND3_X1 U808 ( .A1(G898), .A2(n1138), .A3(G953), .ZN(n1130) );
NOR2_X1 U809 ( .A1(n1139), .A2(n1140), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
NOR3_X1 U811 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
NOR2_X1 U812 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
NOR2_X1 U813 ( .A1(n1149), .A2(n1145), .ZN(n1148) );
INV_X1 U814 ( .A(n1144), .ZN(n1147) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1150), .ZN(G63) );
XNOR2_X1 U816 ( .A(n1151), .B(n1152), .ZN(n1150) );
AND2_X1 U817 ( .A1(G478), .A2(n1153), .ZN(n1152) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1154), .ZN(G60) );
XOR2_X1 U819 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U820 ( .A1(n1106), .A2(n1146), .ZN(n1155) );
XOR2_X1 U821 ( .A(n1157), .B(G104), .Z(G6) );
NAND2_X1 U822 ( .A1(KEYINPUT61), .A2(n1158), .ZN(n1157) );
NAND2_X1 U823 ( .A1(n1159), .A2(n1047), .ZN(n1158) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1160), .ZN(G57) );
XOR2_X1 U825 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U826 ( .A(G101), .B(n1163), .ZN(n1162) );
NAND2_X1 U827 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
NAND3_X1 U828 ( .A1(n1153), .A2(G472), .A3(n1166), .ZN(n1165) );
NAND2_X1 U829 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
INV_X1 U830 ( .A(n1166), .ZN(n1168) );
XNOR2_X1 U831 ( .A(n1169), .B(n1170), .ZN(n1166) );
XNOR2_X1 U832 ( .A(n1171), .B(n1172), .ZN(n1169) );
NOR2_X1 U833 ( .A1(KEYINPUT1), .A2(n1173), .ZN(n1172) );
XOR2_X1 U834 ( .A(KEYINPUT58), .B(n1174), .Z(n1167) );
AND2_X1 U835 ( .A1(G472), .A2(n1153), .ZN(n1174) );
NOR2_X1 U836 ( .A1(n1139), .A2(n1175), .ZN(G54) );
XOR2_X1 U837 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U838 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U839 ( .A(KEYINPUT8), .B(n1180), .Z(n1179) );
NOR2_X1 U840 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U841 ( .A(KEYINPUT28), .B(n1183), .Z(n1182) );
NOR2_X1 U842 ( .A1(G110), .A2(n1184), .ZN(n1183) );
NOR2_X1 U843 ( .A1(G140), .A2(n1185), .ZN(n1181) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1146), .ZN(n1178) );
XOR2_X1 U845 ( .A(n1187), .B(n1123), .Z(n1176) );
NOR2_X1 U846 ( .A1(n1139), .A2(n1188), .ZN(G51) );
XOR2_X1 U847 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR4_X1 U848 ( .A1(n1191), .A2(n1192), .A3(KEYINPUT48), .A4(n1193), .ZN(n1190) );
AND2_X1 U849 ( .A1(n1194), .A2(KEYINPUT22), .ZN(n1193) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1138), .ZN(n1192) );
NOR2_X1 U851 ( .A1(n1194), .A2(n1196), .ZN(n1195) );
NOR4_X1 U852 ( .A1(n1134), .A2(n1196), .A3(KEYINPUT22), .A4(n1194), .ZN(n1191) );
XNOR2_X1 U853 ( .A(n1197), .B(n1198), .ZN(n1194) );
XOR2_X1 U854 ( .A(n1199), .B(KEYINPUT10), .Z(n1197) );
NAND2_X1 U855 ( .A1(KEYINPUT13), .A2(n1200), .ZN(n1199) );
INV_X1 U856 ( .A(KEYINPUT42), .ZN(n1196) );
INV_X1 U857 ( .A(n1138), .ZN(n1134) );
NAND2_X1 U858 ( .A1(n1153), .A2(n1103), .ZN(n1189) );
INV_X1 U859 ( .A(n1146), .ZN(n1153) );
NAND2_X1 U860 ( .A1(G902), .A2(n1052), .ZN(n1146) );
INV_X1 U861 ( .A(n1149), .ZN(n1052) );
NOR3_X1 U862 ( .A1(n1119), .A2(n1137), .A3(n1135), .ZN(n1149) );
NAND3_X1 U863 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1135) );
AND3_X1 U864 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NAND2_X1 U865 ( .A1(n1061), .A2(n1207), .ZN(n1202) );
NAND2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U867 ( .A(KEYINPUT43), .B(n1210), .Z(n1209) );
NOR3_X1 U868 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
INV_X1 U869 ( .A(n1075), .ZN(n1212) );
XOR2_X1 U870 ( .A(KEYINPUT25), .B(n1085), .Z(n1211) );
XNOR2_X1 U871 ( .A(KEYINPUT56), .B(n1214), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1047), .A2(n1215), .ZN(n1201) );
NAND2_X1 U873 ( .A1(n1216), .A2(n1079), .ZN(n1215) );
XOR2_X1 U874 ( .A(n1217), .B(KEYINPUT6), .Z(n1216) );
AND3_X1 U875 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1047) );
NAND4_X1 U876 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1119) );
AND4_X1 U877 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NOR2_X1 U878 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
NOR2_X1 U879 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U880 ( .A(n1233), .B(KEYINPUT15), .Z(n1231) );
NOR3_X1 U881 ( .A1(n1234), .A2(n1235), .A3(n1060), .ZN(n1229) );
NOR2_X1 U882 ( .A1(n1113), .A2(G952), .ZN(n1139) );
XNOR2_X1 U883 ( .A(G146), .B(n1221), .ZN(G48) );
NAND4_X1 U884 ( .A1(n1159), .A2(n1218), .A3(n1236), .A4(n1237), .ZN(n1221) );
XOR2_X1 U885 ( .A(n1238), .B(n1222), .Z(G45) );
NAND3_X1 U886 ( .A1(n1218), .A2(n1075), .A3(n1239), .ZN(n1222) );
AND3_X1 U887 ( .A1(n1099), .A2(n1240), .A3(n1237), .ZN(n1239) );
XOR2_X1 U888 ( .A(G140), .B(n1241), .Z(G42) );
NOR2_X1 U889 ( .A1(KEYINPUT49), .A2(n1228), .ZN(n1241) );
NAND3_X1 U890 ( .A1(n1074), .A2(n1159), .A3(n1242), .ZN(n1228) );
XOR2_X1 U891 ( .A(n1243), .B(n1244), .Z(G39) );
NOR3_X1 U892 ( .A1(n1245), .A2(n1060), .A3(n1234), .ZN(n1244) );
INV_X1 U893 ( .A(n1246), .ZN(n1060) );
XOR2_X1 U894 ( .A(n1236), .B(KEYINPUT23), .Z(n1245) );
NAND2_X1 U895 ( .A1(KEYINPUT27), .A2(n1247), .ZN(n1243) );
INV_X1 U896 ( .A(G137), .ZN(n1247) );
XNOR2_X1 U897 ( .A(G134), .B(n1227), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1046), .A2(n1075), .A3(n1242), .ZN(n1227) );
XNOR2_X1 U899 ( .A(G131), .B(n1226), .ZN(G33) );
NAND3_X1 U900 ( .A1(n1159), .A2(n1075), .A3(n1242), .ZN(n1226) );
INV_X1 U901 ( .A(n1234), .ZN(n1242) );
NAND4_X1 U902 ( .A1(n1248), .A2(n1085), .A3(n1237), .A4(n1064), .ZN(n1234) );
INV_X1 U903 ( .A(n1065), .ZN(n1248) );
INV_X1 U904 ( .A(n1079), .ZN(n1159) );
XOR2_X1 U905 ( .A(G128), .B(n1249), .Z(G30) );
NOR2_X1 U906 ( .A1(n1232), .A2(n1233), .ZN(n1249) );
NAND4_X1 U907 ( .A1(n1046), .A2(n1085), .A3(n1236), .A4(n1237), .ZN(n1233) );
INV_X1 U908 ( .A(n1217), .ZN(n1046) );
XNOR2_X1 U909 ( .A(G101), .B(n1250), .ZN(G3) );
NAND3_X1 U910 ( .A1(n1218), .A2(n1075), .A3(n1251), .ZN(n1250) );
AND2_X1 U911 ( .A1(n1085), .A2(n1061), .ZN(n1218) );
XOR2_X1 U912 ( .A(n1200), .B(n1225), .Z(G27) );
NAND4_X1 U913 ( .A1(n1074), .A2(n1090), .A3(n1061), .A4(n1237), .ZN(n1225) );
NAND2_X1 U914 ( .A1(n1054), .A2(n1252), .ZN(n1237) );
NAND4_X1 U915 ( .A1(n1253), .A2(G953), .A3(G902), .A4(n1115), .ZN(n1252) );
INV_X1 U916 ( .A(G900), .ZN(n1115) );
XOR2_X1 U917 ( .A(n1254), .B(KEYINPUT33), .Z(n1253) );
XOR2_X1 U918 ( .A(n1255), .B(G122), .Z(G24) );
NAND2_X1 U919 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U920 ( .A1(n1137), .A2(n1258), .ZN(n1257) );
INV_X1 U921 ( .A(KEYINPUT3), .ZN(n1258) );
NOR2_X1 U922 ( .A1(n1259), .A2(n1232), .ZN(n1137) );
NAND3_X1 U923 ( .A1(n1061), .A2(n1259), .A3(KEYINPUT3), .ZN(n1256) );
NAND4_X1 U924 ( .A1(n1219), .A2(n1240), .A3(n1099), .A4(n1260), .ZN(n1259) );
NOR2_X1 U925 ( .A1(n1058), .A2(n1059), .ZN(n1260) );
INV_X1 U926 ( .A(n1220), .ZN(n1058) );
XOR2_X1 U927 ( .A(G119), .B(n1261), .Z(G21) );
NOR2_X1 U928 ( .A1(KEYINPUT54), .A2(n1204), .ZN(n1261) );
OR4_X1 U929 ( .A1(n1213), .A2(n1059), .A3(n1232), .A4(n1235), .ZN(n1204) );
INV_X1 U930 ( .A(n1236), .ZN(n1235) );
NAND2_X1 U931 ( .A1(n1262), .A2(n1263), .ZN(n1236) );
NAND3_X1 U932 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
NAND2_X1 U933 ( .A1(KEYINPUT5), .A2(n1074), .ZN(n1262) );
XOR2_X1 U934 ( .A(n1267), .B(n1206), .Z(G18) );
NAND4_X1 U935 ( .A1(n1075), .A2(n1219), .A3(n1061), .A4(n1268), .ZN(n1206) );
NOR2_X1 U936 ( .A1(n1217), .A2(n1059), .ZN(n1268) );
NAND2_X1 U937 ( .A1(n1269), .A2(n1099), .ZN(n1217) );
XOR2_X1 U938 ( .A(n1240), .B(KEYINPUT50), .Z(n1269) );
XNOR2_X1 U939 ( .A(G113), .B(n1205), .ZN(G15) );
NAND4_X1 U940 ( .A1(n1090), .A2(n1061), .A3(n1075), .A4(n1219), .ZN(n1205) );
NAND2_X1 U941 ( .A1(n1270), .A2(n1271), .ZN(n1075) );
NAND3_X1 U942 ( .A1(n1265), .A2(n1272), .A3(n1266), .ZN(n1271) );
INV_X1 U943 ( .A(KEYINPUT5), .ZN(n1266) );
NAND2_X1 U944 ( .A1(KEYINPUT5), .A2(n1220), .ZN(n1270) );
NOR2_X1 U945 ( .A1(n1265), .A2(n1264), .ZN(n1220) );
INV_X1 U946 ( .A(n1272), .ZN(n1264) );
INV_X1 U947 ( .A(n1232), .ZN(n1061) );
NOR2_X1 U948 ( .A1(n1079), .A2(n1059), .ZN(n1090) );
NAND2_X1 U949 ( .A1(n1088), .A2(n1087), .ZN(n1059) );
NAND2_X1 U950 ( .A1(n1273), .A2(n1240), .ZN(n1079) );
INV_X1 U951 ( .A(n1099), .ZN(n1273) );
XOR2_X1 U952 ( .A(G110), .B(n1274), .Z(G12) );
NOR2_X1 U953 ( .A1(n1232), .A2(n1214), .ZN(n1274) );
NAND3_X1 U954 ( .A1(n1074), .A2(n1085), .A3(n1251), .ZN(n1214) );
INV_X1 U955 ( .A(n1213), .ZN(n1251) );
NAND2_X1 U956 ( .A1(n1246), .A2(n1219), .ZN(n1213) );
NAND2_X1 U957 ( .A1(n1054), .A2(n1275), .ZN(n1219) );
NAND4_X1 U958 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1129), .ZN(n1275) );
INV_X1 U959 ( .A(G898), .ZN(n1129) );
NAND3_X1 U960 ( .A1(n1254), .A2(n1113), .A3(G952), .ZN(n1054) );
NAND2_X1 U961 ( .A1(G237), .A2(n1276), .ZN(n1254) );
NOR2_X1 U962 ( .A1(n1099), .A2(n1240), .ZN(n1246) );
NAND3_X1 U963 ( .A1(n1277), .A2(n1278), .A3(n1097), .ZN(n1240) );
NAND2_X1 U964 ( .A1(n1105), .A2(n1106), .ZN(n1097) );
NAND2_X1 U965 ( .A1(n1106), .A2(n1279), .ZN(n1278) );
OR3_X1 U966 ( .A1(n1106), .A2(n1105), .A3(n1279), .ZN(n1277) );
INV_X1 U967 ( .A(KEYINPUT30), .ZN(n1279) );
NOR2_X1 U968 ( .A1(n1156), .A2(G902), .ZN(n1105) );
XNOR2_X1 U969 ( .A(n1280), .B(n1281), .ZN(n1156) );
XNOR2_X1 U970 ( .A(n1282), .B(n1283), .ZN(n1281) );
NAND2_X1 U971 ( .A1(n1284), .A2(KEYINPUT60), .ZN(n1282) );
XOR2_X1 U972 ( .A(n1285), .B(G146), .Z(n1284) );
NAND2_X1 U973 ( .A1(KEYINPUT26), .A2(n1286), .ZN(n1285) );
XOR2_X1 U974 ( .A(n1287), .B(n1288), .Z(n1280) );
XOR2_X1 U975 ( .A(G131), .B(G122), .Z(n1288) );
NAND2_X1 U976 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND2_X1 U977 ( .A1(n1291), .A2(n1238), .ZN(n1290) );
XOR2_X1 U978 ( .A(n1292), .B(KEYINPUT59), .Z(n1289) );
OR2_X1 U979 ( .A1(n1291), .A2(n1238), .ZN(n1292) );
NAND3_X1 U980 ( .A1(n1293), .A2(n1113), .A3(G214), .ZN(n1291) );
INV_X1 U981 ( .A(G475), .ZN(n1106) );
XNOR2_X1 U982 ( .A(n1294), .B(G478), .ZN(n1099) );
NAND2_X1 U983 ( .A1(n1151), .A2(n1295), .ZN(n1294) );
XNOR2_X1 U984 ( .A(n1296), .B(n1297), .ZN(n1151) );
XNOR2_X1 U985 ( .A(n1298), .B(n1299), .ZN(n1297) );
NAND2_X1 U986 ( .A1(G217), .A2(n1300), .ZN(n1298) );
XOR2_X1 U987 ( .A(n1301), .B(n1302), .Z(n1296) );
XOR2_X1 U988 ( .A(G134), .B(G116), .Z(n1302) );
NAND2_X1 U989 ( .A1(n1303), .A2(KEYINPUT38), .ZN(n1301) );
XOR2_X1 U990 ( .A(n1238), .B(n1304), .Z(n1303) );
NOR2_X1 U991 ( .A1(KEYINPUT9), .A2(n1305), .ZN(n1304) );
XOR2_X1 U992 ( .A(KEYINPUT17), .B(G128), .Z(n1305) );
AND2_X1 U993 ( .A1(n1306), .A2(n1087), .ZN(n1085) );
NAND2_X1 U994 ( .A1(G221), .A2(n1307), .ZN(n1087) );
INV_X1 U995 ( .A(n1088), .ZN(n1306) );
XOR2_X1 U996 ( .A(n1186), .B(n1308), .Z(n1088) );
NOR2_X1 U997 ( .A1(KEYINPUT36), .A2(n1107), .ZN(n1308) );
NAND2_X1 U998 ( .A1(n1309), .A2(n1295), .ZN(n1107) );
XOR2_X1 U999 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1000 ( .A(G110), .B(n1312), .Z(n1311) );
XOR2_X1 U1001 ( .A(KEYINPUT51), .B(G140), .Z(n1312) );
XOR2_X1 U1002 ( .A(n1313), .B(n1187), .Z(n1310) );
XNOR2_X1 U1003 ( .A(n1314), .B(n1315), .ZN(n1187) );
XOR2_X1 U1004 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U1005 ( .A(G107), .B(G101), .Z(n1317) );
NOR2_X1 U1006 ( .A1(n1114), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1007 ( .A(KEYINPUT18), .B(G953), .Z(n1318) );
INV_X1 U1008 ( .A(G227), .ZN(n1114) );
XNOR2_X1 U1009 ( .A(n1319), .B(n1170), .ZN(n1314) );
NAND2_X1 U1010 ( .A1(KEYINPUT44), .A2(n1320), .ZN(n1319) );
INV_X1 U1011 ( .A(G104), .ZN(n1320) );
NAND2_X1 U1012 ( .A1(KEYINPUT31), .A2(n1123), .ZN(n1313) );
XOR2_X1 U1013 ( .A(n1238), .B(n1321), .Z(n1123) );
INV_X1 U1014 ( .A(G469), .ZN(n1186) );
NOR2_X1 U1015 ( .A1(n1272), .A2(n1265), .ZN(n1074) );
OR2_X1 U1016 ( .A1(n1322), .A2(n1096), .ZN(n1265) );
NOR2_X1 U1017 ( .A1(n1323), .A2(n1324), .ZN(n1096) );
XOR2_X1 U1018 ( .A(KEYINPUT52), .B(n1098), .Z(n1322) );
NAND2_X1 U1019 ( .A1(n1324), .A2(n1323), .ZN(n1098) );
NAND2_X1 U1020 ( .A1(n1325), .A2(n1295), .ZN(n1323) );
XNOR2_X1 U1021 ( .A(n1173), .B(n1326), .ZN(n1325) );
XOR2_X1 U1022 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1023 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1024 ( .A(n1331), .B(KEYINPUT14), .Z(n1330) );
NAND2_X1 U1025 ( .A1(n1170), .A2(n1171), .ZN(n1331) );
NOR2_X1 U1026 ( .A1(n1170), .A2(n1171), .ZN(n1329) );
XNOR2_X1 U1027 ( .A(n1124), .B(KEYINPUT4), .ZN(n1170) );
XOR2_X1 U1028 ( .A(G131), .B(n1332), .Z(n1124) );
XOR2_X1 U1029 ( .A(G137), .B(G134), .Z(n1332) );
NOR2_X1 U1030 ( .A1(n1333), .A2(n1334), .ZN(n1327) );
XOR2_X1 U1031 ( .A(n1335), .B(KEYINPUT35), .Z(n1334) );
NAND2_X1 U1032 ( .A1(n1336), .A2(n1163), .ZN(n1335) );
NOR2_X1 U1033 ( .A1(n1336), .A2(n1163), .ZN(n1333) );
NAND3_X1 U1034 ( .A1(n1293), .A2(n1113), .A3(n1337), .ZN(n1163) );
XOR2_X1 U1035 ( .A(KEYINPUT37), .B(G210), .Z(n1337) );
XNOR2_X1 U1036 ( .A(KEYINPUT16), .B(G101), .ZN(n1336) );
XOR2_X1 U1037 ( .A(n1338), .B(G113), .Z(n1173) );
NAND2_X1 U1038 ( .A1(KEYINPUT19), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1039 ( .A(G119), .B(G116), .Z(n1339) );
XOR2_X1 U1040 ( .A(G472), .B(KEYINPUT47), .Z(n1324) );
NAND3_X1 U1041 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1272) );
NAND2_X1 U1042 ( .A1(KEYINPUT63), .A2(n1141), .ZN(n1342) );
INV_X1 U1043 ( .A(n1108), .ZN(n1141) );
OR3_X1 U1044 ( .A1(n1343), .A2(KEYINPUT63), .A3(n1109), .ZN(n1341) );
NAND2_X1 U1045 ( .A1(n1109), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1046 ( .A1(KEYINPUT21), .A2(n1108), .ZN(n1343) );
NAND2_X1 U1047 ( .A1(n1144), .A2(n1295), .ZN(n1108) );
NAND3_X1 U1048 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1144) );
OR2_X1 U1049 ( .A1(n1347), .A2(KEYINPUT34), .ZN(n1346) );
NAND3_X1 U1050 ( .A1(KEYINPUT34), .A2(n1347), .A3(n1348), .ZN(n1345) );
INV_X1 U1051 ( .A(n1349), .ZN(n1348) );
NAND2_X1 U1052 ( .A1(n1349), .A2(n1350), .ZN(n1344) );
NAND2_X1 U1053 ( .A1(n1351), .A2(KEYINPUT34), .ZN(n1350) );
XNOR2_X1 U1054 ( .A(n1347), .B(KEYINPUT11), .ZN(n1351) );
XNOR2_X1 U1055 ( .A(n1352), .B(G137), .ZN(n1347) );
NAND2_X1 U1056 ( .A1(G221), .A2(n1300), .ZN(n1352) );
AND2_X1 U1057 ( .A1(G234), .A2(n1113), .ZN(n1300) );
INV_X1 U1058 ( .A(G953), .ZN(n1113) );
XOR2_X1 U1059 ( .A(n1353), .B(n1354), .Z(n1349) );
NOR2_X1 U1060 ( .A1(KEYINPUT55), .A2(n1355), .ZN(n1354) );
XOR2_X1 U1061 ( .A(n1356), .B(G119), .Z(n1355) );
INV_X1 U1062 ( .A(G128), .ZN(n1356) );
XOR2_X1 U1063 ( .A(n1185), .B(n1357), .Z(n1353) );
NOR2_X1 U1064 ( .A1(KEYINPUT7), .A2(n1358), .ZN(n1357) );
NOR2_X1 U1065 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1066 ( .A(n1361), .B(KEYINPUT0), .Z(n1360) );
NAND2_X1 U1067 ( .A1(n1362), .A2(G146), .ZN(n1361) );
XOR2_X1 U1068 ( .A(n1286), .B(KEYINPUT12), .Z(n1362) );
NOR2_X1 U1069 ( .A1(G146), .A2(n1286), .ZN(n1359) );
XNOR2_X1 U1070 ( .A(n1122), .B(KEYINPUT40), .ZN(n1286) );
XOR2_X1 U1071 ( .A(n1200), .B(n1184), .Z(n1122) );
INV_X1 U1072 ( .A(G140), .ZN(n1184) );
INV_X1 U1073 ( .A(G125), .ZN(n1200) );
INV_X1 U1074 ( .A(G110), .ZN(n1185) );
INV_X1 U1075 ( .A(n1145), .ZN(n1109) );
NAND2_X1 U1076 ( .A1(G217), .A2(n1307), .ZN(n1145) );
NAND2_X1 U1077 ( .A1(n1276), .A2(n1295), .ZN(n1307) );
XNOR2_X1 U1078 ( .A(G234), .B(KEYINPUT2), .ZN(n1276) );
NAND2_X1 U1079 ( .A1(n1064), .A2(n1065), .ZN(n1232) );
NAND2_X1 U1080 ( .A1(n1363), .A2(n1364), .ZN(n1065) );
NAND2_X1 U1081 ( .A1(n1104), .A2(n1365), .ZN(n1364) );
XOR2_X1 U1082 ( .A(KEYINPUT46), .B(n1366), .Z(n1363) );
NOR2_X1 U1083 ( .A1(n1104), .A2(n1365), .ZN(n1366) );
XOR2_X1 U1084 ( .A(KEYINPUT32), .B(n1103), .Z(n1365) );
AND2_X1 U1085 ( .A1(G210), .A2(n1367), .ZN(n1103) );
AND2_X1 U1086 ( .A1(n1368), .A2(n1295), .ZN(n1104) );
XOR2_X1 U1087 ( .A(n1138), .B(n1369), .Z(n1368) );
XOR2_X1 U1088 ( .A(G125), .B(n1198), .Z(n1369) );
XOR2_X1 U1089 ( .A(n1171), .B(n1370), .Z(n1198) );
NOR2_X1 U1090 ( .A1(G953), .A2(n1128), .ZN(n1370) );
INV_X1 U1091 ( .A(G224), .ZN(n1128) );
XNOR2_X1 U1092 ( .A(n1371), .B(n1321), .ZN(n1171) );
XOR2_X1 U1093 ( .A(G128), .B(G146), .Z(n1321) );
NAND2_X1 U1094 ( .A1(KEYINPUT62), .A2(n1238), .ZN(n1371) );
INV_X1 U1095 ( .A(G143), .ZN(n1238) );
XOR2_X1 U1096 ( .A(n1372), .B(n1373), .Z(n1138) );
XOR2_X1 U1097 ( .A(n1299), .B(n1283), .Z(n1373) );
XOR2_X1 U1098 ( .A(G104), .B(G113), .Z(n1283) );
XNOR2_X1 U1099 ( .A(n1044), .B(G122), .ZN(n1299) );
INV_X1 U1100 ( .A(G107), .ZN(n1044) );
XOR2_X1 U1101 ( .A(n1374), .B(n1375), .Z(n1372) );
NOR2_X1 U1102 ( .A1(G101), .A2(KEYINPUT29), .ZN(n1375) );
XOR2_X1 U1103 ( .A(n1376), .B(G110), .Z(n1374) );
NAND3_X1 U1104 ( .A1(n1377), .A2(n1378), .A3(n1379), .ZN(n1376) );
OR2_X1 U1105 ( .A1(n1380), .A2(KEYINPUT20), .ZN(n1379) );
NAND3_X1 U1106 ( .A1(KEYINPUT20), .A2(n1380), .A3(G116), .ZN(n1378) );
INV_X1 U1107 ( .A(G119), .ZN(n1380) );
NAND2_X1 U1108 ( .A1(n1381), .A2(n1267), .ZN(n1377) );
INV_X1 U1109 ( .A(G116), .ZN(n1267) );
NAND2_X1 U1110 ( .A1(KEYINPUT20), .A2(n1382), .ZN(n1381) );
XOR2_X1 U1111 ( .A(KEYINPUT45), .B(G119), .Z(n1382) );
NAND2_X1 U1112 ( .A1(G214), .A2(n1367), .ZN(n1064) );
NAND2_X1 U1113 ( .A1(n1293), .A2(n1295), .ZN(n1367) );
INV_X1 U1114 ( .A(G902), .ZN(n1295) );
INV_X1 U1115 ( .A(G237), .ZN(n1293) );
endmodule


