//Key = 1011100011001000101011011010111110011001111111010101110100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317;

XOR2_X1 U733 ( .A(n1005), .B(n1006), .Z(G9) );
NAND2_X1 U734 ( .A1(KEYINPUT8), .A2(G107), .ZN(n1006) );
NOR2_X1 U735 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U736 ( .A1(G953), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1008) );
NOR2_X1 U737 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U738 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U739 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U740 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U741 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U742 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U743 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U744 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1022) );
NOR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U748 ( .A1(n1031), .A2(n1034), .A3(n1025), .ZN(n1018) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR4_X1 U751 ( .A1(n1039), .A2(n1025), .A3(n1021), .A4(n1031), .ZN(n1014) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U753 ( .A1(n1009), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U754 ( .A1(n1042), .A2(n1029), .A3(n1043), .A4(n1044), .ZN(n1009) );
NOR4_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1021), .A4(n1047), .ZN(n1044) );
XOR2_X1 U756 ( .A(KEYINPUT25), .B(n1048), .Z(n1047) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
XNOR2_X1 U758 ( .A(n1051), .B(KEYINPUT46), .ZN(n1050) );
INV_X1 U759 ( .A(n1052), .ZN(n1049) );
XOR2_X1 U760 ( .A(n1053), .B(KEYINPUT12), .Z(n1045) );
NOR3_X1 U761 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1043) );
INV_X1 U762 ( .A(n1057), .ZN(n1056) );
XNOR2_X1 U763 ( .A(n1058), .B(n1059), .ZN(n1042) );
NOR2_X1 U764 ( .A1(KEYINPUT15), .A2(n1060), .ZN(n1058) );
XNOR2_X1 U765 ( .A(G475), .B(KEYINPUT55), .ZN(n1060) );
XOR2_X1 U766 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
AND2_X1 U768 ( .A1(G227), .A2(G900), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1061) );
NAND3_X1 U770 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U771 ( .A1(G953), .A2(n1070), .ZN(n1068) );
XOR2_X1 U772 ( .A(KEYINPUT19), .B(n1071), .Z(n1067) );
OR3_X1 U773 ( .A1(n1071), .A2(G953), .A3(n1069), .ZN(n1065) );
XOR2_X1 U774 ( .A(n1072), .B(n1073), .Z(n1069) );
NAND3_X1 U775 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1072) );
OR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U777 ( .A1(n1078), .A2(n1077), .A3(n1079), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1074) );
NAND2_X1 U779 ( .A1(n1082), .A2(n1077), .ZN(n1081) );
INV_X1 U780 ( .A(KEYINPUT13), .ZN(n1077) );
XNOR2_X1 U781 ( .A(n1078), .B(KEYINPUT44), .ZN(n1082) );
XNOR2_X1 U782 ( .A(n1083), .B(n1084), .ZN(n1078) );
NAND2_X1 U783 ( .A1(KEYINPUT40), .A2(n1085), .ZN(n1083) );
XOR2_X1 U784 ( .A(n1086), .B(n1087), .Z(G69) );
XOR2_X1 U785 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U788 ( .A(KEYINPUT59), .B(n1064), .ZN(n1090) );
NAND2_X1 U789 ( .A1(KEYINPUT26), .A2(n1094), .ZN(n1088) );
NAND2_X1 U790 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U791 ( .A1(G953), .A2(n1097), .ZN(n1096) );
NAND2_X1 U792 ( .A1(G953), .A2(n1098), .ZN(n1086) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1098) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
XNOR2_X1 U797 ( .A(n1105), .B(KEYINPUT3), .ZN(n1099) );
NOR2_X1 U798 ( .A1(n1105), .A2(n1106), .ZN(G63) );
XOR2_X1 U799 ( .A(n1107), .B(n1108), .Z(n1106) );
AND2_X1 U800 ( .A1(G478), .A2(n1109), .ZN(n1107) );
NOR2_X1 U801 ( .A1(n1105), .A2(n1110), .ZN(G60) );
XOR2_X1 U802 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U803 ( .A1(KEYINPUT7), .A2(n1113), .ZN(n1112) );
XNOR2_X1 U804 ( .A(n1114), .B(n1115), .ZN(n1113) );
NAND2_X1 U805 ( .A1(n1109), .A2(G475), .ZN(n1111) );
XNOR2_X1 U806 ( .A(n1116), .B(n1117), .ZN(G6) );
NOR2_X1 U807 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U808 ( .A1(n1105), .A2(n1120), .ZN(G57) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1121) );
XNOR2_X1 U812 ( .A(n1127), .B(n1128), .ZN(n1126) );
AND2_X1 U813 ( .A1(G472), .A2(n1109), .ZN(n1128) );
NAND2_X1 U814 ( .A1(KEYINPUT2), .A2(n1129), .ZN(n1125) );
NOR2_X1 U815 ( .A1(n1105), .A2(n1130), .ZN(G54) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U817 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U818 ( .A(KEYINPUT37), .B(n1135), .Z(n1134) );
NOR2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
AND2_X1 U820 ( .A1(n1137), .A2(n1136), .ZN(n1133) );
AND2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
NAND2_X1 U822 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND3_X1 U824 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1138) );
INV_X1 U825 ( .A(n1141), .ZN(n1144) );
NAND2_X1 U826 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
XNOR2_X1 U827 ( .A(n1147), .B(KEYINPUT28), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1148), .A2(G110), .ZN(n1142) );
INV_X1 U829 ( .A(n1147), .ZN(n1148) );
XOR2_X1 U830 ( .A(n1149), .B(n1079), .Z(n1137) );
XNOR2_X1 U831 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U832 ( .A1(n1152), .A2(KEYINPUT47), .ZN(n1150) );
XNOR2_X1 U833 ( .A(n1153), .B(KEYINPUT9), .ZN(n1152) );
AND2_X1 U834 ( .A1(G469), .A2(n1109), .ZN(n1131) );
NOR2_X1 U835 ( .A1(n1105), .A2(n1154), .ZN(G51) );
XOR2_X1 U836 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U837 ( .A1(KEYINPUT14), .A2(n1157), .ZN(n1156) );
XNOR2_X1 U838 ( .A(n1158), .B(n1159), .ZN(n1157) );
XOR2_X1 U839 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U840 ( .A1(KEYINPUT17), .A2(n1162), .ZN(n1161) );
NAND2_X1 U841 ( .A1(n1109), .A2(n1051), .ZN(n1155) );
INV_X1 U842 ( .A(n1104), .ZN(n1109) );
NAND2_X1 U843 ( .A1(n1163), .A2(n1011), .ZN(n1104) );
NAND3_X1 U844 ( .A1(n1071), .A2(n1092), .A3(n1164), .ZN(n1011) );
XOR2_X1 U845 ( .A(n1093), .B(KEYINPUT10), .Z(n1164) );
AND4_X1 U846 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1092) );
AND4_X1 U847 ( .A1(n1005), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1168) );
INV_X1 U848 ( .A(n1172), .ZN(n1170) );
NAND3_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1040), .ZN(n1005) );
NAND2_X1 U850 ( .A1(n1027), .A2(n1175), .ZN(n1167) );
XNOR2_X1 U851 ( .A(KEYINPUT22), .B(n1119), .ZN(n1175) );
NAND4_X1 U852 ( .A1(n1041), .A2(n1173), .A3(n1036), .A4(n1176), .ZN(n1119) );
INV_X1 U853 ( .A(n1177), .ZN(n1036) );
NAND3_X1 U854 ( .A1(n1178), .A2(n1041), .A3(n1179), .ZN(n1166) );
XNOR2_X1 U855 ( .A(n1033), .B(KEYINPUT29), .ZN(n1179) );
NAND3_X1 U856 ( .A1(n1033), .A2(n1040), .A3(n1178), .ZN(n1165) );
AND2_X1 U857 ( .A1(n1180), .A2(n1181), .ZN(n1071) );
NOR4_X1 U858 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR4_X1 U859 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1180) );
NOR3_X1 U860 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
XNOR2_X1 U861 ( .A(n1193), .B(KEYINPUT33), .ZN(n1191) );
XNOR2_X1 U862 ( .A(G902), .B(KEYINPUT39), .ZN(n1163) );
NOR2_X1 U863 ( .A1(n1064), .A2(G952), .ZN(n1105) );
XNOR2_X1 U864 ( .A(n1194), .B(n1188), .ZN(G48) );
AND3_X1 U865 ( .A1(n1041), .A2(n1027), .A3(n1195), .ZN(n1188) );
NAND2_X1 U866 ( .A1(n1196), .A2(n1197), .ZN(G45) );
NAND2_X1 U867 ( .A1(G143), .A2(n1198), .ZN(n1197) );
XOR2_X1 U868 ( .A(KEYINPUT51), .B(n1199), .Z(n1196) );
NOR2_X1 U869 ( .A1(G143), .A2(n1198), .ZN(n1199) );
INV_X1 U870 ( .A(n1187), .ZN(n1198) );
NOR3_X1 U871 ( .A1(n1190), .A2(n1118), .A3(n1200), .ZN(n1187) );
XOR2_X1 U872 ( .A(G140), .B(n1186), .Z(G42) );
AND3_X1 U873 ( .A1(n1193), .A2(n1032), .A3(n1201), .ZN(n1186) );
NOR3_X1 U874 ( .A1(n1202), .A2(n1203), .A3(n1177), .ZN(n1201) );
XOR2_X1 U875 ( .A(G137), .B(n1185), .Z(G39) );
AND3_X1 U876 ( .A1(n1193), .A2(n1195), .A3(n1204), .ZN(n1185) );
INV_X1 U877 ( .A(n1031), .ZN(n1193) );
XNOR2_X1 U878 ( .A(n1085), .B(n1205), .ZN(G36) );
NOR3_X1 U879 ( .A1(n1190), .A2(n1192), .A3(n1031), .ZN(n1205) );
INV_X1 U880 ( .A(n1040), .ZN(n1192) );
XNOR2_X1 U881 ( .A(G131), .B(n1206), .ZN(G33) );
NOR2_X1 U882 ( .A1(n1184), .A2(KEYINPUT48), .ZN(n1206) );
NOR3_X1 U883 ( .A1(n1031), .A2(n1202), .A3(n1190), .ZN(n1184) );
OR3_X1 U884 ( .A1(n1177), .A2(n1203), .A3(n1207), .ZN(n1190) );
NAND2_X1 U885 ( .A1(n1208), .A2(n1029), .ZN(n1031) );
XNOR2_X1 U886 ( .A(KEYINPUT50), .B(n1028), .ZN(n1208) );
XNOR2_X1 U887 ( .A(n1209), .B(n1183), .ZN(G30) );
AND3_X1 U888 ( .A1(n1040), .A2(n1027), .A3(n1195), .ZN(n1183) );
NOR4_X1 U889 ( .A1(n1177), .A2(n1210), .A3(n1211), .A4(n1203), .ZN(n1195) );
INV_X1 U890 ( .A(n1118), .ZN(n1027) );
XNOR2_X1 U891 ( .A(G101), .B(n1171), .ZN(G3) );
NAND3_X1 U892 ( .A1(n1033), .A2(n1174), .A3(n1204), .ZN(n1171) );
XOR2_X1 U893 ( .A(G125), .B(n1182), .Z(G27) );
AND3_X1 U894 ( .A1(n1032), .A2(n1041), .A3(n1212), .ZN(n1182) );
NOR3_X1 U895 ( .A1(n1021), .A2(n1203), .A3(n1118), .ZN(n1212) );
AND2_X1 U896 ( .A1(n1013), .A2(n1213), .ZN(n1203) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1214), .A4(n1070), .ZN(n1213) );
INV_X1 U898 ( .A(G900), .ZN(n1070) );
INV_X1 U899 ( .A(n1202), .ZN(n1041) );
XNOR2_X1 U900 ( .A(n1215), .B(n1216), .ZN(G24) );
NAND2_X1 U901 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NAND4_X1 U902 ( .A1(n1173), .A2(n1200), .A3(n1178), .A4(n1219), .ZN(n1218) );
INV_X1 U903 ( .A(KEYINPUT18), .ZN(n1219) );
NAND2_X1 U904 ( .A1(n1172), .A2(KEYINPUT18), .ZN(n1217) );
NOR3_X1 U905 ( .A1(n1200), .A2(n1025), .A3(n1220), .ZN(n1172) );
INV_X1 U906 ( .A(n1173), .ZN(n1025) );
NOR2_X1 U907 ( .A1(n1221), .A2(n1046), .ZN(n1173) );
OR2_X1 U908 ( .A1(n1222), .A2(n1053), .ZN(n1200) );
XOR2_X1 U909 ( .A(n1223), .B(n1224), .Z(G21) );
NOR2_X1 U910 ( .A1(KEYINPUT6), .A2(n1093), .ZN(n1224) );
OR4_X1 U911 ( .A1(n1220), .A2(n1017), .A3(n1210), .A4(n1211), .ZN(n1093) );
XNOR2_X1 U912 ( .A(G119), .B(KEYINPUT32), .ZN(n1223) );
XNOR2_X1 U913 ( .A(G116), .B(n1225), .ZN(G18) );
NAND3_X1 U914 ( .A1(n1178), .A2(n1033), .A3(n1226), .ZN(n1225) );
XNOR2_X1 U915 ( .A(n1040), .B(KEYINPUT24), .ZN(n1226) );
NOR2_X1 U916 ( .A1(n1227), .A2(n1053), .ZN(n1040) );
XOR2_X1 U917 ( .A(G113), .B(n1228), .Z(G15) );
NOR4_X1 U918 ( .A1(KEYINPUT11), .A2(n1202), .A3(n1207), .A4(n1220), .ZN(n1228) );
INV_X1 U919 ( .A(n1178), .ZN(n1220) );
NOR3_X1 U920 ( .A1(n1118), .A2(n1229), .A3(n1021), .ZN(n1178) );
NAND2_X1 U921 ( .A1(n1230), .A2(n1038), .ZN(n1021) );
INV_X1 U922 ( .A(n1033), .ZN(n1207) );
NOR2_X1 U923 ( .A1(n1221), .A2(n1211), .ZN(n1033) );
INV_X1 U924 ( .A(n1046), .ZN(n1211) );
NAND2_X1 U925 ( .A1(n1231), .A2(n1227), .ZN(n1202) );
INV_X1 U926 ( .A(n1222), .ZN(n1227) );
XOR2_X1 U927 ( .A(n1169), .B(n1232), .Z(G12) );
NAND2_X1 U928 ( .A1(n1233), .A2(G110), .ZN(n1232) );
XNOR2_X1 U929 ( .A(KEYINPUT63), .B(KEYINPUT52), .ZN(n1233) );
NAND3_X1 U930 ( .A1(n1032), .A2(n1174), .A3(n1204), .ZN(n1169) );
INV_X1 U931 ( .A(n1017), .ZN(n1204) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1222), .ZN(n1017) );
XOR2_X1 U933 ( .A(n1059), .B(G475), .Z(n1222) );
NAND2_X1 U934 ( .A1(n1234), .A2(n1235), .ZN(n1059) );
XNOR2_X1 U935 ( .A(n1115), .B(n1236), .ZN(n1234) );
INV_X1 U936 ( .A(n1114), .ZN(n1236) );
XOR2_X1 U937 ( .A(G104), .B(n1237), .Z(n1114) );
XNOR2_X1 U938 ( .A(n1216), .B(G113), .ZN(n1237) );
XNOR2_X1 U939 ( .A(n1238), .B(n1239), .ZN(n1115) );
NOR2_X1 U940 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U941 ( .A(n1242), .B(KEYINPUT41), .Z(n1241) );
NAND2_X1 U942 ( .A1(G131), .A2(n1243), .ZN(n1242) );
NOR2_X1 U943 ( .A1(G131), .A2(n1243), .ZN(n1240) );
XNOR2_X1 U944 ( .A(n1244), .B(n1245), .ZN(n1243) );
XOR2_X1 U945 ( .A(KEYINPUT62), .B(G143), .Z(n1245) );
NAND2_X1 U946 ( .A1(G214), .A2(n1246), .ZN(n1244) );
NAND2_X1 U947 ( .A1(n1247), .A2(KEYINPUT53), .ZN(n1238) );
XNOR2_X1 U948 ( .A(G146), .B(n1073), .ZN(n1247) );
XOR2_X1 U949 ( .A(n1053), .B(KEYINPUT56), .Z(n1231) );
XOR2_X1 U950 ( .A(n1248), .B(G478), .Z(n1053) );
OR2_X1 U951 ( .A1(n1108), .A2(G902), .ZN(n1248) );
XNOR2_X1 U952 ( .A(n1249), .B(n1250), .ZN(n1108) );
NOR2_X1 U953 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U954 ( .A(KEYINPUT57), .B(n1253), .Z(n1252) );
NOR2_X1 U955 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U956 ( .A(n1256), .B(KEYINPUT42), .Z(n1254) );
NOR2_X1 U957 ( .A1(n1257), .A2(n1256), .ZN(n1251) );
XOR2_X1 U958 ( .A(n1258), .B(n1259), .Z(n1256) );
XNOR2_X1 U959 ( .A(G143), .B(n1209), .ZN(n1259) );
NAND2_X1 U960 ( .A1(KEYINPUT58), .A2(n1085), .ZN(n1258) );
INV_X1 U961 ( .A(G134), .ZN(n1085) );
INV_X1 U962 ( .A(n1255), .ZN(n1257) );
XNOR2_X1 U963 ( .A(n1260), .B(G107), .ZN(n1255) );
NAND2_X1 U964 ( .A1(n1261), .A2(KEYINPUT30), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1262), .B(n1216), .ZN(n1261) );
NAND2_X1 U966 ( .A1(KEYINPUT61), .A2(n1263), .ZN(n1262) );
NAND2_X1 U967 ( .A1(G217), .A2(n1264), .ZN(n1249) );
NOR3_X1 U968 ( .A1(n1177), .A2(n1229), .A3(n1118), .ZN(n1174) );
NAND2_X1 U969 ( .A1(n1028), .A2(n1029), .ZN(n1118) );
NAND2_X1 U970 ( .A1(G214), .A2(n1265), .ZN(n1029) );
OR2_X1 U971 ( .A1(n1054), .A2(n1266), .ZN(n1028) );
AND2_X1 U972 ( .A1(n1051), .A2(n1052), .ZN(n1266) );
NOR2_X1 U973 ( .A1(n1052), .A2(n1051), .ZN(n1054) );
AND2_X1 U974 ( .A1(G210), .A2(n1265), .ZN(n1051) );
NAND2_X1 U975 ( .A1(n1267), .A2(n1235), .ZN(n1265) );
INV_X1 U976 ( .A(G237), .ZN(n1267) );
NAND2_X1 U977 ( .A1(n1268), .A2(n1235), .ZN(n1052) );
XOR2_X1 U978 ( .A(n1160), .B(n1269), .Z(n1268) );
XOR2_X1 U979 ( .A(n1162), .B(n1270), .Z(n1269) );
NAND2_X1 U980 ( .A1(KEYINPUT31), .A2(n1158), .ZN(n1270) );
XOR2_X1 U981 ( .A(G125), .B(n1271), .Z(n1158) );
NAND2_X1 U982 ( .A1(G224), .A2(n1064), .ZN(n1162) );
XNOR2_X1 U983 ( .A(n1095), .B(KEYINPUT4), .ZN(n1160) );
XNOR2_X1 U984 ( .A(n1272), .B(n1273), .ZN(n1095) );
XOR2_X1 U985 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U986 ( .A(G116), .B(n1276), .ZN(n1275) );
NAND2_X1 U987 ( .A1(KEYINPUT20), .A2(n1216), .ZN(n1276) );
INV_X1 U988 ( .A(G122), .ZN(n1216) );
NOR2_X1 U989 ( .A1(G113), .A2(KEYINPUT54), .ZN(n1274) );
XOR2_X1 U990 ( .A(n1277), .B(n1278), .Z(n1272) );
XOR2_X1 U991 ( .A(n1279), .B(n1280), .Z(n1277) );
NAND2_X1 U992 ( .A1(KEYINPUT0), .A2(n1127), .ZN(n1279) );
INV_X1 U993 ( .A(G101), .ZN(n1127) );
INV_X1 U994 ( .A(n1176), .ZN(n1229) );
NAND2_X1 U995 ( .A1(n1013), .A2(n1281), .ZN(n1176) );
NAND4_X1 U996 ( .A1(G953), .A2(G902), .A3(n1214), .A4(n1097), .ZN(n1281) );
INV_X1 U997 ( .A(G898), .ZN(n1097) );
NAND3_X1 U998 ( .A1(n1214), .A2(n1064), .A3(G952), .ZN(n1013) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1214) );
NAND2_X1 U1000 ( .A1(n1037), .A2(n1038), .ZN(n1177) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1282), .ZN(n1038) );
INV_X1 U1002 ( .A(n1230), .ZN(n1037) );
XOR2_X1 U1003 ( .A(n1283), .B(G469), .Z(n1230) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1235), .ZN(n1283) );
XOR2_X1 U1005 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U1006 ( .A(n1287), .B(n1288), .ZN(n1286) );
XNOR2_X1 U1007 ( .A(n1141), .B(n1147), .ZN(n1288) );
XOR2_X1 U1008 ( .A(G140), .B(KEYINPUT5), .Z(n1147) );
NAND2_X1 U1009 ( .A1(G227), .A2(n1064), .ZN(n1141) );
INV_X1 U1010 ( .A(n1153), .ZN(n1287) );
XOR2_X1 U1011 ( .A(n1289), .B(n1290), .Z(n1285) );
XNOR2_X1 U1012 ( .A(G110), .B(n1151), .ZN(n1290) );
NAND2_X1 U1013 ( .A1(n1291), .A2(n1292), .ZN(n1151) );
NAND2_X1 U1014 ( .A1(G101), .A2(n1280), .ZN(n1292) );
XOR2_X1 U1015 ( .A(KEYINPUT23), .B(n1293), .Z(n1291) );
NOR2_X1 U1016 ( .A1(G101), .A2(n1280), .ZN(n1293) );
XNOR2_X1 U1017 ( .A(n1116), .B(G107), .ZN(n1280) );
INV_X1 U1018 ( .A(G104), .ZN(n1116) );
NAND2_X1 U1019 ( .A1(KEYINPUT21), .A2(n1079), .ZN(n1289) );
INV_X1 U1020 ( .A(n1080), .ZN(n1079) );
XOR2_X1 U1021 ( .A(G143), .B(n1294), .Z(n1080) );
NOR2_X1 U1022 ( .A1(n1046), .A2(n1210), .ZN(n1032) );
XOR2_X1 U1023 ( .A(n1221), .B(KEYINPUT35), .Z(n1210) );
NAND2_X1 U1024 ( .A1(n1295), .A2(n1057), .ZN(n1221) );
NAND2_X1 U1025 ( .A1(n1296), .A2(n1103), .ZN(n1057) );
XNOR2_X1 U1026 ( .A(n1055), .B(KEYINPUT38), .ZN(n1295) );
NOR2_X1 U1027 ( .A1(n1103), .A2(n1296), .ZN(n1055) );
NOR2_X1 U1028 ( .A1(n1102), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1029 ( .A(KEYINPUT45), .B(G902), .ZN(n1297) );
XNOR2_X1 U1030 ( .A(n1298), .B(n1299), .ZN(n1102) );
XOR2_X1 U1031 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1032 ( .A(G137), .B(n1302), .Z(n1301) );
NOR2_X1 U1033 ( .A1(KEYINPUT1), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1034 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1035 ( .A(KEYINPUT16), .B(n1194), .ZN(n1305) );
NAND2_X1 U1036 ( .A1(n1306), .A2(KEYINPUT49), .ZN(n1304) );
XNOR2_X1 U1037 ( .A(n1073), .B(KEYINPUT60), .ZN(n1306) );
XOR2_X1 U1038 ( .A(G125), .B(G140), .Z(n1073) );
AND2_X1 U1039 ( .A1(n1264), .A2(G221), .ZN(n1300) );
AND2_X1 U1040 ( .A1(G234), .A2(n1064), .ZN(n1264) );
INV_X1 U1041 ( .A(G953), .ZN(n1064) );
XOR2_X1 U1042 ( .A(n1307), .B(n1278), .Z(n1298) );
XNOR2_X1 U1043 ( .A(G119), .B(n1146), .ZN(n1278) );
INV_X1 U1044 ( .A(G110), .ZN(n1146) );
NAND2_X1 U1045 ( .A1(KEYINPUT36), .A2(n1209), .ZN(n1307) );
INV_X1 U1046 ( .A(G128), .ZN(n1209) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1282), .ZN(n1103) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1235), .ZN(n1282) );
INV_X1 U1049 ( .A(G902), .ZN(n1235) );
XOR2_X1 U1050 ( .A(G472), .B(n1308), .Z(n1046) );
NOR2_X1 U1051 ( .A1(G902), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1052 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1053 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1054 ( .A(n1314), .B(KEYINPUT43), .Z(n1313) );
NAND2_X1 U1055 ( .A1(n1123), .A2(n1124), .ZN(n1314) );
NOR2_X1 U1056 ( .A1(n1123), .A2(n1124), .ZN(n1312) );
XNOR2_X1 U1057 ( .A(n1315), .B(n1316), .ZN(n1124) );
XNOR2_X1 U1058 ( .A(n1263), .B(G113), .ZN(n1316) );
INV_X1 U1059 ( .A(G116), .ZN(n1263) );
XNOR2_X1 U1060 ( .A(G119), .B(KEYINPUT27), .ZN(n1315) );
XNOR2_X1 U1061 ( .A(n1153), .B(n1271), .ZN(n1123) );
XOR2_X1 U1062 ( .A(n1294), .B(n1317), .Z(n1271) );
NOR2_X1 U1063 ( .A1(G143), .A2(KEYINPUT34), .ZN(n1317) );
XNOR2_X1 U1064 ( .A(G128), .B(n1194), .ZN(n1294) );
INV_X1 U1065 ( .A(G146), .ZN(n1194) );
XOR2_X1 U1066 ( .A(G134), .B(n1084), .Z(n1153) );
XOR2_X1 U1067 ( .A(G137), .B(G131), .Z(n1084) );
XNOR2_X1 U1068 ( .A(n1129), .B(G101), .ZN(n1310) );
AND2_X1 U1069 ( .A1(G210), .A2(n1246), .ZN(n1129) );
NOR2_X1 U1070 ( .A1(G237), .A2(G953), .ZN(n1246) );
endmodule


