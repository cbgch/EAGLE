//Key = 0100100010101100011010001011001111010001011000101011111010001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
n1434, n1435, n1436;

XNOR2_X1 U803 ( .A(G107), .B(n1104), .ZN(G9) );
NOR2_X1 U804 ( .A1(n1105), .A2(n1106), .ZN(G75) );
AND3_X1 U805 ( .A1(n1107), .A2(G952), .A3(n1108), .ZN(n1106) );
AND3_X1 U806 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1107) );
NAND2_X1 U807 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U808 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND4_X1 U809 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
NAND2_X1 U810 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U811 ( .A(n1122), .B(KEYINPUT15), .Z(n1120) );
NAND2_X1 U812 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U813 ( .A1(n1125), .A2(n1126), .ZN(n1114) );
NAND2_X1 U814 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U815 ( .A1(n1118), .A2(n1129), .A3(n1117), .ZN(n1128) );
INV_X1 U816 ( .A(n1130), .ZN(n1129) );
NAND2_X1 U817 ( .A1(n1116), .A2(n1131), .ZN(n1127) );
NAND2_X1 U818 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U819 ( .A1(n1118), .A2(n1134), .ZN(n1133) );
NAND2_X1 U820 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U821 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U822 ( .A1(n1117), .A2(n1139), .ZN(n1132) );
OR2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
INV_X1 U824 ( .A(n1142), .ZN(n1125) );
INV_X1 U825 ( .A(n1143), .ZN(n1112) );
NOR3_X1 U826 ( .A1(n1144), .A2(G953), .A3(n1145), .ZN(n1105) );
INV_X1 U827 ( .A(n1109), .ZN(n1145) );
NAND4_X1 U828 ( .A1(n1146), .A2(n1117), .A3(n1147), .A4(n1148), .ZN(n1109) );
NOR4_X1 U829 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1142), .ZN(n1148) );
XOR2_X1 U830 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U831 ( .A1(G472), .A2(KEYINPUT3), .ZN(n1153) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1147) );
XOR2_X1 U833 ( .A(KEYINPUT32), .B(n1156), .Z(n1155) );
NOR2_X1 U834 ( .A1(KEYINPUT22), .A2(G478), .ZN(n1156) );
XNOR2_X1 U835 ( .A(n1157), .B(n1158), .ZN(n1146) );
XNOR2_X1 U836 ( .A(KEYINPUT44), .B(n1159), .ZN(n1158) );
XOR2_X1 U837 ( .A(KEYINPUT14), .B(G952), .Z(n1144) );
XOR2_X1 U838 ( .A(n1160), .B(n1161), .Z(G72) );
NOR2_X1 U839 ( .A1(KEYINPUT19), .A2(n1162), .ZN(n1161) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1110), .ZN(n1162) );
AND2_X1 U841 ( .A1(G227), .A2(G900), .ZN(n1163) );
NOR2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NOR3_X1 U843 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
NOR2_X1 U844 ( .A1(KEYINPUT49), .A2(n1169), .ZN(n1168) );
NOR2_X1 U845 ( .A1(G900), .A2(n1110), .ZN(n1167) );
INV_X1 U846 ( .A(n1170), .ZN(n1166) );
NOR3_X1 U847 ( .A1(n1169), .A2(n1171), .A3(n1172), .ZN(n1164) );
NOR2_X1 U848 ( .A1(G953), .A2(n1173), .ZN(n1172) );
NOR2_X1 U849 ( .A1(KEYINPUT49), .A2(n1170), .ZN(n1173) );
XNOR2_X1 U850 ( .A(n1174), .B(n1175), .ZN(n1170) );
XOR2_X1 U851 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U852 ( .A(n1178), .B(G131), .ZN(n1177) );
NOR2_X1 U853 ( .A1(KEYINPUT29), .A2(n1179), .ZN(n1176) );
XNOR2_X1 U854 ( .A(n1180), .B(n1181), .ZN(n1174) );
NOR2_X1 U855 ( .A1(KEYINPUT49), .A2(n1110), .ZN(n1171) );
INV_X1 U856 ( .A(n1182), .ZN(n1169) );
NAND2_X1 U857 ( .A1(n1183), .A2(n1184), .ZN(G69) );
NAND3_X1 U858 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
OR2_X1 U859 ( .A1(n1110), .A2(G224), .ZN(n1187) );
NAND2_X1 U860 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
XOR2_X1 U861 ( .A(n1190), .B(n1191), .Z(n1188) );
NOR2_X1 U862 ( .A1(G953), .A2(n1192), .ZN(n1191) );
NOR2_X1 U863 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U864 ( .A(n1195), .B(KEYINPUT18), .ZN(n1193) );
NAND4_X1 U865 ( .A1(G953), .A2(n1196), .A3(n1190), .A4(n1189), .ZN(n1183) );
INV_X1 U866 ( .A(KEYINPUT9), .ZN(n1189) );
NAND3_X1 U867 ( .A1(n1197), .A2(n1198), .A3(n1186), .ZN(n1190) );
INV_X1 U868 ( .A(n1199), .ZN(n1186) );
NAND2_X1 U869 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NAND2_X1 U870 ( .A1(n1202), .A2(n1203), .ZN(n1197) );
XNOR2_X1 U871 ( .A(KEYINPUT16), .B(n1201), .ZN(n1202) );
XOR2_X1 U872 ( .A(n1204), .B(n1205), .Z(n1201) );
NAND2_X1 U873 ( .A1(G898), .A2(G224), .ZN(n1196) );
NOR2_X1 U874 ( .A1(n1206), .A2(n1207), .ZN(G66) );
XOR2_X1 U875 ( .A(n1208), .B(n1209), .Z(n1207) );
NAND2_X1 U876 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
NOR2_X1 U877 ( .A1(n1206), .A2(n1212), .ZN(G63) );
XOR2_X1 U878 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND2_X1 U879 ( .A1(n1210), .A2(G478), .ZN(n1213) );
NOR2_X1 U880 ( .A1(n1206), .A2(n1215), .ZN(G60) );
NOR3_X1 U881 ( .A1(n1157), .A2(n1216), .A3(n1217), .ZN(n1215) );
AND3_X1 U882 ( .A1(n1218), .A2(G475), .A3(n1210), .ZN(n1217) );
NOR2_X1 U883 ( .A1(n1219), .A2(n1218), .ZN(n1216) );
NOR2_X1 U884 ( .A1(n1108), .A2(n1159), .ZN(n1219) );
XNOR2_X1 U885 ( .A(G104), .B(n1220), .ZN(G6) );
NOR2_X1 U886 ( .A1(n1221), .A2(KEYINPUT40), .ZN(n1220) );
NOR2_X1 U887 ( .A1(n1206), .A2(n1222), .ZN(G57) );
XOR2_X1 U888 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U889 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U890 ( .A(n1227), .B(n1228), .Z(n1223) );
NOR2_X1 U891 ( .A1(KEYINPUT43), .A2(n1229), .ZN(n1228) );
NAND2_X1 U892 ( .A1(n1210), .A2(G472), .ZN(n1227) );
NOR2_X1 U893 ( .A1(n1206), .A2(n1230), .ZN(G54) );
XOR2_X1 U894 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U895 ( .A(n1233), .B(n1234), .Z(n1232) );
NAND2_X1 U896 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
OR2_X1 U897 ( .A1(n1237), .A2(n1229), .ZN(n1236) );
NAND2_X1 U898 ( .A1(n1238), .A2(n1237), .ZN(n1235) );
NAND2_X1 U899 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
XOR2_X1 U900 ( .A(n1241), .B(KEYINPUT5), .Z(n1239) );
XNOR2_X1 U901 ( .A(n1229), .B(KEYINPUT27), .ZN(n1238) );
NAND2_X1 U902 ( .A1(n1210), .A2(G469), .ZN(n1233) );
XOR2_X1 U903 ( .A(n1242), .B(n1243), .Z(n1231) );
XNOR2_X1 U904 ( .A(G110), .B(n1244), .ZN(n1243) );
NOR2_X1 U905 ( .A1(KEYINPUT38), .A2(G140), .ZN(n1244) );
NOR2_X1 U906 ( .A1(n1206), .A2(n1245), .ZN(G51) );
XOR2_X1 U907 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U908 ( .A(n1248), .B(n1249), .Z(n1247) );
NAND2_X1 U909 ( .A1(n1210), .A2(n1250), .ZN(n1249) );
NOR2_X1 U910 ( .A1(n1251), .A2(n1108), .ZN(n1210) );
NOR3_X1 U911 ( .A1(n1194), .A2(n1195), .A3(n1182), .ZN(n1108) );
NAND4_X1 U912 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1182) );
NOR4_X1 U913 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1255) );
NOR2_X1 U914 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XNOR2_X1 U915 ( .A(KEYINPUT53), .B(n1135), .ZN(n1261) );
AND3_X1 U916 ( .A1(n1140), .A2(n1262), .A3(n1263), .ZN(n1258) );
NOR2_X1 U917 ( .A1(n1264), .A2(n1265), .ZN(n1254) );
NOR2_X1 U918 ( .A1(n1142), .A2(n1266), .ZN(n1265) );
NOR2_X1 U919 ( .A1(n1130), .A2(n1267), .ZN(n1264) );
NOR2_X1 U920 ( .A1(n1268), .A2(n1262), .ZN(n1130) );
OR2_X1 U921 ( .A1(n1269), .A2(KEYINPUT11), .ZN(n1253) );
NAND4_X1 U922 ( .A1(n1268), .A2(n1141), .A3(n1270), .A4(KEYINPUT11), .ZN(n1252) );
NOR3_X1 U923 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND4_X1 U924 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1194) );
AND4_X1 U925 ( .A1(n1278), .A2(n1104), .A3(n1279), .A4(n1280), .ZN(n1277) );
NAND3_X1 U926 ( .A1(n1262), .A2(n1118), .A3(n1281), .ZN(n1104) );
NOR2_X1 U927 ( .A1(n1221), .A2(n1282), .ZN(n1276) );
NOR2_X1 U928 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
AND3_X1 U929 ( .A1(n1281), .A2(n1118), .A3(n1268), .ZN(n1221) );
NAND4_X1 U930 ( .A1(n1140), .A2(n1117), .A3(n1285), .A4(n1121), .ZN(n1275) );
AND3_X1 U931 ( .A1(n1262), .A2(n1284), .A3(n1286), .ZN(n1285) );
INV_X1 U932 ( .A(KEYINPUT24), .ZN(n1284) );
NAND2_X1 U933 ( .A1(n1287), .A2(n1272), .ZN(n1274) );
XOR2_X1 U934 ( .A(n1288), .B(KEYINPUT31), .Z(n1287) );
NAND2_X1 U935 ( .A1(n1289), .A2(KEYINPUT63), .ZN(n1248) );
XNOR2_X1 U936 ( .A(n1290), .B(n1291), .ZN(n1289) );
XOR2_X1 U937 ( .A(G125), .B(n1292), .Z(n1291) );
NOR2_X1 U938 ( .A1(KEYINPUT0), .A2(n1293), .ZN(n1292) );
NOR2_X1 U939 ( .A1(n1110), .A2(G952), .ZN(n1206) );
NAND3_X1 U940 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(G48) );
NAND2_X1 U941 ( .A1(G146), .A2(n1297), .ZN(n1296) );
NAND2_X1 U942 ( .A1(n1298), .A2(n1299), .ZN(n1295) );
INV_X1 U943 ( .A(KEYINPUT39), .ZN(n1299) );
NAND2_X1 U944 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
XNOR2_X1 U945 ( .A(KEYINPUT25), .B(n1297), .ZN(n1300) );
NAND2_X1 U946 ( .A1(KEYINPUT39), .A2(n1302), .ZN(n1294) );
NAND2_X1 U947 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U948 ( .A1(KEYINPUT25), .A2(n1297), .ZN(n1304) );
OR3_X1 U949 ( .A1(G146), .A2(KEYINPUT25), .A3(n1297), .ZN(n1303) );
NAND2_X1 U950 ( .A1(n1305), .A2(n1306), .ZN(n1297) );
XNOR2_X1 U951 ( .A(n1268), .B(KEYINPUT20), .ZN(n1305) );
XNOR2_X1 U952 ( .A(n1307), .B(n1308), .ZN(G45) );
NOR3_X1 U953 ( .A1(n1260), .A2(KEYINPUT59), .A3(n1135), .ZN(n1308) );
NAND3_X1 U954 ( .A1(n1140), .A2(n1272), .A3(n1309), .ZN(n1260) );
NOR3_X1 U955 ( .A1(n1310), .A2(n1273), .A3(n1311), .ZN(n1309) );
XOR2_X1 U956 ( .A(G140), .B(n1257), .Z(G42) );
AND3_X1 U957 ( .A1(n1263), .A2(n1141), .A3(n1268), .ZN(n1257) );
XOR2_X1 U958 ( .A(G137), .B(n1256), .Z(G39) );
AND4_X1 U959 ( .A1(n1263), .A2(n1116), .A3(n1312), .A4(n1313), .ZN(n1256) );
XOR2_X1 U960 ( .A(n1314), .B(n1315), .Z(G36) );
XNOR2_X1 U961 ( .A(G134), .B(KEYINPUT6), .ZN(n1315) );
NAND3_X1 U962 ( .A1(n1263), .A2(n1262), .A3(n1316), .ZN(n1314) );
XNOR2_X1 U963 ( .A(n1140), .B(KEYINPUT54), .ZN(n1316) );
NOR3_X1 U964 ( .A1(n1135), .A2(n1273), .A3(n1142), .ZN(n1263) );
XNOR2_X1 U965 ( .A(n1317), .B(n1318), .ZN(G33) );
NOR2_X1 U966 ( .A1(n1319), .A2(n1142), .ZN(n1318) );
NAND2_X1 U967 ( .A1(n1124), .A2(n1320), .ZN(n1142) );
XOR2_X1 U968 ( .A(n1266), .B(KEYINPUT34), .Z(n1319) );
NAND4_X1 U969 ( .A1(n1140), .A2(n1268), .A3(n1321), .A4(n1322), .ZN(n1266) );
XOR2_X1 U970 ( .A(n1323), .B(n1324), .Z(G30) );
NAND2_X1 U971 ( .A1(KEYINPUT61), .A2(G128), .ZN(n1324) );
NAND2_X1 U972 ( .A1(n1306), .A2(n1262), .ZN(n1323) );
INV_X1 U973 ( .A(n1267), .ZN(n1306) );
NAND3_X1 U974 ( .A1(n1321), .A2(n1312), .A3(n1325), .ZN(n1267) );
XOR2_X1 U975 ( .A(n1278), .B(n1326), .Z(G3) );
XNOR2_X1 U976 ( .A(KEYINPUT42), .B(n1327), .ZN(n1326) );
NAND3_X1 U977 ( .A1(n1116), .A2(n1281), .A3(n1140), .ZN(n1278) );
NAND2_X1 U978 ( .A1(n1328), .A2(n1329), .ZN(G27) );
NAND2_X1 U979 ( .A1(G125), .A2(n1269), .ZN(n1329) );
XOR2_X1 U980 ( .A(KEYINPUT52), .B(n1330), .Z(n1328) );
NOR2_X1 U981 ( .A1(G125), .A2(n1269), .ZN(n1330) );
NAND4_X1 U982 ( .A1(n1325), .A2(n1268), .A3(n1331), .A4(n1117), .ZN(n1269) );
NOR3_X1 U983 ( .A1(n1273), .A2(n1332), .A3(n1121), .ZN(n1325) );
INV_X1 U984 ( .A(n1322), .ZN(n1273) );
NAND2_X1 U985 ( .A1(n1143), .A2(n1333), .ZN(n1322) );
NAND4_X1 U986 ( .A1(G902), .A2(G953), .A3(n1334), .A4(n1335), .ZN(n1333) );
INV_X1 U987 ( .A(G900), .ZN(n1335) );
XNOR2_X1 U988 ( .A(G122), .B(n1280), .ZN(G24) );
NAND4_X1 U989 ( .A1(n1336), .A2(n1118), .A3(n1337), .A4(n1338), .ZN(n1280) );
NOR2_X1 U990 ( .A1(n1313), .A2(n1312), .ZN(n1118) );
XNOR2_X1 U991 ( .A(G119), .B(n1279), .ZN(G21) );
NAND4_X1 U992 ( .A1(n1336), .A2(n1116), .A3(n1312), .A4(n1313), .ZN(n1279) );
XNOR2_X1 U993 ( .A(G116), .B(n1283), .ZN(G18) );
NAND3_X1 U994 ( .A1(n1140), .A2(n1262), .A3(n1336), .ZN(n1283) );
NOR3_X1 U995 ( .A1(n1121), .A2(n1339), .A3(n1271), .ZN(n1336) );
NOR2_X1 U996 ( .A1(n1338), .A2(n1310), .ZN(n1262) );
INV_X1 U997 ( .A(n1337), .ZN(n1310) );
XOR2_X1 U998 ( .A(G113), .B(n1340), .Z(G15) );
NOR2_X1 U999 ( .A1(n1121), .A2(n1288), .ZN(n1340) );
NAND4_X1 U1000 ( .A1(n1140), .A2(n1268), .A3(n1117), .A4(n1286), .ZN(n1288) );
INV_X1 U1001 ( .A(n1271), .ZN(n1117) );
NAND2_X1 U1002 ( .A1(n1138), .A2(n1341), .ZN(n1271) );
NOR2_X1 U1003 ( .A1(n1337), .A2(n1311), .ZN(n1268) );
INV_X1 U1004 ( .A(n1338), .ZN(n1311) );
NOR2_X1 U1005 ( .A1(n1313), .A2(n1331), .ZN(n1140) );
INV_X1 U1006 ( .A(n1312), .ZN(n1331) );
INV_X1 U1007 ( .A(n1332), .ZN(n1313) );
XNOR2_X1 U1008 ( .A(n1342), .B(n1195), .ZN(G12) );
AND3_X1 U1009 ( .A1(n1141), .A2(n1281), .A3(n1116), .ZN(n1195) );
NOR2_X1 U1010 ( .A1(n1337), .A2(n1338), .ZN(n1116) );
XOR2_X1 U1011 ( .A(n1343), .B(n1159), .Z(n1338) );
INV_X1 U1012 ( .A(G475), .ZN(n1159) );
NAND2_X1 U1013 ( .A1(KEYINPUT48), .A2(n1157), .ZN(n1343) );
NOR2_X1 U1014 ( .A1(n1218), .A2(G902), .ZN(n1157) );
XNOR2_X1 U1015 ( .A(n1344), .B(n1345), .ZN(n1218) );
XOR2_X1 U1016 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1017 ( .A(G113), .B(G104), .Z(n1347) );
XNOR2_X1 U1018 ( .A(n1307), .B(G131), .ZN(n1346) );
XOR2_X1 U1019 ( .A(n1348), .B(n1349), .Z(n1344) );
XOR2_X1 U1020 ( .A(n1350), .B(n1351), .Z(n1349) );
NAND2_X1 U1021 ( .A1(n1352), .A2(G214), .ZN(n1351) );
NAND2_X1 U1022 ( .A1(n1353), .A2(n1354), .ZN(n1350) );
NAND2_X1 U1023 ( .A1(n1355), .A2(n1301), .ZN(n1354) );
XOR2_X1 U1024 ( .A(KEYINPUT35), .B(n1356), .Z(n1353) );
NOR2_X1 U1025 ( .A1(n1301), .A2(n1355), .ZN(n1356) );
NAND2_X1 U1026 ( .A1(KEYINPUT4), .A2(n1357), .ZN(n1348) );
XNOR2_X1 U1027 ( .A(n1154), .B(G478), .ZN(n1337) );
NAND2_X1 U1028 ( .A1(n1358), .A2(n1251), .ZN(n1154) );
XNOR2_X1 U1029 ( .A(n1214), .B(KEYINPUT50), .ZN(n1358) );
XNOR2_X1 U1030 ( .A(n1359), .B(n1360), .ZN(n1214) );
XNOR2_X1 U1031 ( .A(n1361), .B(n1362), .ZN(n1360) );
XNOR2_X1 U1032 ( .A(n1178), .B(G122), .ZN(n1362) );
XOR2_X1 U1033 ( .A(n1363), .B(n1364), .Z(n1359) );
AND3_X1 U1034 ( .A1(G217), .A2(n1110), .A3(G234), .ZN(n1364) );
XNOR2_X1 U1035 ( .A(G107), .B(n1365), .ZN(n1363) );
NOR2_X1 U1036 ( .A1(KEYINPUT47), .A2(n1366), .ZN(n1365) );
XNOR2_X1 U1037 ( .A(G128), .B(G143), .ZN(n1366) );
NOR3_X1 U1038 ( .A1(n1121), .A2(n1339), .A3(n1135), .ZN(n1281) );
INV_X1 U1039 ( .A(n1321), .ZN(n1135) );
NOR2_X1 U1040 ( .A1(n1138), .A2(n1137), .ZN(n1321) );
INV_X1 U1041 ( .A(n1341), .ZN(n1137) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1367), .ZN(n1341) );
XOR2_X1 U1043 ( .A(n1368), .B(G469), .Z(n1138) );
NAND2_X1 U1044 ( .A1(n1251), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1045 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1046 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
XNOR2_X1 U1047 ( .A(n1374), .B(n1229), .ZN(n1373) );
XOR2_X1 U1048 ( .A(n1242), .B(n1375), .Z(n1372) );
XOR2_X1 U1049 ( .A(n1376), .B(KEYINPUT7), .Z(n1370) );
NAND2_X1 U1050 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
XNOR2_X1 U1051 ( .A(n1375), .B(n1242), .ZN(n1378) );
NAND2_X1 U1052 ( .A1(G227), .A2(n1110), .ZN(n1242) );
NOR2_X1 U1053 ( .A1(KEYINPUT21), .A2(n1379), .ZN(n1375) );
XNOR2_X1 U1054 ( .A(G140), .B(n1342), .ZN(n1379) );
XNOR2_X1 U1055 ( .A(n1374), .B(n1380), .ZN(n1377) );
INV_X1 U1056 ( .A(n1229), .ZN(n1380) );
NAND2_X1 U1057 ( .A1(n1381), .A2(n1240), .ZN(n1374) );
NAND2_X1 U1058 ( .A1(n1382), .A2(n1180), .ZN(n1240) );
XOR2_X1 U1059 ( .A(n1241), .B(KEYINPUT23), .Z(n1381) );
OR2_X1 U1060 ( .A1(n1180), .A2(n1382), .ZN(n1241) );
XNOR2_X1 U1061 ( .A(n1383), .B(n1384), .ZN(n1382) );
XNOR2_X1 U1062 ( .A(G101), .B(KEYINPUT62), .ZN(n1383) );
XNOR2_X1 U1063 ( .A(n1385), .B(n1386), .ZN(n1180) );
XNOR2_X1 U1064 ( .A(n1387), .B(n1301), .ZN(n1385) );
NAND2_X1 U1065 ( .A1(KEYINPUT60), .A2(n1307), .ZN(n1387) );
INV_X1 U1066 ( .A(n1286), .ZN(n1339) );
NAND2_X1 U1067 ( .A1(n1143), .A2(n1388), .ZN(n1286) );
NAND3_X1 U1068 ( .A1(n1199), .A2(n1334), .A3(G902), .ZN(n1388) );
NOR2_X1 U1069 ( .A1(n1110), .A2(G898), .ZN(n1199) );
NAND3_X1 U1070 ( .A1(n1334), .A2(n1110), .A3(G952), .ZN(n1143) );
NAND2_X1 U1071 ( .A1(G237), .A2(G234), .ZN(n1334) );
INV_X1 U1072 ( .A(n1272), .ZN(n1121) );
NOR2_X1 U1073 ( .A1(n1124), .A2(n1123), .ZN(n1272) );
INV_X1 U1074 ( .A(n1320), .ZN(n1123) );
NAND2_X1 U1075 ( .A1(G214), .A2(n1389), .ZN(n1320) );
XOR2_X1 U1076 ( .A(n1390), .B(n1250), .Z(n1124) );
AND2_X1 U1077 ( .A1(G210), .A2(n1389), .ZN(n1250) );
NAND2_X1 U1078 ( .A1(n1391), .A2(n1251), .ZN(n1389) );
INV_X1 U1079 ( .A(G237), .ZN(n1391) );
NAND2_X1 U1080 ( .A1(n1392), .A2(n1251), .ZN(n1390) );
XOR2_X1 U1081 ( .A(n1393), .B(n1394), .Z(n1392) );
XNOR2_X1 U1082 ( .A(n1246), .B(n1395), .ZN(n1394) );
XNOR2_X1 U1083 ( .A(n1396), .B(n1203), .ZN(n1246) );
INV_X1 U1084 ( .A(n1200), .ZN(n1203) );
XNOR2_X1 U1085 ( .A(G110), .B(n1357), .ZN(n1200) );
INV_X1 U1086 ( .A(G122), .ZN(n1357) );
XOR2_X1 U1087 ( .A(n1397), .B(n1204), .Z(n1396) );
XNOR2_X1 U1088 ( .A(n1398), .B(G113), .ZN(n1204) );
NAND2_X1 U1089 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
NAND2_X1 U1090 ( .A1(G119), .A2(n1361), .ZN(n1400) );
XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n1401), .Z(n1399) );
NOR2_X1 U1092 ( .A1(G119), .A2(n1361), .ZN(n1401) );
INV_X1 U1093 ( .A(G116), .ZN(n1361) );
NAND2_X1 U1094 ( .A1(KEYINPUT12), .A2(n1205), .ZN(n1397) );
XOR2_X1 U1095 ( .A(n1402), .B(G101), .Z(n1205) );
NAND2_X1 U1096 ( .A1(KEYINPUT13), .A2(n1384), .ZN(n1402) );
XNOR2_X1 U1097 ( .A(G104), .B(G107), .ZN(n1384) );
XOR2_X1 U1098 ( .A(n1293), .B(n1403), .Z(n1393) );
NOR2_X1 U1099 ( .A1(KEYINPUT37), .A2(n1404), .ZN(n1403) );
XNOR2_X1 U1100 ( .A(G125), .B(KEYINPUT30), .ZN(n1404) );
NAND2_X1 U1101 ( .A1(G224), .A2(n1110), .ZN(n1293) );
NOR2_X1 U1102 ( .A1(n1312), .A2(n1332), .ZN(n1141) );
NOR2_X1 U1103 ( .A1(n1405), .A2(n1150), .ZN(n1332) );
NOR2_X1 U1104 ( .A1(n1406), .A2(n1211), .ZN(n1150) );
XOR2_X1 U1105 ( .A(n1149), .B(KEYINPUT36), .Z(n1405) );
AND2_X1 U1106 ( .A1(n1211), .A2(n1406), .ZN(n1149) );
NAND2_X1 U1107 ( .A1(n1209), .A2(n1407), .ZN(n1406) );
XNOR2_X1 U1108 ( .A(KEYINPUT56), .B(n1251), .ZN(n1407) );
XOR2_X1 U1109 ( .A(n1408), .B(n1409), .Z(n1209) );
XOR2_X1 U1110 ( .A(n1410), .B(n1411), .Z(n1409) );
XOR2_X1 U1111 ( .A(G119), .B(n1412), .Z(n1411) );
NOR2_X1 U1112 ( .A1(KEYINPUT55), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1113 ( .A(n1414), .B(n1415), .Z(n1413) );
XNOR2_X1 U1114 ( .A(n1301), .B(n1355), .ZN(n1415) );
XOR2_X1 U1115 ( .A(n1181), .B(KEYINPUT41), .Z(n1355) );
XOR2_X1 U1116 ( .A(G125), .B(G140), .Z(n1181) );
XOR2_X1 U1117 ( .A(KEYINPUT58), .B(KEYINPUT2), .Z(n1414) );
AND3_X1 U1118 ( .A1(G221), .A2(n1110), .A3(G234), .ZN(n1410) );
INV_X1 U1119 ( .A(G953), .ZN(n1110) );
XNOR2_X1 U1120 ( .A(n1416), .B(n1417), .ZN(n1408) );
INV_X1 U1121 ( .A(n1179), .ZN(n1417) );
XNOR2_X1 U1122 ( .A(n1418), .B(n1419), .ZN(n1416) );
NAND2_X1 U1123 ( .A1(KEYINPUT8), .A2(G128), .ZN(n1419) );
NAND2_X1 U1124 ( .A1(KEYINPUT26), .A2(n1342), .ZN(n1418) );
AND2_X1 U1125 ( .A1(G217), .A2(n1367), .ZN(n1211) );
NAND2_X1 U1126 ( .A1(G234), .A2(n1251), .ZN(n1367) );
XNOR2_X1 U1127 ( .A(n1152), .B(G472), .ZN(n1312) );
NAND2_X1 U1128 ( .A1(n1420), .A2(n1251), .ZN(n1152) );
INV_X1 U1129 ( .A(G902), .ZN(n1251) );
XNOR2_X1 U1130 ( .A(n1229), .B(n1421), .ZN(n1420) );
XNOR2_X1 U1131 ( .A(n1422), .B(n1225), .ZN(n1421) );
XOR2_X1 U1132 ( .A(n1423), .B(n1395), .Z(n1225) );
INV_X1 U1133 ( .A(n1290), .ZN(n1395) );
XNOR2_X1 U1134 ( .A(n1424), .B(n1386), .ZN(n1290) );
XOR2_X1 U1135 ( .A(G128), .B(KEYINPUT33), .Z(n1386) );
XNOR2_X1 U1136 ( .A(n1425), .B(n1307), .ZN(n1424) );
INV_X1 U1137 ( .A(G143), .ZN(n1307) );
NAND2_X1 U1138 ( .A1(KEYINPUT10), .A2(n1301), .ZN(n1425) );
INV_X1 U1139 ( .A(G146), .ZN(n1301) );
NAND2_X1 U1140 ( .A1(n1426), .A2(n1427), .ZN(n1423) );
NAND2_X1 U1141 ( .A1(n1428), .A2(G113), .ZN(n1427) );
XOR2_X1 U1142 ( .A(KEYINPUT17), .B(n1429), .Z(n1426) );
NOR2_X1 U1143 ( .A1(G113), .A2(n1428), .ZN(n1429) );
XNOR2_X1 U1144 ( .A(G116), .B(n1430), .ZN(n1428) );
NOR2_X1 U1145 ( .A1(G119), .A2(KEYINPUT45), .ZN(n1430) );
NAND2_X1 U1146 ( .A1(KEYINPUT1), .A2(n1226), .ZN(n1422) );
AND2_X1 U1147 ( .A1(n1431), .A2(n1432), .ZN(n1226) );
NAND2_X1 U1148 ( .A1(n1433), .A2(n1327), .ZN(n1432) );
INV_X1 U1149 ( .A(G101), .ZN(n1327) );
NAND2_X1 U1150 ( .A1(n1352), .A2(G210), .ZN(n1433) );
NAND3_X1 U1151 ( .A1(n1352), .A2(G210), .A3(G101), .ZN(n1431) );
NOR2_X1 U1152 ( .A1(G953), .A2(G237), .ZN(n1352) );
XOR2_X1 U1153 ( .A(n1179), .B(n1434), .Z(n1229) );
XNOR2_X1 U1154 ( .A(n1435), .B(n1436), .ZN(n1434) );
NOR2_X1 U1155 ( .A1(KEYINPUT57), .A2(n1317), .ZN(n1436) );
INV_X1 U1156 ( .A(G131), .ZN(n1317) );
NAND2_X1 U1157 ( .A1(KEYINPUT46), .A2(n1178), .ZN(n1435) );
INV_X1 U1158 ( .A(G134), .ZN(n1178) );
XOR2_X1 U1159 ( .A(G137), .B(KEYINPUT28), .Z(n1179) );
INV_X1 U1160 ( .A(G110), .ZN(n1342) );
endmodule


