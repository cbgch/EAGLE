//Key = 1101001010000101101000110110000110111110100011010111010001011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U748 ( .A(G107), .B(n1036), .ZN(G9) );
NOR2_X1 U749 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR4_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR4_X1 U752 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1043) );
NAND3_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1045) );
NAND3_X1 U754 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1051), .A2(n1055), .ZN(n1054) );
NAND2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U757 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
INV_X1 U761 ( .A(n1068), .ZN(n1067) );
NAND3_X1 U762 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1066) );
OR2_X1 U763 ( .A1(n1071), .A2(n1070), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1061) );
NAND3_X1 U765 ( .A1(n1072), .A2(n1074), .A3(n1063), .ZN(n1056) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U767 ( .A1(n1060), .A2(n1077), .ZN(n1076) );
OR2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U769 ( .A1(n1058), .A2(n1080), .ZN(n1075) );
NAND2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U771 ( .A1(n1049), .A2(n1044), .A3(n1050), .ZN(n1082) );
INV_X1 U772 ( .A(KEYINPUT14), .ZN(n1044) );
INV_X1 U773 ( .A(n1083), .ZN(n1051) );
NOR3_X1 U774 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1037) );
INV_X1 U775 ( .A(n1052), .ZN(n1084) );
NAND4_X1 U776 ( .A1(n1085), .A2(n1070), .A3(n1086), .A4(n1087), .ZN(n1052) );
NOR4_X1 U777 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1087) );
XOR2_X1 U778 ( .A(n1092), .B(KEYINPUT40), .Z(n1089) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1088) );
XOR2_X1 U780 ( .A(KEYINPUT62), .B(G472), .Z(n1094) );
NOR2_X1 U781 ( .A1(n1050), .A2(n1069), .ZN(n1086) );
XNOR2_X1 U782 ( .A(n1095), .B(n1096), .ZN(n1085) );
NOR2_X1 U783 ( .A1(n1097), .A2(KEYINPUT12), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(G72) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1053), .ZN(n1099) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U788 ( .A1(n1103), .A2(n1053), .ZN(n1102) );
XOR2_X1 U789 ( .A(n1104), .B(n1042), .Z(n1103) );
NAND3_X1 U790 ( .A1(n1105), .A2(n1104), .A3(G953), .ZN(n1101) );
XNOR2_X1 U791 ( .A(n1106), .B(n1107), .ZN(n1104) );
XNOR2_X1 U792 ( .A(n1108), .B(KEYINPUT63), .ZN(n1107) );
NAND2_X1 U793 ( .A1(KEYINPUT31), .A2(n1109), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1110), .B(n1111), .Z(n1106) );
XOR2_X1 U795 ( .A(KEYINPUT16), .B(n1112), .Z(n1105) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(G69) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1053), .ZN(n1114) );
AND2_X1 U798 ( .A1(G224), .A2(G898), .ZN(n1115) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND3_X1 U800 ( .A1(n1118), .A2(n1119), .A3(n1040), .ZN(n1117) );
NAND2_X1 U801 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U803 ( .A1(G898), .A2(n1123), .ZN(n1121) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1053), .ZN(n1118) );
OR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1124) );
INV_X1 U806 ( .A(KEYINPUT38), .ZN(n1122) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1125), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U809 ( .A1(G898), .A2(n1128), .ZN(n1127) );
NAND2_X1 U810 ( .A1(n1040), .A2(n1129), .ZN(n1128) );
NAND2_X1 U811 ( .A1(KEYINPUT38), .A2(G953), .ZN(n1129) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1053), .ZN(n1126) );
NAND2_X1 U813 ( .A1(KEYINPUT38), .A2(n1040), .ZN(n1130) );
XNOR2_X1 U814 ( .A(n1131), .B(n1132), .ZN(n1123) );
XOR2_X1 U815 ( .A(KEYINPUT22), .B(n1133), .Z(n1132) );
NOR2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1134), .A2(n1140), .ZN(G63) );
XNOR2_X1 U820 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U821 ( .A(n1143), .B(KEYINPUT34), .Z(n1142) );
NAND2_X1 U822 ( .A1(n1138), .A2(G478), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1134), .A2(n1144), .ZN(G60) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U825 ( .A(KEYINPUT19), .B(n1147), .Z(n1146) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
AND2_X1 U827 ( .A1(n1149), .A2(n1148), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1138), .A2(G475), .ZN(n1149) );
XNOR2_X1 U829 ( .A(G104), .B(n1150), .ZN(G6) );
NOR2_X1 U830 ( .A1(n1134), .A2(n1151), .ZN(G57) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U833 ( .A(n1156), .B(KEYINPUT33), .Z(n1152) );
NAND2_X1 U834 ( .A1(n1138), .A2(G472), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1134), .A2(n1157), .ZN(G54) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U837 ( .A(n1160), .B(n1161), .ZN(n1159) );
NAND2_X1 U838 ( .A1(n1138), .A2(G469), .ZN(n1160) );
INV_X1 U839 ( .A(n1162), .ZN(n1138) );
XOR2_X1 U840 ( .A(n1163), .B(n1164), .Z(n1158) );
XOR2_X1 U841 ( .A(n1165), .B(KEYINPUT11), .Z(n1164) );
NAND2_X1 U842 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U843 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U844 ( .A(n1170), .B(KEYINPUT48), .Z(n1166) );
NAND2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1163) );
NAND2_X1 U847 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U848 ( .A1(n1134), .A2(n1177), .ZN(G51) );
XOR2_X1 U849 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U850 ( .A(n1180), .B(n1111), .Z(n1179) );
XOR2_X1 U851 ( .A(G125), .B(n1169), .Z(n1111) );
XNOR2_X1 U852 ( .A(KEYINPUT56), .B(n1181), .ZN(n1178) );
NOR2_X1 U853 ( .A1(n1182), .A2(KEYINPUT42), .ZN(n1181) );
NOR2_X1 U854 ( .A1(n1183), .A2(n1162), .ZN(n1182) );
NAND2_X1 U855 ( .A1(G902), .A2(n1184), .ZN(n1162) );
OR2_X1 U856 ( .A1(n1040), .A2(n1042), .ZN(n1184) );
NAND4_X1 U857 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1042) );
AND4_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1193), .A2(n1060), .ZN(n1187) );
NAND3_X1 U860 ( .A1(n1078), .A2(n1194), .A3(n1195), .ZN(n1186) );
NAND2_X1 U861 ( .A1(n1196), .A2(n1073), .ZN(n1185) );
NAND2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(n1073) );
INV_X1 U863 ( .A(n1199), .ZN(n1196) );
NAND4_X1 U864 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1040) );
AND4_X1 U865 ( .A1(n1204), .A2(n1205), .A3(n1150), .A4(n1036), .ZN(n1203) );
NAND3_X1 U866 ( .A1(n1206), .A2(n1058), .A3(n1207), .ZN(n1036) );
NAND3_X1 U867 ( .A1(n1207), .A2(n1058), .A3(n1208), .ZN(n1150) );
NAND2_X1 U868 ( .A1(n1209), .A2(n1210), .ZN(n1202) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND3_X1 U870 ( .A1(n1213), .A2(n1058), .A3(n1214), .ZN(n1212) );
XNOR2_X1 U871 ( .A(KEYINPUT47), .B(n1215), .ZN(n1211) );
NAND3_X1 U872 ( .A1(n1207), .A2(n1216), .A3(n1063), .ZN(n1200) );
XOR2_X1 U873 ( .A(KEYINPUT27), .B(n1079), .Z(n1216) );
NOR2_X1 U874 ( .A1(n1053), .A2(G952), .ZN(n1134) );
XOR2_X1 U875 ( .A(G146), .B(n1217), .Z(G48) );
NOR2_X1 U876 ( .A1(n1218), .A2(n1199), .ZN(n1217) );
XOR2_X1 U877 ( .A(n1197), .B(KEYINPUT30), .Z(n1218) );
XNOR2_X1 U878 ( .A(G143), .B(n1192), .ZN(G45) );
NAND4_X1 U879 ( .A1(n1219), .A2(n1214), .A3(n1079), .A4(n1209), .ZN(n1192) );
XOR2_X1 U880 ( .A(n1109), .B(n1191), .Z(G42) );
NAND2_X1 U881 ( .A1(n1220), .A2(n1078), .ZN(n1191) );
XOR2_X1 U882 ( .A(n1190), .B(n1221), .Z(G39) );
NAND2_X1 U883 ( .A1(KEYINPUT60), .A2(G137), .ZN(n1221) );
NAND3_X1 U884 ( .A1(n1219), .A2(n1222), .A3(n1060), .ZN(n1190) );
XOR2_X1 U885 ( .A(n1223), .B(n1224), .Z(G36) );
NAND2_X1 U886 ( .A1(n1225), .A2(n1060), .ZN(n1224) );
XNOR2_X1 U887 ( .A(n1193), .B(KEYINPUT25), .ZN(n1225) );
AND3_X1 U888 ( .A1(n1079), .A2(n1206), .A3(n1219), .ZN(n1193) );
XNOR2_X1 U889 ( .A(G131), .B(n1226), .ZN(G33) );
NOR2_X1 U890 ( .A1(n1227), .A2(KEYINPUT20), .ZN(n1226) );
INV_X1 U891 ( .A(n1189), .ZN(n1227) );
NAND2_X1 U892 ( .A1(n1220), .A2(n1079), .ZN(n1189) );
AND3_X1 U893 ( .A1(n1219), .A2(n1208), .A3(n1060), .ZN(n1220) );
NOR2_X1 U894 ( .A1(n1228), .A2(n1050), .ZN(n1060) );
INV_X1 U895 ( .A(n1049), .ZN(n1228) );
INV_X1 U896 ( .A(n1197), .ZN(n1208) );
XOR2_X1 U897 ( .A(G128), .B(n1229), .Z(G30) );
NOR2_X1 U898 ( .A1(n1198), .A2(n1199), .ZN(n1229) );
NAND4_X1 U899 ( .A1(n1230), .A2(n1219), .A3(n1209), .A4(n1090), .ZN(n1199) );
AND2_X1 U900 ( .A1(n1068), .A2(n1194), .ZN(n1219) );
INV_X1 U901 ( .A(n1206), .ZN(n1198) );
XOR2_X1 U902 ( .A(n1231), .B(n1232), .Z(G3) );
NAND3_X1 U903 ( .A1(n1063), .A2(n1207), .A3(n1079), .ZN(n1232) );
NAND3_X1 U904 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(G27) );
OR2_X1 U905 ( .A1(n1236), .A2(G125), .ZN(n1235) );
NAND2_X1 U906 ( .A1(KEYINPUT2), .A2(n1237), .ZN(n1234) );
NAND2_X1 U907 ( .A1(G125), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U908 ( .A(KEYINPUT3), .B(n1236), .ZN(n1238) );
NAND2_X1 U909 ( .A1(n1239), .A2(n1240), .ZN(n1233) );
INV_X1 U910 ( .A(KEYINPUT2), .ZN(n1240) );
NAND2_X1 U911 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
NAND3_X1 U912 ( .A1(KEYINPUT3), .A2(G125), .A3(n1236), .ZN(n1242) );
OR2_X1 U913 ( .A1(n1236), .A2(KEYINPUT3), .ZN(n1241) );
NAND3_X1 U914 ( .A1(n1243), .A2(n1194), .A3(n1195), .ZN(n1236) );
NAND2_X1 U915 ( .A1(n1083), .A2(n1244), .ZN(n1194) );
NAND4_X1 U916 ( .A1(G953), .A2(G902), .A3(n1112), .A4(n1245), .ZN(n1244) );
XOR2_X1 U917 ( .A(G900), .B(KEYINPUT18), .Z(n1112) );
XOR2_X1 U918 ( .A(KEYINPUT4), .B(n1078), .Z(n1243) );
XOR2_X1 U919 ( .A(n1246), .B(n1247), .Z(G24) );
NAND4_X1 U920 ( .A1(n1213), .A2(n1058), .A3(n1248), .A4(n1249), .ZN(n1247) );
XOR2_X1 U921 ( .A(KEYINPUT24), .B(n1214), .Z(n1249) );
AND2_X1 U922 ( .A1(n1250), .A2(n1091), .ZN(n1214) );
XOR2_X1 U923 ( .A(KEYINPUT9), .B(n1209), .Z(n1248) );
INV_X1 U924 ( .A(n1048), .ZN(n1058) );
NAND2_X1 U925 ( .A1(n1251), .A2(n1252), .ZN(n1048) );
XOR2_X1 U926 ( .A(KEYINPUT44), .B(n1090), .Z(n1251) );
XOR2_X1 U927 ( .A(G119), .B(n1253), .Z(G21) );
NOR3_X1 U928 ( .A1(n1215), .A2(KEYINPUT5), .A3(n1081), .ZN(n1253) );
NAND2_X1 U929 ( .A1(n1222), .A2(n1213), .ZN(n1215) );
NOR3_X1 U930 ( .A1(n1046), .A2(n1254), .A3(n1252), .ZN(n1222) );
INV_X1 U931 ( .A(n1063), .ZN(n1046) );
XOR2_X1 U932 ( .A(n1255), .B(n1205), .Z(G18) );
NAND4_X1 U933 ( .A1(n1079), .A2(n1213), .A3(n1206), .A4(n1209), .ZN(n1205) );
NOR2_X1 U934 ( .A1(n1091), .A2(n1256), .ZN(n1206) );
AND2_X1 U935 ( .A1(n1072), .A2(n1257), .ZN(n1213) );
XOR2_X1 U936 ( .A(n1258), .B(n1201), .Z(G15) );
NAND3_X1 U937 ( .A1(n1079), .A2(n1257), .A3(n1195), .ZN(n1201) );
NOR3_X1 U938 ( .A1(n1081), .A2(n1047), .A3(n1197), .ZN(n1195) );
NAND2_X1 U939 ( .A1(n1256), .A2(n1091), .ZN(n1197) );
INV_X1 U940 ( .A(n1072), .ZN(n1047) );
NAND2_X1 U941 ( .A1(n1259), .A2(n1260), .ZN(n1072) );
NAND3_X1 U942 ( .A1(n1070), .A2(n1261), .A3(n1071), .ZN(n1260) );
INV_X1 U943 ( .A(KEYINPUT55), .ZN(n1071) );
NAND2_X1 U944 ( .A1(KEYINPUT55), .A2(n1068), .ZN(n1259) );
INV_X1 U945 ( .A(n1209), .ZN(n1081) );
NOR2_X1 U946 ( .A1(n1252), .A2(n1090), .ZN(n1079) );
INV_X1 U947 ( .A(n1254), .ZN(n1090) );
INV_X1 U948 ( .A(n1230), .ZN(n1252) );
XOR2_X1 U949 ( .A(n1262), .B(n1204), .Z(G12) );
NAND3_X1 U950 ( .A1(n1063), .A2(n1207), .A3(n1078), .ZN(n1204) );
NOR2_X1 U951 ( .A1(n1254), .A2(n1230), .ZN(n1078) );
XOR2_X1 U952 ( .A(n1093), .B(n1263), .Z(n1230) );
NOR2_X1 U953 ( .A1(G472), .A2(KEYINPUT39), .ZN(n1263) );
NAND2_X1 U954 ( .A1(n1264), .A2(n1265), .ZN(n1093) );
XOR2_X1 U955 ( .A(n1154), .B(n1266), .Z(n1264) );
XNOR2_X1 U956 ( .A(n1267), .B(KEYINPUT10), .ZN(n1266) );
NAND2_X1 U957 ( .A1(KEYINPUT32), .A2(n1155), .ZN(n1267) );
XOR2_X1 U958 ( .A(n1268), .B(n1231), .Z(n1155) );
INV_X1 U959 ( .A(G101), .ZN(n1231) );
NAND2_X1 U960 ( .A1(n1269), .A2(G210), .ZN(n1268) );
XNOR2_X1 U961 ( .A(n1270), .B(n1271), .ZN(n1154) );
XOR2_X1 U962 ( .A(n1169), .B(n1272), .Z(n1271) );
XOR2_X1 U963 ( .A(n1273), .B(KEYINPUT45), .Z(n1270) );
XOR2_X1 U964 ( .A(n1274), .B(n1139), .Z(n1254) );
AND2_X1 U965 ( .A1(G217), .A2(n1275), .ZN(n1139) );
NAND2_X1 U966 ( .A1(n1137), .A2(n1265), .ZN(n1274) );
XNOR2_X1 U967 ( .A(n1276), .B(n1277), .ZN(n1137) );
NOR2_X1 U968 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U969 ( .A1(n1280), .A2(G137), .ZN(n1279) );
NOR3_X1 U970 ( .A1(n1281), .A2(G953), .A3(n1282), .ZN(n1280) );
NOR4_X1 U971 ( .A1(G953), .A2(n1283), .A3(n1282), .A4(n1281), .ZN(n1278) );
INV_X1 U972 ( .A(G221), .ZN(n1281) );
INV_X1 U973 ( .A(G234), .ZN(n1282) );
XNOR2_X1 U974 ( .A(G137), .B(KEYINPUT54), .ZN(n1283) );
NAND2_X1 U975 ( .A1(KEYINPUT8), .A2(n1284), .ZN(n1276) );
XOR2_X1 U976 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U977 ( .A(n1287), .B(n1288), .ZN(n1286) );
NAND2_X1 U978 ( .A1(KEYINPUT6), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U979 ( .A(G125), .B(n1290), .ZN(n1289) );
NAND2_X1 U980 ( .A1(KEYINPUT35), .A2(G140), .ZN(n1290) );
XOR2_X1 U981 ( .A(G119), .B(G110), .Z(n1285) );
AND3_X1 U982 ( .A1(n1068), .A2(n1257), .A3(n1209), .ZN(n1207) );
NOR2_X1 U983 ( .A1(n1049), .A2(n1050), .ZN(n1209) );
AND2_X1 U984 ( .A1(G214), .A2(n1291), .ZN(n1050) );
XOR2_X1 U985 ( .A(n1095), .B(n1097), .Z(n1049) );
INV_X1 U986 ( .A(n1183), .ZN(n1097) );
NAND2_X1 U987 ( .A1(G210), .A2(n1291), .ZN(n1183) );
NAND2_X1 U988 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
INV_X1 U989 ( .A(G237), .ZN(n1292) );
NAND2_X1 U990 ( .A1(n1294), .A2(n1265), .ZN(n1095) );
XOR2_X1 U991 ( .A(n1295), .B(n1180), .Z(n1294) );
XNOR2_X1 U992 ( .A(n1296), .B(n1133), .ZN(n1180) );
XOR2_X1 U993 ( .A(G110), .B(G122), .Z(n1133) );
XOR2_X1 U994 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U995 ( .A1(KEYINPUT21), .A2(n1299), .ZN(n1298) );
XOR2_X1 U996 ( .A(KEYINPUT28), .B(n1300), .Z(n1299) );
INV_X1 U997 ( .A(n1131), .ZN(n1300) );
XOR2_X1 U998 ( .A(n1301), .B(n1302), .Z(n1131) );
XNOR2_X1 U999 ( .A(n1272), .B(n1303), .ZN(n1301) );
NOR2_X1 U1000 ( .A1(G104), .A2(KEYINPUT29), .ZN(n1303) );
XNOR2_X1 U1001 ( .A(n1258), .B(n1304), .ZN(n1272) );
XOR2_X1 U1002 ( .A(G119), .B(G116), .Z(n1304) );
NAND2_X1 U1003 ( .A1(G224), .A2(n1053), .ZN(n1297) );
XOR2_X1 U1004 ( .A(n1305), .B(KEYINPUT51), .Z(n1295) );
NAND2_X1 U1005 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1006 ( .A1(G125), .A2(n1171), .ZN(n1307) );
XOR2_X1 U1007 ( .A(n1308), .B(KEYINPUT17), .Z(n1306) );
OR2_X1 U1008 ( .A1(n1171), .A2(G125), .ZN(n1308) );
NAND2_X1 U1009 ( .A1(n1083), .A2(n1309), .ZN(n1257) );
NAND4_X1 U1010 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1310), .ZN(n1309) );
INV_X1 U1011 ( .A(G898), .ZN(n1310) );
NAND3_X1 U1012 ( .A1(n1245), .A2(n1053), .A3(G952), .ZN(n1083) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1245) );
NOR2_X1 U1014 ( .A1(n1070), .A2(n1069), .ZN(n1068) );
INV_X1 U1015 ( .A(n1261), .ZN(n1069) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1275), .ZN(n1261) );
NAND2_X1 U1017 ( .A1(G234), .A2(n1293), .ZN(n1275) );
INV_X1 U1018 ( .A(G902), .ZN(n1293) );
XNOR2_X1 U1019 ( .A(n1311), .B(n1312), .ZN(n1070) );
XOR2_X1 U1020 ( .A(KEYINPUT37), .B(G469), .Z(n1312) );
NAND2_X1 U1021 ( .A1(n1313), .A2(n1265), .ZN(n1311) );
XOR2_X1 U1022 ( .A(n1314), .B(n1315), .Z(n1313) );
NOR2_X1 U1023 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1024 ( .A(n1318), .B(KEYINPUT1), .Z(n1317) );
NAND2_X1 U1025 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1026 ( .A(n1161), .B(KEYINPUT61), .ZN(n1319) );
NOR2_X1 U1027 ( .A1(n1320), .A2(n1161), .ZN(n1316) );
XNOR2_X1 U1028 ( .A(n1273), .B(KEYINPUT50), .ZN(n1161) );
XOR2_X1 U1029 ( .A(n1110), .B(KEYINPUT49), .Z(n1273) );
XNOR2_X1 U1030 ( .A(G131), .B(n1321), .ZN(n1110) );
XOR2_X1 U1031 ( .A(G137), .B(G134), .Z(n1321) );
XOR2_X1 U1032 ( .A(n1322), .B(n1172), .Z(n1320) );
INV_X1 U1033 ( .A(n1168), .ZN(n1172) );
XNOR2_X1 U1034 ( .A(G104), .B(n1302), .ZN(n1168) );
XOR2_X1 U1035 ( .A(G101), .B(n1323), .Z(n1302) );
NAND2_X1 U1036 ( .A1(KEYINPUT57), .A2(n1169), .ZN(n1322) );
INV_X1 U1037 ( .A(n1171), .ZN(n1169) );
XNOR2_X1 U1038 ( .A(G143), .B(n1288), .ZN(n1171) );
XNOR2_X1 U1039 ( .A(G146), .B(n1324), .ZN(n1288) );
NAND4_X1 U1040 ( .A1(KEYINPUT23), .A2(n1173), .A3(n1325), .A4(n1326), .ZN(n1314) );
NAND3_X1 U1041 ( .A1(KEYINPUT13), .A2(n1175), .A3(n1176), .ZN(n1326) );
OR2_X1 U1042 ( .A1(n1176), .A2(KEYINPUT13), .ZN(n1325) );
OR2_X1 U1043 ( .A1(n1176), .A2(n1175), .ZN(n1173) );
XOR2_X1 U1044 ( .A(n1262), .B(n1109), .Z(n1175) );
INV_X1 U1045 ( .A(G140), .ZN(n1109) );
NAND2_X1 U1046 ( .A1(G227), .A2(n1053), .ZN(n1176) );
NOR2_X1 U1047 ( .A1(n1250), .A2(n1091), .ZN(n1063) );
XNOR2_X1 U1048 ( .A(n1327), .B(G475), .ZN(n1091) );
NAND2_X1 U1049 ( .A1(n1148), .A2(n1265), .ZN(n1327) );
XNOR2_X1 U1050 ( .A(n1328), .B(n1329), .ZN(n1148) );
XOR2_X1 U1051 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1052 ( .A(G131), .B(G104), .Z(n1331) );
XOR2_X1 U1053 ( .A(KEYINPUT0), .B(G143), .Z(n1330) );
XOR2_X1 U1054 ( .A(n1332), .B(n1333), .Z(n1328) );
NOR3_X1 U1055 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1333) );
AND2_X1 U1056 ( .A1(n1246), .A2(KEYINPUT58), .ZN(n1336) );
NOR3_X1 U1057 ( .A1(KEYINPUT58), .A2(G113), .A3(n1246), .ZN(n1335) );
NOR2_X1 U1058 ( .A1(n1337), .A2(n1258), .ZN(n1334) );
INV_X1 U1059 ( .A(G113), .ZN(n1258) );
NOR2_X1 U1060 ( .A1(KEYINPUT58), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1061 ( .A(n1246), .B(KEYINPUT52), .Z(n1338) );
INV_X1 U1062 ( .A(G122), .ZN(n1246) );
XOR2_X1 U1063 ( .A(n1339), .B(n1340), .Z(n1332) );
AND2_X1 U1064 ( .A1(G214), .A2(n1269), .ZN(n1340) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1269) );
NAND2_X1 U1066 ( .A1(n1341), .A2(n1342), .ZN(n1339) );
NAND2_X1 U1067 ( .A1(G146), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1068 ( .A(KEYINPUT59), .B(n1344), .Z(n1341) );
NOR2_X1 U1069 ( .A1(G146), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1070 ( .A(KEYINPUT43), .B(n1343), .Z(n1345) );
XOR2_X1 U1071 ( .A(G140), .B(G125), .Z(n1343) );
INV_X1 U1072 ( .A(n1256), .ZN(n1250) );
XOR2_X1 U1073 ( .A(n1092), .B(KEYINPUT7), .Z(n1256) );
XOR2_X1 U1074 ( .A(n1346), .B(G478), .Z(n1092) );
NAND2_X1 U1075 ( .A1(n1141), .A2(n1265), .ZN(n1346) );
XOR2_X1 U1076 ( .A(G902), .B(KEYINPUT36), .Z(n1265) );
XNOR2_X1 U1077 ( .A(n1347), .B(n1348), .ZN(n1141) );
XOR2_X1 U1078 ( .A(n1349), .B(n1323), .Z(n1348) );
XOR2_X1 U1079 ( .A(G107), .B(KEYINPUT26), .Z(n1323) );
AND3_X1 U1080 ( .A1(G217), .A2(n1053), .A3(G234), .ZN(n1349) );
INV_X1 U1081 ( .A(G953), .ZN(n1053) );
XOR2_X1 U1082 ( .A(n1350), .B(n1351), .Z(n1347) );
NOR2_X1 U1083 ( .A1(KEYINPUT46), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1084 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1085 ( .A(n1355), .B(G143), .Z(n1354) );
NAND2_X1 U1086 ( .A1(KEYINPUT15), .A2(n1324), .ZN(n1355) );
XNOR2_X1 U1087 ( .A(G128), .B(KEYINPUT41), .ZN(n1324) );
NAND2_X1 U1088 ( .A1(KEYINPUT53), .A2(n1223), .ZN(n1353) );
INV_X1 U1089 ( .A(G134), .ZN(n1223) );
XOR2_X1 U1090 ( .A(n1255), .B(G122), .Z(n1350) );
INV_X1 U1091 ( .A(G116), .ZN(n1255) );
INV_X1 U1092 ( .A(G110), .ZN(n1262) );
endmodule


