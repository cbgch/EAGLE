//Key = 0101001011111000001101010001001011000011111001011111010101111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427;

XNOR2_X1 U786 ( .A(G107), .B(n1086), .ZN(G9) );
NAND4_X1 U787 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1086) );
NOR2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U789 ( .A(KEYINPUT14), .B(n1093), .Z(n1087) );
NOR2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(G75) );
NOR4_X1 U791 ( .A1(G953), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1095) );
XOR2_X1 U792 ( .A(n1099), .B(KEYINPUT33), .Z(n1097) );
NAND2_X1 U793 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U795 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NAND2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NAND2_X1 U797 ( .A1(n1089), .A2(n1109), .ZN(n1108) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
OR2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U800 ( .A1(n1110), .A2(n1114), .A3(n1089), .ZN(n1102) );
NAND2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND3_X1 U802 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NAND3_X1 U804 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1117) );
INV_X1 U805 ( .A(n1093), .ZN(n1123) );
NAND3_X1 U806 ( .A1(G221), .A2(n1125), .A3(n1126), .ZN(n1122) );
NOR3_X1 U807 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1094) );
AND4_X1 U808 ( .A1(n1106), .A2(n1104), .A3(n1127), .A4(n1128), .ZN(n1096) );
NOR4_X1 U809 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1128) );
XOR2_X1 U810 ( .A(n1133), .B(n1134), .Z(n1131) );
XOR2_X1 U811 ( .A(KEYINPUT25), .B(n1135), .Z(n1134) );
NOR2_X1 U812 ( .A1(KEYINPUT28), .A2(n1136), .ZN(n1135) );
XNOR2_X1 U813 ( .A(n1137), .B(KEYINPUT40), .ZN(n1130) );
XNOR2_X1 U814 ( .A(n1138), .B(n1139), .ZN(n1127) );
NOR2_X1 U815 ( .A1(KEYINPUT36), .A2(n1140), .ZN(n1139) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(G72) );
NOR2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
AND2_X1 U818 ( .A1(G227), .A2(G900), .ZN(n1143) );
NAND2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
NAND3_X1 U820 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
INV_X1 U821 ( .A(n1150), .ZN(n1148) );
OR2_X1 U822 ( .A1(n1147), .A2(n1149), .ZN(n1145) );
NAND2_X1 U823 ( .A1(n1144), .A2(n1151), .ZN(n1149) );
NAND2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1147) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U828 ( .A1(G125), .A2(n1160), .ZN(n1159) );
XOR2_X1 U829 ( .A(KEYINPUT1), .B(n1161), .Z(n1158) );
NOR2_X1 U830 ( .A1(G125), .A2(n1162), .ZN(n1161) );
XOR2_X1 U831 ( .A(KEYINPUT57), .B(G140), .Z(n1162) );
NAND3_X1 U832 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1156) );
INV_X1 U833 ( .A(n1166), .ZN(n1165) );
NAND2_X1 U834 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
INV_X1 U835 ( .A(KEYINPUT51), .ZN(n1168) );
XOR2_X1 U836 ( .A(G131), .B(n1169), .Z(n1167) );
NOR2_X1 U837 ( .A1(G134), .A2(n1170), .ZN(n1169) );
NAND2_X1 U838 ( .A1(KEYINPUT51), .A2(n1171), .ZN(n1163) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(G69) );
NOR2_X1 U840 ( .A1(n1174), .A2(n1144), .ZN(n1173) );
AND2_X1 U841 ( .A1(G224), .A2(G898), .ZN(n1174) );
XOR2_X1 U842 ( .A(n1175), .B(n1176), .Z(n1172) );
NOR2_X1 U843 ( .A1(KEYINPUT31), .A2(n1177), .ZN(n1176) );
NOR3_X1 U844 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NOR2_X1 U845 ( .A1(G898), .A2(n1144), .ZN(n1180) );
AND2_X1 U846 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
XOR2_X1 U847 ( .A(KEYINPUT5), .B(n1183), .Z(n1178) );
NOR2_X1 U848 ( .A1(n1182), .A2(n1181), .ZN(n1183) );
NAND2_X1 U849 ( .A1(n1144), .A2(n1184), .ZN(n1175) );
NAND3_X1 U850 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
XNOR2_X1 U851 ( .A(KEYINPUT59), .B(n1188), .ZN(n1186) );
NOR3_X1 U852 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(G66) );
AND2_X1 U853 ( .A1(KEYINPUT60), .A2(n1192), .ZN(n1191) );
NOR3_X1 U854 ( .A1(KEYINPUT60), .A2(n1144), .A3(n1193), .ZN(n1190) );
INV_X1 U855 ( .A(G952), .ZN(n1193) );
XOR2_X1 U856 ( .A(n1194), .B(n1195), .Z(n1189) );
NOR2_X1 U857 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NOR2_X1 U858 ( .A1(n1192), .A2(n1198), .ZN(G63) );
NOR3_X1 U859 ( .A1(n1138), .A2(n1199), .A3(n1200), .ZN(n1198) );
NOR4_X1 U860 ( .A1(n1201), .A2(n1197), .A3(KEYINPUT24), .A4(n1140), .ZN(n1200) );
NOR2_X1 U861 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
NOR3_X1 U862 ( .A1(n1140), .A2(KEYINPUT24), .A3(n1204), .ZN(n1203) );
INV_X1 U863 ( .A(n1098), .ZN(n1204) );
INV_X1 U864 ( .A(G478), .ZN(n1140) );
NOR2_X1 U865 ( .A1(n1192), .A2(n1205), .ZN(G60) );
XOR2_X1 U866 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U867 ( .A(KEYINPUT39), .B(n1208), .Z(n1207) );
NOR2_X1 U868 ( .A1(n1209), .A2(n1197), .ZN(n1208) );
INV_X1 U869 ( .A(G475), .ZN(n1209) );
XOR2_X1 U870 ( .A(n1210), .B(n1211), .Z(G6) );
NOR2_X1 U871 ( .A1(KEYINPUT34), .A2(n1212), .ZN(n1211) );
INV_X1 U872 ( .A(G104), .ZN(n1212) );
NOR3_X1 U873 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1210) );
NAND3_X1 U874 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1213) );
NAND2_X1 U875 ( .A1(KEYINPUT32), .A2(n1219), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1216) );
INV_X1 U877 ( .A(KEYINPUT32), .ZN(n1221) );
NAND2_X1 U878 ( .A1(n1093), .A2(n1092), .ZN(n1220) );
NOR2_X1 U879 ( .A1(n1192), .A2(n1222), .ZN(G57) );
XOR2_X1 U880 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U882 ( .A(n1227), .B(KEYINPUT30), .Z(n1226) );
NAND2_X1 U883 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
XOR2_X1 U885 ( .A(n1230), .B(KEYINPUT55), .Z(n1229) );
NOR2_X1 U886 ( .A1(n1197), .A2(n1231), .ZN(n1228) );
NAND2_X1 U887 ( .A1(n1232), .A2(n1233), .ZN(n1223) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U889 ( .A(KEYINPUT61), .B(n1236), .Z(n1232) );
NOR2_X1 U890 ( .A1(n1235), .A2(n1234), .ZN(n1236) );
NOR2_X1 U891 ( .A1(n1192), .A2(n1237), .ZN(G54) );
XOR2_X1 U892 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U893 ( .A(n1240), .B(n1154), .ZN(n1239) );
XOR2_X1 U894 ( .A(n1241), .B(n1242), .Z(n1238) );
XNOR2_X1 U895 ( .A(n1243), .B(n1244), .ZN(n1241) );
NOR2_X1 U896 ( .A1(n1245), .A2(n1197), .ZN(n1244) );
INV_X1 U897 ( .A(G469), .ZN(n1245) );
NOR2_X1 U898 ( .A1(n1192), .A2(n1246), .ZN(G51) );
XOR2_X1 U899 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U900 ( .A(n1249), .B(n1250), .Z(n1247) );
NOR2_X1 U901 ( .A1(n1251), .A2(n1197), .ZN(n1250) );
NAND2_X1 U902 ( .A1(G902), .A2(n1098), .ZN(n1197) );
NAND4_X1 U903 ( .A1(n1252), .A2(n1253), .A3(n1187), .A4(n1152), .ZN(n1098) );
AND4_X1 U904 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1152) );
NAND3_X1 U905 ( .A1(n1258), .A2(n1112), .A3(n1259), .ZN(n1254) );
XNOR2_X1 U906 ( .A(n1260), .B(KEYINPUT6), .ZN(n1259) );
AND3_X1 U907 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1187) );
NAND4_X1 U908 ( .A1(n1264), .A2(n1089), .A3(n1109), .A4(n1088), .ZN(n1263) );
NAND2_X1 U909 ( .A1(n1091), .A2(n1265), .ZN(n1109) );
XNOR2_X1 U910 ( .A(n1153), .B(KEYINPUT42), .ZN(n1253) );
AND4_X1 U911 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1153) );
NOR2_X1 U912 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
NOR2_X1 U913 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
INV_X1 U914 ( .A(KEYINPUT8), .ZN(n1272) );
NOR2_X1 U915 ( .A1(KEYINPUT8), .A2(n1274), .ZN(n1270) );
NAND4_X1 U916 ( .A1(n1275), .A2(n1276), .A3(n1264), .A4(n1277), .ZN(n1274) );
XOR2_X1 U917 ( .A(n1278), .B(KEYINPUT19), .Z(n1252) );
NAND2_X1 U918 ( .A1(n1185), .A2(n1188), .ZN(n1278) );
AND3_X1 U919 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1185) );
NAND3_X1 U920 ( .A1(n1260), .A2(n1089), .A3(n1282), .ZN(n1281) );
NAND3_X1 U921 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1279) );
XOR2_X1 U922 ( .A(KEYINPUT11), .B(n1214), .Z(n1284) );
NAND2_X1 U923 ( .A1(n1286), .A2(KEYINPUT27), .ZN(n1249) );
XOR2_X1 U924 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U925 ( .A(KEYINPUT2), .B(G125), .Z(n1288) );
NAND2_X1 U926 ( .A1(KEYINPUT3), .A2(n1289), .ZN(n1287) );
NOR2_X1 U927 ( .A1(n1144), .A2(G952), .ZN(n1192) );
XNOR2_X1 U928 ( .A(G146), .B(n1255), .ZN(G48) );
NAND3_X1 U929 ( .A1(n1276), .A2(n1218), .A3(n1258), .ZN(n1255) );
XNOR2_X1 U930 ( .A(G143), .B(n1290), .ZN(G45) );
NAND4_X1 U931 ( .A1(KEYINPUT53), .A2(n1260), .A3(n1258), .A4(n1112), .ZN(n1290) );
XOR2_X1 U932 ( .A(n1160), .B(n1256), .Z(G42) );
NAND3_X1 U933 ( .A1(n1113), .A2(n1218), .A3(n1291), .ZN(n1256) );
XNOR2_X1 U934 ( .A(n1292), .B(n1257), .ZN(G39) );
NAND2_X1 U935 ( .A1(n1291), .A2(n1283), .ZN(n1257) );
XOR2_X1 U936 ( .A(n1170), .B(KEYINPUT9), .Z(n1292) );
XOR2_X1 U937 ( .A(G134), .B(n1293), .Z(G36) );
NOR2_X1 U938 ( .A1(KEYINPUT26), .A2(n1267), .ZN(n1293) );
NAND3_X1 U939 ( .A1(n1112), .A2(n1277), .A3(n1291), .ZN(n1267) );
XOR2_X1 U940 ( .A(n1294), .B(n1269), .Z(G33) );
NAND3_X1 U941 ( .A1(n1112), .A2(n1218), .A3(n1291), .ZN(n1269) );
AND3_X1 U942 ( .A1(n1093), .A2(n1295), .A3(n1104), .ZN(n1291) );
NOR2_X1 U943 ( .A1(n1296), .A2(n1120), .ZN(n1104) );
INV_X1 U944 ( .A(n1124), .ZN(n1120) );
XNOR2_X1 U945 ( .A(G128), .B(n1273), .ZN(G30) );
NAND3_X1 U946 ( .A1(n1276), .A2(n1277), .A3(n1258), .ZN(n1273) );
NOR2_X1 U947 ( .A1(n1219), .A2(n1275), .ZN(n1258) );
INV_X1 U948 ( .A(n1295), .ZN(n1275) );
XOR2_X1 U949 ( .A(n1235), .B(n1261), .Z(G3) );
NAND2_X1 U950 ( .A1(n1112), .A2(n1297), .ZN(n1261) );
XOR2_X1 U951 ( .A(n1298), .B(n1268), .Z(G27) );
NAND4_X1 U952 ( .A1(n1285), .A2(n1113), .A3(n1218), .A4(n1295), .ZN(n1268) );
NAND2_X1 U953 ( .A1(n1299), .A2(n1300), .ZN(n1295) );
NAND3_X1 U954 ( .A1(G902), .A2(n1301), .A3(n1150), .ZN(n1300) );
NOR2_X1 U955 ( .A1(n1144), .A2(G900), .ZN(n1150) );
XOR2_X1 U956 ( .A(KEYINPUT45), .B(n1100), .Z(n1299) );
INV_X1 U957 ( .A(n1302), .ZN(n1100) );
INV_X1 U958 ( .A(n1115), .ZN(n1285) );
XOR2_X1 U959 ( .A(n1303), .B(G122), .Z(G24) );
NAND2_X1 U960 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND4_X1 U961 ( .A1(n1306), .A2(n1260), .A3(n1282), .A4(n1307), .ZN(n1305) );
INV_X1 U962 ( .A(KEYINPUT54), .ZN(n1307) );
NAND3_X1 U963 ( .A1(n1308), .A2(n1309), .A3(KEYINPUT54), .ZN(n1304) );
NAND4_X1 U964 ( .A1(n1306), .A2(n1260), .A3(n1106), .A4(n1088), .ZN(n1309) );
NOR2_X1 U965 ( .A1(n1310), .A2(n1311), .ZN(n1260) );
XOR2_X1 U966 ( .A(n1215), .B(KEYINPUT41), .Z(n1306) );
INV_X1 U967 ( .A(n1089), .ZN(n1215) );
NOR2_X1 U968 ( .A1(n1312), .A2(n1313), .ZN(n1089) );
XOR2_X1 U969 ( .A(G119), .B(n1314), .Z(G21) );
AND2_X1 U970 ( .A1(n1283), .A2(n1282), .ZN(n1314) );
AND2_X1 U971 ( .A1(n1276), .A2(n1110), .ZN(n1283) );
AND2_X1 U972 ( .A1(n1313), .A2(n1312), .ZN(n1276) );
INV_X1 U973 ( .A(n1315), .ZN(n1312) );
NAND3_X1 U974 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(G18) );
NAND2_X1 U975 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND3_X1 U976 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(n1320) );
NAND2_X1 U977 ( .A1(KEYINPUT13), .A2(n1324), .ZN(n1323) );
OR2_X1 U978 ( .A1(n1325), .A2(KEYINPUT12), .ZN(n1322) );
NAND2_X1 U979 ( .A1(KEYINPUT12), .A2(n1326), .ZN(n1321) );
NAND2_X1 U980 ( .A1(G116), .A2(n1327), .ZN(n1326) );
NAND2_X1 U981 ( .A1(KEYINPUT44), .A2(n1328), .ZN(n1327) );
INV_X1 U982 ( .A(n1280), .ZN(n1319) );
NAND4_X1 U983 ( .A1(n1280), .A2(n1324), .A3(G116), .A4(n1328), .ZN(n1317) );
INV_X1 U984 ( .A(KEYINPUT13), .ZN(n1328) );
INV_X1 U985 ( .A(KEYINPUT44), .ZN(n1324) );
NAND2_X1 U986 ( .A1(KEYINPUT13), .A2(n1329), .ZN(n1316) );
NAND2_X1 U987 ( .A1(G116), .A2(n1330), .ZN(n1329) );
NAND2_X1 U988 ( .A1(KEYINPUT44), .A2(n1280), .ZN(n1330) );
NAND3_X1 U989 ( .A1(n1112), .A2(n1277), .A3(n1282), .ZN(n1280) );
INV_X1 U990 ( .A(n1091), .ZN(n1277) );
NAND2_X1 U991 ( .A1(n1331), .A2(n1311), .ZN(n1091) );
XNOR2_X1 U992 ( .A(n1188), .B(n1332), .ZN(G15) );
NOR2_X1 U993 ( .A1(KEYINPUT52), .A2(n1333), .ZN(n1332) );
NAND3_X1 U994 ( .A1(n1112), .A2(n1218), .A3(n1282), .ZN(n1188) );
NOR2_X1 U995 ( .A1(n1115), .A2(n1214), .ZN(n1282) );
INV_X1 U996 ( .A(n1088), .ZN(n1214) );
NAND2_X1 U997 ( .A1(n1106), .A2(n1308), .ZN(n1115) );
INV_X1 U998 ( .A(n1121), .ZN(n1106) );
NAND2_X1 U999 ( .A1(n1126), .A2(n1334), .ZN(n1121) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1125), .ZN(n1334) );
NOR2_X1 U1001 ( .A1(n1313), .A2(n1315), .ZN(n1112) );
XNOR2_X1 U1002 ( .A(n1262), .B(n1335), .ZN(G12) );
NOR2_X1 U1003 ( .A1(KEYINPUT7), .A2(n1336), .ZN(n1335) );
NAND2_X1 U1004 ( .A1(n1297), .A2(n1113), .ZN(n1262) );
AND2_X1 U1005 ( .A1(n1315), .A2(n1313), .ZN(n1113) );
XNOR2_X1 U1006 ( .A(n1133), .B(n1136), .ZN(n1313) );
INV_X1 U1007 ( .A(n1196), .ZN(n1136) );
NAND2_X1 U1008 ( .A1(G217), .A2(n1125), .ZN(n1196) );
OR2_X1 U1009 ( .A1(n1195), .A2(G902), .ZN(n1133) );
XNOR2_X1 U1010 ( .A(n1337), .B(n1338), .ZN(n1195) );
XOR2_X1 U1011 ( .A(G119), .B(n1339), .Z(n1338) );
XOR2_X1 U1012 ( .A(G137), .B(G128), .Z(n1339) );
XOR2_X1 U1013 ( .A(n1340), .B(n1341), .Z(n1337) );
AND3_X1 U1014 ( .A1(G221), .A2(n1144), .A3(G234), .ZN(n1341) );
XOR2_X1 U1015 ( .A(n1342), .B(G110), .Z(n1340) );
NAND3_X1 U1016 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1342) );
OR2_X1 U1017 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND3_X1 U1018 ( .A1(n1348), .A2(n1346), .A3(n1349), .ZN(n1344) );
INV_X1 U1019 ( .A(KEYINPUT4), .ZN(n1346) );
OR2_X1 U1020 ( .A1(n1349), .A2(n1348), .ZN(n1343) );
AND2_X1 U1021 ( .A1(KEYINPUT10), .A2(n1347), .ZN(n1348) );
XOR2_X1 U1022 ( .A(G146), .B(KEYINPUT47), .Z(n1349) );
NOR2_X1 U1023 ( .A1(n1129), .A2(n1137), .ZN(n1315) );
AND2_X1 U1024 ( .A1(n1350), .A2(n1231), .ZN(n1137) );
NOR2_X1 U1025 ( .A1(n1231), .A2(n1350), .ZN(n1129) );
AND2_X1 U1026 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1027 ( .A(n1230), .B(n1353), .Z(n1351) );
XOR2_X1 U1028 ( .A(n1234), .B(n1354), .Z(n1353) );
NAND2_X1 U1029 ( .A1(KEYINPUT49), .A2(n1235), .ZN(n1354) );
INV_X1 U1030 ( .A(G101), .ZN(n1235) );
NAND3_X1 U1031 ( .A1(n1355), .A2(n1144), .A3(G210), .ZN(n1234) );
XOR2_X1 U1032 ( .A(n1356), .B(n1357), .Z(n1230) );
INV_X1 U1033 ( .A(n1358), .ZN(n1357) );
XOR2_X1 U1034 ( .A(n1289), .B(n1243), .Z(n1356) );
INV_X1 U1035 ( .A(G472), .ZN(n1231) );
AND3_X1 U1036 ( .A1(n1110), .A2(n1088), .A3(n1264), .ZN(n1297) );
INV_X1 U1037 ( .A(n1219), .ZN(n1264) );
NAND2_X1 U1038 ( .A1(n1308), .A2(n1093), .ZN(n1219) );
NOR2_X1 U1039 ( .A1(n1126), .A2(n1359), .ZN(n1093) );
AND2_X1 U1040 ( .A1(G221), .A2(n1125), .ZN(n1359) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1360), .ZN(n1125) );
XOR2_X1 U1042 ( .A(KEYINPUT48), .B(G902), .Z(n1360) );
XOR2_X1 U1043 ( .A(n1361), .B(G469), .Z(n1126) );
NAND2_X1 U1044 ( .A1(n1362), .A2(n1352), .ZN(n1361) );
XOR2_X1 U1045 ( .A(n1363), .B(n1364), .Z(n1362) );
XOR2_X1 U1046 ( .A(n1365), .B(n1366), .Z(n1364) );
NOR2_X1 U1047 ( .A1(KEYINPUT20), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1048 ( .A(n1240), .B(n1368), .Z(n1367) );
XOR2_X1 U1049 ( .A(KEYINPUT29), .B(KEYINPUT15), .Z(n1368) );
XOR2_X1 U1050 ( .A(n1369), .B(n1370), .Z(n1240) );
XOR2_X1 U1051 ( .A(G140), .B(G110), .Z(n1370) );
NAND2_X1 U1052 ( .A1(G227), .A2(n1144), .ZN(n1369) );
NAND3_X1 U1053 ( .A1(n1371), .A2(n1372), .A3(n1373), .ZN(n1365) );
NAND2_X1 U1054 ( .A1(n1154), .A2(n1242), .ZN(n1373) );
NAND2_X1 U1055 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
INV_X1 U1056 ( .A(KEYINPUT58), .ZN(n1375) );
NAND2_X1 U1057 ( .A1(n1376), .A2(n1377), .ZN(n1374) );
XNOR2_X1 U1058 ( .A(KEYINPUT37), .B(n1154), .ZN(n1377) );
NAND2_X1 U1059 ( .A1(KEYINPUT58), .A2(n1378), .ZN(n1371) );
NAND2_X1 U1060 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
NAND2_X1 U1061 ( .A1(KEYINPUT37), .A2(n1154), .ZN(n1380) );
OR3_X1 U1062 ( .A1(n1242), .A2(KEYINPUT37), .A3(n1154), .ZN(n1379) );
XOR2_X1 U1063 ( .A(n1289), .B(KEYINPUT18), .Z(n1154) );
INV_X1 U1064 ( .A(n1376), .ZN(n1242) );
XNOR2_X1 U1065 ( .A(G107), .B(n1381), .ZN(n1376) );
XNOR2_X1 U1066 ( .A(n1243), .B(KEYINPUT62), .ZN(n1363) );
NOR2_X1 U1067 ( .A1(n1171), .A2(n1166), .ZN(n1243) );
NOR3_X1 U1068 ( .A1(n1382), .A2(G137), .A3(n1294), .ZN(n1166) );
NAND2_X1 U1069 ( .A1(n1383), .A2(n1384), .ZN(n1171) );
NAND3_X1 U1070 ( .A1(n1294), .A2(n1382), .A3(n1170), .ZN(n1384) );
INV_X1 U1071 ( .A(G137), .ZN(n1170) );
INV_X1 U1072 ( .A(G134), .ZN(n1382) );
NAND2_X1 U1073 ( .A1(n1385), .A2(G137), .ZN(n1383) );
XOR2_X1 U1074 ( .A(G134), .B(G131), .Z(n1385) );
INV_X1 U1075 ( .A(n1092), .ZN(n1308) );
NAND2_X1 U1076 ( .A1(n1296), .A2(n1124), .ZN(n1092) );
NAND2_X1 U1077 ( .A1(G214), .A2(n1386), .ZN(n1124) );
INV_X1 U1078 ( .A(n1119), .ZN(n1296) );
XNOR2_X1 U1079 ( .A(n1387), .B(n1251), .ZN(n1119) );
NAND2_X1 U1080 ( .A1(G210), .A2(n1386), .ZN(n1251) );
NAND2_X1 U1081 ( .A1(n1355), .A2(n1352), .ZN(n1386) );
NAND2_X1 U1082 ( .A1(n1388), .A2(n1352), .ZN(n1387) );
XNOR2_X1 U1083 ( .A(n1389), .B(n1248), .ZN(n1388) );
XOR2_X1 U1084 ( .A(n1181), .B(n1390), .Z(n1248) );
XOR2_X1 U1085 ( .A(n1391), .B(n1392), .Z(n1390) );
NOR2_X1 U1086 ( .A1(KEYINPUT0), .A2(n1182), .ZN(n1392) );
XNOR2_X1 U1087 ( .A(n1336), .B(G122), .ZN(n1182) );
INV_X1 U1088 ( .A(G110), .ZN(n1336) );
NOR2_X1 U1089 ( .A1(G953), .A2(n1393), .ZN(n1391) );
XOR2_X1 U1090 ( .A(KEYINPUT38), .B(G224), .Z(n1393) );
XNOR2_X1 U1091 ( .A(n1358), .B(n1394), .ZN(n1181) );
XOR2_X1 U1092 ( .A(n1395), .B(n1381), .Z(n1394) );
XOR2_X1 U1093 ( .A(G104), .B(G101), .Z(n1381) );
NOR2_X1 U1094 ( .A1(G107), .A2(KEYINPUT63), .ZN(n1395) );
XOR2_X1 U1095 ( .A(n1333), .B(n1396), .Z(n1358) );
XOR2_X1 U1096 ( .A(G119), .B(G116), .Z(n1396) );
NAND2_X1 U1097 ( .A1(KEYINPUT21), .A2(n1397), .ZN(n1389) );
XOR2_X1 U1098 ( .A(n1298), .B(n1289), .Z(n1397) );
XNOR2_X1 U1099 ( .A(G128), .B(n1398), .ZN(n1289) );
NAND2_X1 U1100 ( .A1(n1302), .A2(n1399), .ZN(n1088) );
NAND4_X1 U1101 ( .A1(G953), .A2(G902), .A3(n1301), .A4(n1400), .ZN(n1399) );
INV_X1 U1102 ( .A(G898), .ZN(n1400) );
NAND3_X1 U1103 ( .A1(n1301), .A2(n1144), .A3(n1401), .ZN(n1302) );
XOR2_X1 U1104 ( .A(KEYINPUT16), .B(G952), .Z(n1401) );
NAND2_X1 U1105 ( .A1(G237), .A2(G234), .ZN(n1301) );
NAND2_X1 U1106 ( .A1(n1402), .A2(n1403), .ZN(n1110) );
OR3_X1 U1107 ( .A1(n1331), .A2(n1132), .A3(KEYINPUT17), .ZN(n1403) );
NAND2_X1 U1108 ( .A1(KEYINPUT17), .A2(n1218), .ZN(n1402) );
INV_X1 U1109 ( .A(n1265), .ZN(n1218) );
NAND2_X1 U1110 ( .A1(n1132), .A2(n1310), .ZN(n1265) );
INV_X1 U1111 ( .A(n1331), .ZN(n1310) );
XNOR2_X1 U1112 ( .A(n1138), .B(n1404), .ZN(n1331) );
XOR2_X1 U1113 ( .A(KEYINPUT23), .B(G478), .Z(n1404) );
NOR2_X1 U1114 ( .A1(n1202), .A2(G902), .ZN(n1138) );
INV_X1 U1115 ( .A(n1201), .ZN(n1202) );
NAND3_X1 U1116 ( .A1(n1405), .A2(n1406), .A3(n1407), .ZN(n1201) );
NAND4_X1 U1117 ( .A1(G234), .A2(G217), .A3(n1408), .A4(n1144), .ZN(n1407) );
NAND2_X1 U1118 ( .A1(KEYINPUT50), .A2(n1409), .ZN(n1408) );
OR2_X1 U1119 ( .A1(n1410), .A2(KEYINPUT35), .ZN(n1409) );
OR2_X1 U1120 ( .A1(n1410), .A2(KEYINPUT50), .ZN(n1406) );
NAND3_X1 U1121 ( .A1(n1410), .A2(n1411), .A3(KEYINPUT50), .ZN(n1405) );
NAND4_X1 U1122 ( .A1(G234), .A2(G217), .A3(n1144), .A4(n1412), .ZN(n1411) );
INV_X1 U1123 ( .A(KEYINPUT35), .ZN(n1412) );
XNOR2_X1 U1124 ( .A(n1413), .B(n1414), .ZN(n1410) );
XNOR2_X1 U1125 ( .A(G107), .B(n1415), .ZN(n1414) );
NAND2_X1 U1126 ( .A1(n1416), .A2(n1417), .ZN(n1415) );
XOR2_X1 U1127 ( .A(G143), .B(G128), .Z(n1417) );
XNOR2_X1 U1128 ( .A(KEYINPUT43), .B(KEYINPUT22), .ZN(n1416) );
XOR2_X1 U1129 ( .A(n1325), .B(n1418), .Z(n1413) );
XOR2_X1 U1130 ( .A(G134), .B(G122), .Z(n1418) );
INV_X1 U1131 ( .A(G116), .ZN(n1325) );
INV_X1 U1132 ( .A(n1311), .ZN(n1132) );
XOR2_X1 U1133 ( .A(n1419), .B(G475), .Z(n1311) );
NAND2_X1 U1134 ( .A1(n1206), .A2(n1352), .ZN(n1419) );
INV_X1 U1135 ( .A(G902), .ZN(n1352) );
XNOR2_X1 U1136 ( .A(n1420), .B(n1421), .ZN(n1206) );
XOR2_X1 U1137 ( .A(G122), .B(G104), .Z(n1421) );
XNOR2_X1 U1138 ( .A(n1422), .B(n1423), .ZN(n1420) );
NOR2_X1 U1139 ( .A1(KEYINPUT46), .A2(n1333), .ZN(n1423) );
INV_X1 U1140 ( .A(G113), .ZN(n1333) );
NOR2_X1 U1141 ( .A1(KEYINPUT56), .A2(n1424), .ZN(n1422) );
XOR2_X1 U1142 ( .A(n1425), .B(n1426), .Z(n1424) );
XOR2_X1 U1143 ( .A(n1398), .B(n1347), .Z(n1426) );
XOR2_X1 U1144 ( .A(n1160), .B(n1298), .Z(n1347) );
INV_X1 U1145 ( .A(G125), .ZN(n1298) );
INV_X1 U1146 ( .A(G140), .ZN(n1160) );
XOR2_X1 U1147 ( .A(G143), .B(G146), .Z(n1398) );
XOR2_X1 U1148 ( .A(n1294), .B(n1427), .Z(n1425) );
AND3_X1 U1149 ( .A1(G214), .A2(n1144), .A3(n1355), .ZN(n1427) );
INV_X1 U1150 ( .A(G237), .ZN(n1355) );
INV_X1 U1151 ( .A(G953), .ZN(n1144) );
INV_X1 U1152 ( .A(G131), .ZN(n1294) );
endmodule


