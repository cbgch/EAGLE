//Key = 1101011101001001001100010001100011000000100011000100001000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;

XNOR2_X1 U735 ( .A(G107), .B(n1020), .ZN(G9) );
NOR2_X1 U736 ( .A1(KEYINPUT51), .A2(n1021), .ZN(n1020) );
NOR4_X1 U737 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
XNOR2_X1 U738 ( .A(KEYINPUT30), .B(n1026), .ZN(n1025) );
NAND2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1023) );
NOR2_X1 U740 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U741 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
NOR2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U745 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U748 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U750 ( .A1(n1050), .A2(n1051), .ZN(n1044) );
NOR2_X1 U751 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
INV_X1 U752 ( .A(n1022), .ZN(n1053) );
NOR3_X1 U753 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1052) );
NOR2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1040) );
NOR2_X1 U755 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1054), .ZN(n1061) );
INV_X1 U758 ( .A(KEYINPUT45), .ZN(n1054) );
NOR3_X1 U759 ( .A1(n1058), .A2(n1064), .A3(n1043), .ZN(n1036) );
NAND2_X1 U760 ( .A1(n1065), .A2(n1028), .ZN(n1058) );
NOR3_X1 U761 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1031) );
NOR4_X1 U763 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U764 ( .A(n1074), .B(G472), .Z(n1073) );
NAND2_X1 U765 ( .A1(KEYINPUT19), .A2(n1075), .ZN(n1074) );
XNOR2_X1 U766 ( .A(n1076), .B(n1077), .ZN(n1072) );
NAND2_X1 U767 ( .A1(KEYINPUT32), .A2(n1078), .ZN(n1076) );
INV_X1 U768 ( .A(n1079), .ZN(n1070) );
NOR3_X1 U769 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1068) );
NOR3_X1 U770 ( .A1(n1083), .A2(KEYINPUT31), .A3(n1084), .ZN(n1082) );
AND2_X1 U771 ( .A1(n1083), .A2(KEYINPUT31), .ZN(n1081) );
XOR2_X1 U772 ( .A(G478), .B(n1085), .Z(n1080) );
XOR2_X1 U773 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U774 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U776 ( .A1(n1092), .A2(G953), .ZN(n1091) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1090) );
XOR2_X1 U778 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U779 ( .A1(G125), .A2(KEYINPUT37), .ZN(n1096) );
XOR2_X1 U780 ( .A(n1097), .B(n1098), .Z(n1093) );
XOR2_X1 U781 ( .A(KEYINPUT25), .B(G143), .Z(n1098) );
NAND2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U784 ( .A1(n1103), .A2(n1099), .ZN(n1086) );
AND2_X1 U785 ( .A1(G227), .A2(G900), .ZN(n1103) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U788 ( .A1(G953), .A2(n1108), .ZN(n1107) );
NAND2_X1 U789 ( .A1(G898), .A2(G224), .ZN(n1108) );
INV_X1 U790 ( .A(n1109), .ZN(n1106) );
NAND2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U793 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(n1109) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U796 ( .A(n1099), .B(KEYINPUT40), .Z(n1117) );
NAND2_X1 U797 ( .A1(n1118), .A2(n1111), .ZN(n1114) );
INV_X1 U798 ( .A(n1119), .ZN(n1111) );
XOR2_X1 U799 ( .A(n1120), .B(n1121), .Z(n1118) );
NOR2_X1 U800 ( .A1(KEYINPUT11), .A2(n1122), .ZN(n1120) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U804 ( .A1(n1083), .A2(n1129), .ZN(n1128) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1130), .ZN(G63) );
NOR3_X1 U806 ( .A1(n1085), .A2(n1131), .A3(n1132), .ZN(n1130) );
AND3_X1 U807 ( .A1(n1133), .A2(G478), .A3(n1134), .ZN(n1132) );
NOR2_X1 U808 ( .A1(n1135), .A2(n1133), .ZN(n1131) );
AND2_X1 U809 ( .A1(n1033), .A2(G478), .ZN(n1135) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1136), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR3_X1 U812 ( .A1(n1129), .A2(KEYINPUT35), .A3(n1139), .ZN(n1138) );
INV_X1 U813 ( .A(G475), .ZN(n1139) );
XOR2_X1 U814 ( .A(n1140), .B(n1141), .Z(G6) );
NAND2_X1 U815 ( .A1(KEYINPUT0), .A2(n1142), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1125), .A2(n1143), .ZN(G57) );
XOR2_X1 U817 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U818 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U819 ( .A1(KEYINPUT26), .A2(n1148), .ZN(n1147) );
AND2_X1 U820 ( .A1(G472), .A2(n1134), .ZN(n1146) );
NOR2_X1 U821 ( .A1(n1125), .A2(n1149), .ZN(G54) );
XOR2_X1 U822 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U823 ( .A1(KEYINPUT42), .A2(n1152), .ZN(n1151) );
NOR3_X1 U824 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NOR2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
INV_X1 U826 ( .A(n1158), .ZN(n1157) );
NOR2_X1 U827 ( .A1(KEYINPUT60), .A2(n1159), .ZN(n1156) );
XNOR2_X1 U828 ( .A(n1160), .B(KEYINPUT12), .ZN(n1159) );
NOR3_X1 U829 ( .A1(n1158), .A2(KEYINPUT60), .A3(n1160), .ZN(n1154) );
XNOR2_X1 U830 ( .A(n1161), .B(n1162), .ZN(n1158) );
NOR3_X1 U831 ( .A1(n1163), .A2(KEYINPUT14), .A3(n1164), .ZN(n1162) );
NOR2_X1 U832 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U833 ( .A(n1167), .B(KEYINPUT44), .Z(n1166) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
NOR2_X1 U835 ( .A1(G140), .A2(n1170), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1171), .A2(n1097), .ZN(n1163) );
NOR2_X1 U837 ( .A1(n1170), .A2(n1169), .ZN(n1171) );
XOR2_X1 U838 ( .A(KEYINPUT2), .B(G110), .Z(n1169) );
INV_X1 U839 ( .A(KEYINPUT23), .ZN(n1170) );
AND2_X1 U840 ( .A1(n1160), .A2(KEYINPUT60), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1134), .A2(G469), .ZN(n1150) );
INV_X1 U842 ( .A(n1129), .ZN(n1134) );
NOR2_X1 U843 ( .A1(n1125), .A2(n1172), .ZN(G51) );
XOR2_X1 U844 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U846 ( .A1(n1177), .A2(n1129), .ZN(n1176) );
NAND2_X1 U847 ( .A1(G902), .A2(n1033), .ZN(n1129) );
NAND3_X1 U848 ( .A1(n1101), .A2(n1178), .A3(n1116), .ZN(n1033) );
AND4_X1 U849 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1116) );
NOR4_X1 U850 ( .A1(n1183), .A2(n1141), .A3(n1184), .A4(n1185), .ZN(n1182) );
NOR4_X1 U851 ( .A1(n1186), .A2(n1051), .A3(n1187), .A4(n1188), .ZN(n1185) );
XOR2_X1 U852 ( .A(n1022), .B(KEYINPUT59), .Z(n1186) );
NOR4_X1 U853 ( .A1(n1022), .A2(n1189), .A3(n1190), .A4(n1039), .ZN(n1184) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1026), .ZN(n1189) );
XOR2_X1 U855 ( .A(KEYINPUT52), .B(n1060), .Z(n1191) );
NOR4_X1 U856 ( .A1(n1192), .A2(n1188), .A3(n1022), .A4(n1051), .ZN(n1141) );
INV_X1 U857 ( .A(n1028), .ZN(n1051) );
INV_X1 U858 ( .A(n1193), .ZN(n1183) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1195), .ZN(n1181) );
NOR4_X1 U860 ( .A1(n1188), .A2(n1192), .A3(n1190), .A4(n1196), .ZN(n1194) );
XOR2_X1 U861 ( .A(KEYINPUT6), .B(n1065), .Z(n1196) );
XNOR2_X1 U862 ( .A(KEYINPUT15), .B(n1102), .ZN(n1178) );
AND4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1101) );
NOR3_X1 U864 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
INV_X1 U865 ( .A(n1204), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1064), .A2(n1205), .ZN(n1201) );
NOR2_X1 U867 ( .A1(n1206), .A2(n1027), .ZN(n1064) );
NOR2_X1 U868 ( .A1(KEYINPUT24), .A2(n1207), .ZN(n1175) );
XOR2_X1 U869 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U870 ( .A1(KEYINPUT55), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U871 ( .A(G125), .B(n1211), .ZN(n1208) );
NOR2_X1 U872 ( .A1(n1099), .A2(G952), .ZN(n1125) );
NAND2_X1 U873 ( .A1(n1212), .A2(n1213), .ZN(G48) );
OR4_X1 U874 ( .A1(n1214), .A2(n1205), .A3(n1215), .A4(KEYINPUT21), .ZN(n1213) );
NAND3_X1 U875 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1212) );
OR2_X1 U876 ( .A1(n1205), .A2(n1215), .ZN(n1218) );
XOR2_X1 U877 ( .A(n1192), .B(KEYINPUT39), .Z(n1215) );
OR3_X1 U878 ( .A1(n1214), .A2(KEYINPUT21), .A3(KEYINPUT8), .ZN(n1217) );
NAND2_X1 U879 ( .A1(n1214), .A2(KEYINPUT8), .ZN(n1216) );
XOR2_X1 U880 ( .A(G146), .B(KEYINPUT56), .Z(n1214) );
XOR2_X1 U881 ( .A(n1219), .B(n1204), .Z(G45) );
NAND3_X1 U882 ( .A1(n1220), .A2(n1049), .A3(n1221), .ZN(n1204) );
XOR2_X1 U883 ( .A(G140), .B(n1202), .Z(G42) );
AND3_X1 U884 ( .A1(n1048), .A2(n1206), .A3(n1222), .ZN(n1202) );
XOR2_X1 U885 ( .A(n1199), .B(n1223), .Z(G39) );
XOR2_X1 U886 ( .A(KEYINPUT49), .B(G137), .Z(n1223) );
NAND4_X1 U887 ( .A1(n1222), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1199) );
XNOR2_X1 U888 ( .A(G134), .B(n1197), .ZN(G36) );
NAND3_X1 U889 ( .A1(n1049), .A2(n1027), .A3(n1222), .ZN(n1197) );
INV_X1 U890 ( .A(n1187), .ZN(n1027) );
XNOR2_X1 U891 ( .A(G131), .B(n1102), .ZN(G33) );
NAND3_X1 U892 ( .A1(n1049), .A2(n1206), .A3(n1222), .ZN(n1102) );
NOR3_X1 U893 ( .A1(n1022), .A2(n1227), .A3(n1043), .ZN(n1222) );
INV_X1 U894 ( .A(n1067), .ZN(n1043) );
NOR2_X1 U895 ( .A1(n1062), .A2(n1063), .ZN(n1067) );
INV_X1 U896 ( .A(n1228), .ZN(n1063) );
XOR2_X1 U897 ( .A(G128), .B(n1229), .Z(G30) );
NOR2_X1 U898 ( .A1(n1187), .A2(n1205), .ZN(n1229) );
NAND3_X1 U899 ( .A1(n1225), .A2(n1226), .A3(n1221), .ZN(n1205) );
NOR3_X1 U900 ( .A1(n1022), .A2(n1227), .A3(n1024), .ZN(n1221) );
XOR2_X1 U901 ( .A(G101), .B(n1230), .Z(G3) );
AND2_X1 U902 ( .A1(n1049), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U903 ( .A(G125), .B(n1198), .ZN(G27) );
NAND4_X1 U904 ( .A1(n1048), .A2(n1206), .A3(n1232), .A4(n1065), .ZN(n1198) );
NOR2_X1 U905 ( .A1(n1227), .A2(n1024), .ZN(n1232) );
AND2_X1 U906 ( .A1(n1035), .A2(n1233), .ZN(n1227) );
NAND4_X1 U907 ( .A1(n1092), .A2(G902), .A3(G953), .A4(n1234), .ZN(n1233) );
XNOR2_X1 U908 ( .A(G900), .B(KEYINPUT36), .ZN(n1092) );
XOR2_X1 U909 ( .A(n1235), .B(n1193), .Z(G24) );
NAND3_X1 U910 ( .A1(n1236), .A2(n1028), .A3(n1220), .ZN(n1193) );
AND2_X1 U911 ( .A1(n1237), .A2(n1238), .ZN(n1220) );
XNOR2_X1 U912 ( .A(KEYINPUT50), .B(n1066), .ZN(n1237) );
NOR2_X1 U913 ( .A1(n1225), .A2(n1239), .ZN(n1028) );
XOR2_X1 U914 ( .A(KEYINPUT34), .B(n1226), .Z(n1239) );
XNOR2_X1 U915 ( .A(G119), .B(n1179), .ZN(G21) );
NAND4_X1 U916 ( .A1(n1236), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1179) );
INV_X1 U917 ( .A(n1039), .ZN(n1224) );
XNOR2_X1 U918 ( .A(G116), .B(n1180), .ZN(G18) );
OR2_X1 U919 ( .A1(n1240), .A2(n1187), .ZN(n1180) );
NAND2_X1 U920 ( .A1(n1066), .A2(n1238), .ZN(n1187) );
XNOR2_X1 U921 ( .A(n1241), .B(KEYINPUT33), .ZN(n1238) );
XOR2_X1 U922 ( .A(G113), .B(n1242), .Z(G15) );
NOR2_X1 U923 ( .A1(n1192), .A2(n1240), .ZN(n1242) );
NAND2_X1 U924 ( .A1(n1236), .A2(n1049), .ZN(n1240) );
INV_X1 U925 ( .A(n1190), .ZN(n1049) );
NAND2_X1 U926 ( .A1(n1243), .A2(n1225), .ZN(n1190) );
NOR2_X1 U927 ( .A1(n1188), .A2(n1047), .ZN(n1236) );
INV_X1 U928 ( .A(n1065), .ZN(n1047) );
NOR2_X1 U929 ( .A1(n1056), .A2(n1071), .ZN(n1065) );
INV_X1 U930 ( .A(n1206), .ZN(n1192) );
NOR2_X1 U931 ( .A1(n1241), .A2(n1066), .ZN(n1206) );
XOR2_X1 U932 ( .A(G110), .B(n1195), .Z(G12) );
AND2_X1 U933 ( .A1(n1231), .A2(n1048), .ZN(n1195) );
NOR2_X1 U934 ( .A1(n1225), .A2(n1243), .ZN(n1048) );
INV_X1 U935 ( .A(n1226), .ZN(n1243) );
NAND2_X1 U936 ( .A1(n1244), .A2(n1079), .ZN(n1226) );
NAND2_X1 U937 ( .A1(n1084), .A2(n1083), .ZN(n1079) );
OR2_X1 U938 ( .A1(n1083), .A2(n1084), .ZN(n1244) );
NOR2_X1 U939 ( .A1(n1127), .A2(G902), .ZN(n1084) );
XOR2_X1 U940 ( .A(n1245), .B(n1246), .Z(n1127) );
XOR2_X1 U941 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U942 ( .A1(G137), .A2(KEYINPUT20), .ZN(n1248) );
AND2_X1 U943 ( .A1(G221), .A2(n1249), .ZN(n1247) );
NAND2_X1 U944 ( .A1(n1250), .A2(n1251), .ZN(n1245) );
NAND2_X1 U945 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U946 ( .A(KEYINPUT41), .ZN(n1253) );
XNOR2_X1 U947 ( .A(n1254), .B(n1255), .ZN(n1252) );
NAND2_X1 U948 ( .A1(n1256), .A2(KEYINPUT41), .ZN(n1250) );
XOR2_X1 U949 ( .A(n1254), .B(n1257), .Z(n1256) );
NAND2_X1 U950 ( .A1(G146), .A2(n1258), .ZN(n1257) );
NAND3_X1 U951 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1254) );
OR2_X1 U952 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND3_X1 U953 ( .A1(n1263), .A2(n1262), .A3(G110), .ZN(n1260) );
NAND2_X1 U954 ( .A1(n1264), .A2(n1167), .ZN(n1259) );
INV_X1 U955 ( .A(G110), .ZN(n1167) );
NAND2_X1 U956 ( .A1(n1265), .A2(n1262), .ZN(n1264) );
INV_X1 U957 ( .A(KEYINPUT53), .ZN(n1262) );
XNOR2_X1 U958 ( .A(n1263), .B(KEYINPUT27), .ZN(n1265) );
XOR2_X1 U959 ( .A(G119), .B(n1266), .Z(n1263) );
XOR2_X1 U960 ( .A(KEYINPUT13), .B(G128), .Z(n1266) );
NAND2_X1 U961 ( .A1(G217), .A2(n1267), .ZN(n1083) );
XNOR2_X1 U962 ( .A(n1075), .B(G472), .ZN(n1225) );
NAND2_X1 U963 ( .A1(n1268), .A2(n1269), .ZN(n1075) );
XOR2_X1 U964 ( .A(n1144), .B(n1148), .Z(n1268) );
AND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1148) );
NAND2_X1 U966 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
INV_X1 U967 ( .A(G101), .ZN(n1273) );
NAND2_X1 U968 ( .A1(n1274), .A2(G210), .ZN(n1272) );
NAND3_X1 U969 ( .A1(n1274), .A2(G210), .A3(G101), .ZN(n1270) );
XOR2_X1 U970 ( .A(n1275), .B(n1276), .Z(n1144) );
XNOR2_X1 U971 ( .A(n1277), .B(n1278), .ZN(n1276) );
XOR2_X1 U972 ( .A(KEYINPUT38), .B(G113), .Z(n1278) );
XOR2_X1 U973 ( .A(n1279), .B(n1280), .Z(n1275) );
NOR3_X1 U974 ( .A1(n1188), .A2(n1022), .A3(n1039), .ZN(n1231) );
NAND2_X1 U975 ( .A1(n1066), .A2(n1281), .ZN(n1039) );
INV_X1 U976 ( .A(n1241), .ZN(n1281) );
NAND2_X1 U977 ( .A1(n1282), .A2(n1283), .ZN(n1241) );
OR2_X1 U978 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U979 ( .A(n1286), .B(KEYINPUT17), .Z(n1282) );
NAND2_X1 U980 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
INV_X1 U981 ( .A(G478), .ZN(n1284) );
XOR2_X1 U982 ( .A(n1085), .B(KEYINPUT63), .Z(n1285) );
NOR2_X1 U983 ( .A1(n1133), .A2(G902), .ZN(n1085) );
XNOR2_X1 U984 ( .A(n1287), .B(n1288), .ZN(n1133) );
XOR2_X1 U985 ( .A(n1289), .B(n1290), .Z(n1288) );
NAND2_X1 U986 ( .A1(G217), .A2(n1249), .ZN(n1290) );
AND2_X1 U987 ( .A1(G234), .A2(n1099), .ZN(n1249) );
NAND2_X1 U988 ( .A1(n1291), .A2(KEYINPUT28), .ZN(n1289) );
XNOR2_X1 U989 ( .A(G107), .B(n1292), .ZN(n1291) );
XOR2_X1 U990 ( .A(G122), .B(G116), .Z(n1292) );
XNOR2_X1 U991 ( .A(G134), .B(n1293), .ZN(n1287) );
NOR2_X1 U992 ( .A1(KEYINPUT22), .A2(n1294), .ZN(n1293) );
XOR2_X1 U993 ( .A(n1295), .B(G143), .Z(n1294) );
INV_X1 U994 ( .A(G128), .ZN(n1295) );
XOR2_X1 U995 ( .A(n1296), .B(G475), .Z(n1066) );
NAND2_X1 U996 ( .A1(n1137), .A2(n1269), .ZN(n1296) );
XNOR2_X1 U997 ( .A(n1297), .B(n1298), .ZN(n1137) );
NOR2_X1 U998 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U999 ( .A(KEYINPUT61), .B(n1301), .Z(n1300) );
NOR2_X1 U1000 ( .A1(n1255), .A2(n1302), .ZN(n1301) );
AND2_X1 U1001 ( .A1(n1302), .A2(n1255), .ZN(n1299) );
XOR2_X1 U1002 ( .A(G146), .B(n1258), .Z(n1255) );
XOR2_X1 U1003 ( .A(G125), .B(G140), .Z(n1258) );
NAND2_X1 U1004 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U1005 ( .A1(n1305), .A2(G131), .ZN(n1304) );
XOR2_X1 U1006 ( .A(n1306), .B(KEYINPUT62), .Z(n1303) );
OR2_X1 U1007 ( .A1(n1305), .A2(G131), .ZN(n1306) );
XNOR2_X1 U1008 ( .A(n1307), .B(n1219), .ZN(n1305) );
NAND2_X1 U1009 ( .A1(n1274), .A2(G214), .ZN(n1307) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1274) );
NAND3_X1 U1011 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1297) );
OR2_X1 U1012 ( .A1(n1142), .A2(KEYINPUT18), .ZN(n1310) );
NAND3_X1 U1013 ( .A1(KEYINPUT18), .A2(n1142), .A3(n1311), .ZN(n1309) );
INV_X1 U1014 ( .A(n1312), .ZN(n1311) );
INV_X1 U1015 ( .A(G104), .ZN(n1142) );
NAND2_X1 U1016 ( .A1(n1312), .A2(n1313), .ZN(n1308) );
NAND2_X1 U1017 ( .A1(KEYINPUT18), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1018 ( .A(KEYINPUT3), .B(G104), .Z(n1314) );
XOR2_X1 U1019 ( .A(n1315), .B(G113), .Z(n1312) );
NAND2_X1 U1020 ( .A1(KEYINPUT5), .A2(n1235), .ZN(n1315) );
NAND2_X1 U1021 ( .A1(n1316), .A2(n1056), .ZN(n1022) );
XNOR2_X1 U1022 ( .A(n1077), .B(n1317), .ZN(n1056) );
NOR2_X1 U1023 ( .A1(KEYINPUT29), .A2(n1078), .ZN(n1317) );
INV_X1 U1024 ( .A(G469), .ZN(n1078) );
NAND2_X1 U1025 ( .A1(n1318), .A2(n1269), .ZN(n1077) );
XOR2_X1 U1026 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1027 ( .A(n1321), .B(n1322), .ZN(n1320) );
NOR2_X1 U1028 ( .A1(G110), .A2(KEYINPUT48), .ZN(n1322) );
NOR2_X1 U1029 ( .A1(KEYINPUT47), .A2(n1160), .ZN(n1321) );
XNOR2_X1 U1030 ( .A(n1323), .B(n1324), .ZN(n1160) );
XOR2_X1 U1031 ( .A(n1279), .B(n1123), .Z(n1324) );
XOR2_X1 U1032 ( .A(n1095), .B(KEYINPUT43), .Z(n1279) );
XOR2_X1 U1033 ( .A(n1325), .B(n1326), .Z(n1095) );
XOR2_X1 U1034 ( .A(G137), .B(G134), .Z(n1326) );
XNOR2_X1 U1035 ( .A(G131), .B(n1327), .ZN(n1325) );
XOR2_X1 U1036 ( .A(n1219), .B(KEYINPUT10), .Z(n1323) );
XOR2_X1 U1037 ( .A(n1097), .B(n1161), .Z(n1319) );
AND2_X1 U1038 ( .A1(G227), .A2(n1099), .ZN(n1161) );
INV_X1 U1039 ( .A(G140), .ZN(n1097) );
XOR2_X1 U1040 ( .A(KEYINPUT58), .B(n1071), .Z(n1316) );
INV_X1 U1041 ( .A(n1055), .ZN(n1071) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1267), .ZN(n1055) );
NAND2_X1 U1043 ( .A1(n1328), .A2(n1269), .ZN(n1267) );
NAND2_X1 U1044 ( .A1(n1060), .A2(n1026), .ZN(n1188) );
NAND2_X1 U1045 ( .A1(n1035), .A2(n1329), .ZN(n1026) );
NAND3_X1 U1046 ( .A1(n1119), .A2(n1234), .A3(G902), .ZN(n1329) );
NOR2_X1 U1047 ( .A1(n1099), .A2(G898), .ZN(n1119) );
NAND3_X1 U1048 ( .A1(n1234), .A2(n1099), .A3(G952), .ZN(n1035) );
INV_X1 U1049 ( .A(G953), .ZN(n1099) );
NAND2_X1 U1050 ( .A1(G237), .A2(n1328), .ZN(n1234) );
XOR2_X1 U1051 ( .A(G234), .B(KEYINPUT46), .Z(n1328) );
INV_X1 U1052 ( .A(n1024), .ZN(n1060) );
NAND2_X1 U1053 ( .A1(n1062), .A2(n1228), .ZN(n1024) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1330), .ZN(n1228) );
XOR2_X1 U1055 ( .A(n1331), .B(n1177), .Z(n1062) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1330), .ZN(n1177) );
NAND2_X1 U1057 ( .A1(n1332), .A2(n1269), .ZN(n1330) );
INV_X1 U1058 ( .A(G237), .ZN(n1332) );
NAND2_X1 U1059 ( .A1(n1333), .A2(n1269), .ZN(n1331) );
INV_X1 U1060 ( .A(G902), .ZN(n1269) );
XNOR2_X1 U1061 ( .A(n1334), .B(n1173), .ZN(n1333) );
XNOR2_X1 U1062 ( .A(n1335), .B(n1121), .ZN(n1173) );
XOR2_X1 U1063 ( .A(n1336), .B(n1235), .Z(n1121) );
INV_X1 U1064 ( .A(G122), .ZN(n1235) );
NAND2_X1 U1065 ( .A1(KEYINPUT9), .A2(G110), .ZN(n1336) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1335) );
INV_X1 U1067 ( .A(n1123), .ZN(n1338) );
XOR2_X1 U1068 ( .A(n1339), .B(n1340), .Z(n1123) );
XOR2_X1 U1069 ( .A(G104), .B(G101), .Z(n1340) );
XNOR2_X1 U1070 ( .A(G107), .B(KEYINPUT16), .ZN(n1339) );
NAND2_X1 U1071 ( .A1(KEYINPUT54), .A2(n1124), .ZN(n1337) );
XOR2_X1 U1072 ( .A(G113), .B(n1341), .Z(n1124) );
NOR2_X1 U1073 ( .A1(KEYINPUT4), .A2(n1280), .ZN(n1341) );
XOR2_X1 U1074 ( .A(G116), .B(G119), .Z(n1280) );
NAND3_X1 U1075 ( .A1(n1342), .A2(n1343), .A3(n1344), .ZN(n1334) );
NAND2_X1 U1076 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
OR3_X1 U1077 ( .A1(n1346), .A2(n1345), .A3(KEYINPUT57), .ZN(n1343) );
AND2_X1 U1078 ( .A1(KEYINPUT7), .A2(n1211), .ZN(n1345) );
NAND2_X1 U1079 ( .A1(KEYINPUT57), .A2(n1347), .ZN(n1342) );
OR2_X1 U1080 ( .A1(n1346), .A2(n1211), .ZN(n1347) );
NOR2_X1 U1081 ( .A1(n1113), .A2(G953), .ZN(n1211) );
INV_X1 U1082 ( .A(G224), .ZN(n1113) );
XOR2_X1 U1083 ( .A(n1210), .B(G125), .Z(n1346) );
XNOR2_X1 U1084 ( .A(n1277), .B(n1327), .ZN(n1210) );
XOR2_X1 U1085 ( .A(G128), .B(G146), .Z(n1327) );
NAND2_X1 U1086 ( .A1(KEYINPUT1), .A2(n1219), .ZN(n1277) );
INV_X1 U1087 ( .A(G143), .ZN(n1219) );
endmodule


