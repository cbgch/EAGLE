//Key = 1111000100010110011101010001101110110111101111100111010001101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287;

XOR2_X1 U709 ( .A(G107), .B(n970), .Z(G9) );
NOR2_X1 U710 ( .A1(n971), .A2(n972), .ZN(G75) );
XOR2_X1 U711 ( .A(KEYINPUT55), .B(n973), .Z(n972) );
NOR4_X1 U712 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .ZN(n973) );
NOR3_X1 U713 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NOR2_X1 U714 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR2_X1 U715 ( .A1(n983), .A2(n984), .ZN(n982) );
NOR3_X1 U716 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n983) );
AND3_X1 U717 ( .A1(n988), .A2(n989), .A3(G214), .ZN(n987) );
INV_X1 U718 ( .A(n990), .ZN(n988) );
NOR2_X1 U719 ( .A1(n991), .A2(n992), .ZN(n985) );
NOR3_X1 U720 ( .A1(n993), .A2(n991), .A3(n994), .ZN(n981) );
NAND3_X1 U721 ( .A1(n995), .A2(n992), .A3(G221), .ZN(n993) );
INV_X1 U722 ( .A(KEYINPUT52), .ZN(n992) );
NOR2_X1 U723 ( .A1(n996), .A2(n991), .ZN(n975) );
NOR3_X1 U724 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NOR4_X1 U725 ( .A1(n1000), .A2(n984), .A3(n980), .A4(n1001), .ZN(n999) );
NOR2_X1 U726 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR2_X1 U727 ( .A1(n1004), .A2(n978), .ZN(n998) );
NOR3_X1 U728 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NOR2_X1 U729 ( .A1(n1008), .A2(n984), .ZN(n1007) );
INV_X1 U730 ( .A(n1009), .ZN(n984) );
AND2_X1 U731 ( .A1(n1010), .A2(KEYINPUT0), .ZN(n1006) );
NOR2_X1 U732 ( .A1(n1011), .A2(n980), .ZN(n1005) );
NOR2_X1 U733 ( .A1(n1012), .A2(KEYINPUT0), .ZN(n997) );
NOR2_X1 U734 ( .A1(n1013), .A2(n978), .ZN(n1012) );
OR2_X1 U735 ( .A1(n1001), .A2(n1014), .ZN(n978) );
OR2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n974) );
NOR3_X1 U737 ( .A1(n1015), .A2(G952), .A3(n976), .ZN(n971) );
AND4_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1009), .A4(n1019), .ZN(n976) );
NOR3_X1 U739 ( .A1(n991), .A2(n1020), .A3(n1021), .ZN(n1019) );
XOR2_X1 U740 ( .A(n1022), .B(KEYINPUT34), .Z(n1020) );
INV_X1 U741 ( .A(n1023), .ZN(n991) );
OR2_X1 U742 ( .A1(n1024), .A2(KEYINPUT23), .ZN(n1018) );
NAND2_X1 U743 ( .A1(KEYINPUT23), .A2(n980), .ZN(n1017) );
XOR2_X1 U744 ( .A(n1025), .B(n1026), .Z(G72) );
XOR2_X1 U745 ( .A(n1027), .B(n1028), .Z(n1026) );
NOR2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
XOR2_X1 U747 ( .A(n1031), .B(n1032), .Z(n1030) );
NOR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR3_X1 U749 ( .A1(n1035), .A2(KEYINPUT63), .A3(n1036), .ZN(n1034) );
NOR2_X1 U750 ( .A1(G125), .A2(n1037), .ZN(n1033) );
NOR2_X1 U751 ( .A1(KEYINPUT63), .A2(n1036), .ZN(n1037) );
NAND2_X1 U752 ( .A1(n1038), .A2(KEYINPUT28), .ZN(n1031) );
XOR2_X1 U753 ( .A(n1039), .B(n1040), .Z(n1038) );
XNOR2_X1 U754 ( .A(n1041), .B(n1042), .ZN(n1040) );
INV_X1 U755 ( .A(G131), .ZN(n1041) );
NOR2_X1 U756 ( .A1(n1043), .A2(n1044), .ZN(n1039) );
NOR2_X1 U757 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XNOR2_X1 U758 ( .A(KEYINPUT20), .B(n1047), .ZN(n1045) );
INV_X1 U759 ( .A(G134), .ZN(n1047) );
NOR2_X1 U760 ( .A1(G137), .A2(n1048), .ZN(n1043) );
XNOR2_X1 U761 ( .A(G134), .B(KEYINPUT24), .ZN(n1048) );
NAND2_X1 U762 ( .A1(n1049), .A2(n1050), .ZN(n1027) );
NAND2_X1 U763 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U764 ( .A(n1053), .B(KEYINPUT6), .Z(n1051) );
XNOR2_X1 U765 ( .A(KEYINPUT44), .B(n1054), .ZN(n1049) );
NAND3_X1 U766 ( .A1(G953), .A2(n1055), .A3(KEYINPUT30), .ZN(n1025) );
NAND2_X1 U767 ( .A1(G900), .A2(G227), .ZN(n1055) );
NAND2_X1 U768 ( .A1(n1056), .A2(n1057), .ZN(G69) );
NAND2_X1 U769 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U770 ( .A1(n1060), .A2(n1061), .ZN(n1056) );
NAND2_X1 U771 ( .A1(n1062), .A2(n1059), .ZN(n1061) );
NAND2_X1 U772 ( .A1(G953), .A2(n1063), .ZN(n1059) );
INV_X1 U773 ( .A(G224), .ZN(n1063) );
INV_X1 U774 ( .A(n1064), .ZN(n1062) );
INV_X1 U775 ( .A(n1058), .ZN(n1060) );
XNOR2_X1 U776 ( .A(n1065), .B(n1066), .ZN(n1058) );
NOR2_X1 U777 ( .A1(n1064), .A2(n1067), .ZN(n1066) );
XOR2_X1 U778 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U779 ( .A1(n1070), .A2(n1054), .ZN(n1065) );
NOR2_X1 U780 ( .A1(n1071), .A2(n1072), .ZN(G66) );
XOR2_X1 U781 ( .A(n1073), .B(n1074), .Z(n1072) );
XNOR2_X1 U782 ( .A(n1075), .B(KEYINPUT43), .ZN(n1074) );
NAND3_X1 U783 ( .A1(n1076), .A2(n1077), .A3(KEYINPUT37), .ZN(n1075) );
NOR2_X1 U784 ( .A1(n1071), .A2(n1078), .ZN(G63) );
XOR2_X1 U785 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U786 ( .A1(n1076), .A2(G478), .ZN(n1079) );
NOR2_X1 U787 ( .A1(n1071), .A2(n1081), .ZN(G60) );
XOR2_X1 U788 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND2_X1 U789 ( .A1(n1076), .A2(G475), .ZN(n1082) );
XOR2_X1 U790 ( .A(G104), .B(n1084), .Z(G6) );
NOR2_X1 U791 ( .A1(n1071), .A2(n1085), .ZN(G57) );
XOR2_X1 U792 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U793 ( .A(n1088), .B(n1089), .Z(n1087) );
XNOR2_X1 U794 ( .A(n1090), .B(n1091), .ZN(n1086) );
XOR2_X1 U795 ( .A(n1092), .B(n1093), .Z(n1090) );
NOR2_X1 U796 ( .A1(KEYINPUT10), .A2(n1094), .ZN(n1093) );
NAND2_X1 U797 ( .A1(n1076), .A2(G472), .ZN(n1092) );
NOR2_X1 U798 ( .A1(n1071), .A2(n1095), .ZN(G54) );
XOR2_X1 U799 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U800 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U801 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U802 ( .A1(KEYINPUT33), .A2(n1102), .ZN(n1101) );
XNOR2_X1 U803 ( .A(G140), .B(KEYINPUT3), .ZN(n1102) );
NAND3_X1 U804 ( .A1(n1076), .A2(G469), .A3(n1103), .ZN(n1100) );
XNOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT1), .ZN(n1103) );
NAND2_X1 U806 ( .A1(n1104), .A2(KEYINPUT14), .ZN(n1098) );
XOR2_X1 U807 ( .A(n1105), .B(KEYINPUT35), .Z(n1104) );
XNOR2_X1 U808 ( .A(n1106), .B(n1107), .ZN(n1096) );
XNOR2_X1 U809 ( .A(n1108), .B(n1109), .ZN(n1106) );
NOR2_X1 U810 ( .A1(n1071), .A2(n1110), .ZN(G51) );
NOR2_X1 U811 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U812 ( .A(KEYINPUT12), .B(n1113), .Z(n1112) );
NOR2_X1 U813 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U814 ( .A(n1116), .B(KEYINPUT32), .Z(n1114) );
NOR2_X1 U815 ( .A1(n1117), .A2(n1116), .ZN(n1111) );
NAND2_X1 U816 ( .A1(n1076), .A2(n1118), .ZN(n1116) );
AND2_X1 U817 ( .A1(G902), .A2(n1016), .ZN(n1076) );
NAND3_X1 U818 ( .A1(n1119), .A2(n1053), .A3(n1052), .ZN(n1016) );
AND4_X1 U819 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1052) );
AND4_X1 U820 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
NAND3_X1 U821 ( .A1(n1024), .A2(n986), .A3(n1128), .ZN(n1122) );
NAND3_X1 U822 ( .A1(n1129), .A2(n1023), .A3(n1130), .ZN(n1120) );
INV_X1 U823 ( .A(n1070), .ZN(n1119) );
NAND4_X1 U824 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1070) );
NOR4_X1 U825 ( .A1(n1135), .A2(n1136), .A3(n970), .A4(n1084), .ZN(n1134) );
AND3_X1 U826 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1084) );
AND3_X1 U827 ( .A1(n1137), .A2(n1138), .A3(n1024), .ZN(n970) );
OR2_X1 U828 ( .A1(n1140), .A2(KEYINPUT56), .ZN(n1133) );
NAND2_X1 U829 ( .A1(n986), .A2(n1141), .ZN(n1132) );
NAND2_X1 U830 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U831 ( .A1(KEYINPUT56), .A2(n1144), .ZN(n1143) );
NAND3_X1 U832 ( .A1(n1009), .A2(n1145), .A3(n1146), .ZN(n1144) );
XOR2_X1 U833 ( .A(n1147), .B(KEYINPUT25), .Z(n1142) );
NAND2_X1 U834 ( .A1(n1148), .A2(n1149), .ZN(n1131) );
NAND3_X1 U835 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
OR3_X1 U836 ( .A1(n1153), .A2(n1154), .A3(n1014), .ZN(n1152) );
OR2_X1 U837 ( .A1(n1155), .A2(KEYINPUT29), .ZN(n1151) );
NAND3_X1 U838 ( .A1(n1139), .A2(n1156), .A3(KEYINPUT29), .ZN(n1150) );
NOR2_X1 U839 ( .A1(n1054), .A2(G952), .ZN(n1071) );
XOR2_X1 U840 ( .A(n1053), .B(n1157), .Z(G48) );
XNOR2_X1 U841 ( .A(G146), .B(KEYINPUT8), .ZN(n1157) );
NAND3_X1 U842 ( .A1(n1128), .A2(n986), .A3(n1139), .ZN(n1053) );
XNOR2_X1 U843 ( .A(n1121), .B(n1158), .ZN(G45) );
NOR2_X1 U844 ( .A1(KEYINPUT36), .A2(n1159), .ZN(n1158) );
NAND3_X1 U845 ( .A1(n1003), .A2(n1129), .A3(n1160), .ZN(n1121) );
NOR3_X1 U846 ( .A1(n1161), .A2(n1154), .A3(n1153), .ZN(n1160) );
XNOR2_X1 U847 ( .A(G140), .B(n1127), .ZN(G42) );
NAND4_X1 U848 ( .A1(n1002), .A2(n1139), .A3(n1129), .A4(n1023), .ZN(n1127) );
XNOR2_X1 U849 ( .A(G137), .B(n1125), .ZN(G39) );
NAND3_X1 U850 ( .A1(n1128), .A2(n1023), .A3(n1162), .ZN(n1125) );
NAND3_X1 U851 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(G36) );
OR2_X1 U852 ( .A1(G134), .A2(KEYINPUT61), .ZN(n1165) );
NAND3_X1 U853 ( .A1(KEYINPUT61), .A2(G134), .A3(n1126), .ZN(n1164) );
NAND2_X1 U854 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NAND2_X1 U855 ( .A1(n1168), .A2(KEYINPUT61), .ZN(n1167) );
XNOR2_X1 U856 ( .A(G134), .B(KEYINPUT40), .ZN(n1168) );
INV_X1 U857 ( .A(n1126), .ZN(n1166) );
NAND4_X1 U858 ( .A1(n1003), .A2(n1129), .A3(n1023), .A4(n1024), .ZN(n1126) );
XNOR2_X1 U859 ( .A(G131), .B(n1169), .ZN(G33) );
NAND4_X1 U860 ( .A1(n1170), .A2(n1130), .A3(n1023), .A4(n1171), .ZN(n1169) );
NOR2_X1 U861 ( .A1(n990), .A2(n1172), .ZN(n1023) );
AND2_X1 U862 ( .A1(G214), .A2(n989), .ZN(n1172) );
INV_X1 U863 ( .A(n1155), .ZN(n1130) );
XOR2_X1 U864 ( .A(n1173), .B(KEYINPUT9), .Z(n1170) );
XNOR2_X1 U865 ( .A(G128), .B(n1174), .ZN(G30) );
NAND3_X1 U866 ( .A1(n1128), .A2(n1024), .A3(n1175), .ZN(n1174) );
XNOR2_X1 U867 ( .A(n986), .B(KEYINPUT58), .ZN(n1175) );
INV_X1 U868 ( .A(n1008), .ZN(n1024) );
AND3_X1 U869 ( .A1(n1176), .A2(n1177), .A3(n1129), .ZN(n1128) );
AND2_X1 U870 ( .A1(n1171), .A2(n1173), .ZN(n1129) );
XNOR2_X1 U871 ( .A(n1178), .B(n1136), .ZN(G3) );
AND3_X1 U872 ( .A1(n1162), .A2(n1138), .A3(n1003), .ZN(n1136) );
AND3_X1 U873 ( .A1(n1171), .A2(n1145), .A3(n986), .ZN(n1138) );
NAND2_X1 U874 ( .A1(n1179), .A2(n1180), .ZN(G27) );
NAND2_X1 U875 ( .A1(n1181), .A2(n1035), .ZN(n1180) );
XOR2_X1 U876 ( .A(KEYINPUT38), .B(n1182), .Z(n1179) );
NOR2_X1 U877 ( .A1(n1181), .A2(n1035), .ZN(n1182) );
INV_X1 U878 ( .A(n1124), .ZN(n1181) );
NAND4_X1 U879 ( .A1(n1010), .A2(n1002), .A3(n986), .A4(n1173), .ZN(n1124) );
NAND2_X1 U880 ( .A1(n1183), .A2(n1001), .ZN(n1173) );
NAND2_X1 U881 ( .A1(n1029), .A2(n1184), .ZN(n1183) );
NOR2_X1 U882 ( .A1(n1054), .A2(G900), .ZN(n1029) );
INV_X1 U883 ( .A(n1013), .ZN(n1010) );
NAND2_X1 U884 ( .A1(n1139), .A2(n1009), .ZN(n1013) );
XNOR2_X1 U885 ( .A(G122), .B(n1185), .ZN(G24) );
NAND3_X1 U886 ( .A1(KEYINPUT53), .A2(n1148), .A3(n1186), .ZN(n1185) );
NOR3_X1 U887 ( .A1(n1014), .A2(n1154), .A3(n1153), .ZN(n1186) );
INV_X1 U888 ( .A(n1137), .ZN(n1014) );
NOR2_X1 U889 ( .A1(n1021), .A2(n1177), .ZN(n1137) );
XOR2_X1 U890 ( .A(n1140), .B(n1187), .Z(G21) );
NAND2_X1 U891 ( .A1(KEYINPUT42), .A2(G119), .ZN(n1187) );
NAND2_X1 U892 ( .A1(n1146), .A2(n1148), .ZN(n1140) );
INV_X1 U893 ( .A(n1188), .ZN(n1148) );
AND3_X1 U894 ( .A1(n1176), .A2(n1177), .A3(n1162), .ZN(n1146) );
INV_X1 U895 ( .A(n1022), .ZN(n1177) );
XOR2_X1 U896 ( .A(n1135), .B(n1189), .Z(G18) );
NOR2_X1 U897 ( .A1(KEYINPUT59), .A2(n1190), .ZN(n1189) );
NOR3_X1 U898 ( .A1(n1156), .A2(n1008), .A3(n1188), .ZN(n1135) );
NAND2_X1 U899 ( .A1(n1153), .A2(n1191), .ZN(n1008) );
XOR2_X1 U900 ( .A(n1192), .B(n1193), .Z(G15) );
NOR2_X1 U901 ( .A1(n1155), .A2(n1188), .ZN(n1193) );
NAND3_X1 U902 ( .A1(n986), .A2(n1145), .A3(n1009), .ZN(n1188) );
NOR2_X1 U903 ( .A1(n994), .A2(n1194), .ZN(n1009) );
AND2_X1 U904 ( .A1(G221), .A2(n995), .ZN(n1194) );
INV_X1 U905 ( .A(n1161), .ZN(n986) );
NAND2_X1 U906 ( .A1(n1003), .A2(n1139), .ZN(n1155) );
NOR2_X1 U907 ( .A1(n1191), .A2(n1153), .ZN(n1139) );
INV_X1 U908 ( .A(n1156), .ZN(n1003) );
NAND2_X1 U909 ( .A1(n1022), .A2(n1176), .ZN(n1156) );
XOR2_X1 U910 ( .A(n1021), .B(KEYINPUT62), .Z(n1176) );
XNOR2_X1 U911 ( .A(G113), .B(KEYINPUT18), .ZN(n1192) );
XOR2_X1 U912 ( .A(G110), .B(n1195), .Z(G12) );
NOR2_X1 U913 ( .A1(n1161), .A2(n1147), .ZN(n1195) );
NAND4_X1 U914 ( .A1(n1162), .A2(n1002), .A3(n1171), .A4(n1145), .ZN(n1147) );
NAND2_X1 U915 ( .A1(n1196), .A2(n1001), .ZN(n1145) );
NAND3_X1 U916 ( .A1(n1197), .A2(n1198), .A3(G952), .ZN(n1001) );
INV_X1 U917 ( .A(n1015), .ZN(n1197) );
XOR2_X1 U918 ( .A(G953), .B(KEYINPUT22), .Z(n1015) );
NAND2_X1 U919 ( .A1(n1064), .A2(n1184), .ZN(n1196) );
AND2_X1 U920 ( .A1(G902), .A2(n1198), .ZN(n1184) );
NAND2_X1 U921 ( .A1(G237), .A2(n1199), .ZN(n1198) );
NOR2_X1 U922 ( .A1(G898), .A2(n1054), .ZN(n1064) );
INV_X1 U923 ( .A(n1011), .ZN(n1171) );
NAND2_X1 U924 ( .A1(n994), .A2(n1200), .ZN(n1011) );
NAND2_X1 U925 ( .A1(G221), .A2(n995), .ZN(n1200) );
XNOR2_X1 U926 ( .A(n1201), .B(G469), .ZN(n994) );
NAND2_X1 U927 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U928 ( .A(n1204), .B(n1205), .Z(n1202) );
XNOR2_X1 U929 ( .A(n1206), .B(n1105), .ZN(n1205) );
NAND2_X1 U930 ( .A1(G227), .A2(n1054), .ZN(n1105) );
NAND2_X1 U931 ( .A1(KEYINPUT39), .A2(n1107), .ZN(n1206) );
XNOR2_X1 U932 ( .A(n1207), .B(n1036), .ZN(n1204) );
NAND2_X1 U933 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U934 ( .A1(n1210), .A2(n1091), .ZN(n1209) );
XOR2_X1 U935 ( .A(KEYINPUT2), .B(n1211), .Z(n1208) );
NOR2_X1 U936 ( .A1(n1091), .A2(n1210), .ZN(n1211) );
XNOR2_X1 U937 ( .A(KEYINPUT4), .B(n1109), .ZN(n1210) );
XNOR2_X1 U938 ( .A(n1212), .B(n1042), .ZN(n1109) );
XNOR2_X1 U939 ( .A(n1213), .B(n1214), .ZN(n1042) );
NOR2_X1 U940 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U941 ( .A(KEYINPUT16), .B(n1217), .Z(n1216) );
AND2_X1 U942 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR2_X1 U943 ( .A1(n1218), .A2(n1219), .ZN(n1215) );
XOR2_X1 U944 ( .A(G143), .B(KEYINPUT15), .Z(n1219) );
NAND2_X1 U945 ( .A1(KEYINPUT11), .A2(n1220), .ZN(n1213) );
INV_X1 U946 ( .A(n1108), .ZN(n1091) );
NOR2_X1 U947 ( .A1(n1021), .A2(n1022), .ZN(n1002) );
XOR2_X1 U948 ( .A(n1221), .B(n1077), .Z(n1022) );
AND2_X1 U949 ( .A1(G217), .A2(n995), .ZN(n1077) );
NAND2_X1 U950 ( .A1(n1222), .A2(n1199), .ZN(n995) );
XOR2_X1 U951 ( .A(G234), .B(KEYINPUT5), .Z(n1199) );
NAND2_X1 U952 ( .A1(n1073), .A2(n1203), .ZN(n1221) );
XNOR2_X1 U953 ( .A(n1223), .B(n1224), .ZN(n1073) );
XNOR2_X1 U954 ( .A(n1225), .B(KEYINPUT27), .ZN(n1224) );
NAND2_X1 U955 ( .A1(n1226), .A2(KEYINPUT60), .ZN(n1225) );
XOR2_X1 U956 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U957 ( .A(KEYINPUT45), .B(n1046), .ZN(n1228) );
NAND2_X1 U958 ( .A1(G221), .A2(n1229), .ZN(n1227) );
XNOR2_X1 U959 ( .A(n1230), .B(n1231), .ZN(n1223) );
NOR2_X1 U960 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NOR3_X1 U961 ( .A1(G125), .A2(G140), .A3(n1234), .ZN(n1233) );
NOR2_X1 U962 ( .A1(n1235), .A2(n1035), .ZN(n1232) );
NOR2_X1 U963 ( .A1(G140), .A2(n1234), .ZN(n1235) );
INV_X1 U964 ( .A(KEYINPUT21), .ZN(n1234) );
XNOR2_X1 U965 ( .A(n1236), .B(n1237), .ZN(n1021) );
XOR2_X1 U966 ( .A(KEYINPUT54), .B(G472), .Z(n1237) );
NAND2_X1 U967 ( .A1(n1238), .A2(n1203), .ZN(n1236) );
XOR2_X1 U968 ( .A(n1239), .B(n1089), .Z(n1238) );
AND2_X1 U969 ( .A1(n1240), .A2(n1241), .ZN(n1089) );
NAND2_X1 U970 ( .A1(n1242), .A2(n1178), .ZN(n1241) );
INV_X1 U971 ( .A(G101), .ZN(n1178) );
NAND3_X1 U972 ( .A1(n1243), .A2(n1054), .A3(G210), .ZN(n1242) );
NAND4_X1 U973 ( .A1(n1243), .A2(n1054), .A3(G210), .A4(G101), .ZN(n1240) );
NOR2_X1 U974 ( .A1(n1244), .A2(n1245), .ZN(n1239) );
XOR2_X1 U975 ( .A(n1246), .B(KEYINPUT19), .Z(n1245) );
NAND2_X1 U976 ( .A1(n1088), .A2(n1247), .ZN(n1246) );
NOR2_X1 U977 ( .A1(n1088), .A2(n1247), .ZN(n1244) );
NAND3_X1 U978 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
NAND2_X1 U979 ( .A1(KEYINPUT26), .A2(n1251), .ZN(n1250) );
NAND3_X1 U980 ( .A1(n1252), .A2(n1253), .A3(n1108), .ZN(n1249) );
INV_X1 U981 ( .A(KEYINPUT26), .ZN(n1253) );
OR2_X1 U982 ( .A1(n1108), .A2(n1252), .ZN(n1248) );
NOR2_X1 U983 ( .A1(KEYINPUT41), .A2(n1251), .ZN(n1252) );
XOR2_X1 U984 ( .A(n1094), .B(KEYINPUT13), .Z(n1251) );
XOR2_X1 U985 ( .A(n1254), .B(n1255), .Z(n1094) );
XOR2_X1 U986 ( .A(G131), .B(n1256), .Z(n1108) );
XNOR2_X1 U987 ( .A(n1046), .B(G134), .ZN(n1256) );
INV_X1 U988 ( .A(G137), .ZN(n1046) );
XNOR2_X1 U989 ( .A(n1257), .B(G113), .ZN(n1088) );
NAND2_X1 U990 ( .A1(KEYINPUT7), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U991 ( .A(G119), .B(n1190), .ZN(n1258) );
INV_X1 U992 ( .A(n980), .ZN(n1162) );
NAND2_X1 U993 ( .A1(n1154), .A2(n1153), .ZN(n980) );
XOR2_X1 U994 ( .A(n1259), .B(G475), .Z(n1153) );
NAND2_X1 U995 ( .A1(n1083), .A2(n1203), .ZN(n1259) );
XNOR2_X1 U996 ( .A(n1260), .B(n1261), .ZN(n1083) );
XOR2_X1 U997 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U998 ( .A(n1036), .B(G131), .ZN(n1263) );
INV_X1 U999 ( .A(G140), .ZN(n1036) );
XNOR2_X1 U1000 ( .A(n1218), .B(G143), .ZN(n1262) );
INV_X1 U1001 ( .A(G146), .ZN(n1218) );
XOR2_X1 U1002 ( .A(n1264), .B(n1265), .Z(n1260) );
XNOR2_X1 U1003 ( .A(n1035), .B(G104), .ZN(n1265) );
XNOR2_X1 U1004 ( .A(n1266), .B(n1267), .ZN(n1264) );
NAND4_X1 U1005 ( .A1(KEYINPUT31), .A2(G214), .A3(n1243), .A4(n1054), .ZN(n1267) );
NAND2_X1 U1006 ( .A1(KEYINPUT17), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U1007 ( .A(G122), .B(n1269), .ZN(n1268) );
INV_X1 U1008 ( .A(n1191), .ZN(n1154) );
XNOR2_X1 U1009 ( .A(n1270), .B(G478), .ZN(n1191) );
NAND2_X1 U1010 ( .A1(n1080), .A2(n1203), .ZN(n1270) );
XNOR2_X1 U1011 ( .A(n1271), .B(n1272), .ZN(n1080) );
XOR2_X1 U1012 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U1013 ( .A(n1159), .B(G134), .ZN(n1274) );
INV_X1 U1014 ( .A(G143), .ZN(n1159) );
XOR2_X1 U1015 ( .A(KEYINPUT50), .B(KEYINPUT46), .Z(n1273) );
XOR2_X1 U1016 ( .A(n1275), .B(n1276), .Z(n1271) );
XNOR2_X1 U1017 ( .A(n1220), .B(G107), .ZN(n1276) );
XOR2_X1 U1018 ( .A(n1277), .B(n1278), .Z(n1275) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1229), .ZN(n1277) );
AND2_X1 U1020 ( .A1(G234), .A2(n1054), .ZN(n1229) );
NAND2_X1 U1021 ( .A1(n990), .A2(n1279), .ZN(n1161) );
NAND2_X1 U1022 ( .A1(G214), .A2(n989), .ZN(n1279) );
XNOR2_X1 U1023 ( .A(n1280), .B(n1118), .ZN(n990) );
AND2_X1 U1024 ( .A1(G210), .A2(n989), .ZN(n1118) );
NAND2_X1 U1025 ( .A1(n1222), .A2(n1243), .ZN(n989) );
INV_X1 U1026 ( .A(G237), .ZN(n1243) );
XNOR2_X1 U1027 ( .A(G902), .B(KEYINPUT47), .ZN(n1222) );
NAND2_X1 U1028 ( .A1(n1117), .A2(n1203), .ZN(n1280) );
INV_X1 U1029 ( .A(G902), .ZN(n1203) );
INV_X1 U1030 ( .A(n1115), .ZN(n1117) );
XNOR2_X1 U1031 ( .A(n1281), .B(n1282), .ZN(n1115) );
XOR2_X1 U1032 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U1033 ( .A(n1254), .B(n1035), .ZN(n1284) );
INV_X1 U1034 ( .A(G125), .ZN(n1035) );
NAND2_X1 U1035 ( .A1(KEYINPUT51), .A2(G143), .ZN(n1254) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1054), .ZN(n1283) );
INV_X1 U1037 ( .A(G953), .ZN(n1054) );
XOR2_X1 U1038 ( .A(n1068), .B(n1230), .Z(n1281) );
XOR2_X1 U1039 ( .A(n1069), .B(n1255), .Z(n1230) );
XNOR2_X1 U1040 ( .A(n1220), .B(G146), .ZN(n1255) );
INV_X1 U1041 ( .A(G128), .ZN(n1220) );
XNOR2_X1 U1042 ( .A(G119), .B(n1107), .ZN(n1069) );
XNOR2_X1 U1043 ( .A(G110), .B(KEYINPUT49), .ZN(n1107) );
XOR2_X1 U1044 ( .A(n1285), .B(n1286), .Z(n1068) );
XNOR2_X1 U1045 ( .A(KEYINPUT48), .B(n1269), .ZN(n1286) );
INV_X1 U1046 ( .A(G113), .ZN(n1269) );
XOR2_X1 U1047 ( .A(n1212), .B(n1278), .Z(n1285) );
XNOR2_X1 U1048 ( .A(n1190), .B(G122), .ZN(n1278) );
INV_X1 U1049 ( .A(G116), .ZN(n1190) );
XNOR2_X1 U1050 ( .A(G101), .B(n1287), .ZN(n1212) );
XOR2_X1 U1051 ( .A(G107), .B(G104), .Z(n1287) );
endmodule


