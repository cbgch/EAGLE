//Key = 1111010111011100011111011111100110100001011101010000011110110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388;

XOR2_X1 U755 ( .A(G107), .B(n1047), .Z(G9) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U757 ( .A1(G953), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1063) );
NOR2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
INV_X1 U769 ( .A(n1075), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
XNOR2_X1 U771 ( .A(n1078), .B(KEYINPUT44), .ZN(n1076) );
NOR3_X1 U772 ( .A1(n1079), .A2(KEYINPUT13), .A3(n1065), .ZN(n1069) );
AND3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XNOR2_X1 U777 ( .A(KEYINPUT26), .B(n1089), .ZN(n1088) );
NAND2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1080) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U780 ( .A1(KEYINPUT13), .A2(n1094), .ZN(n1092) );
INV_X1 U781 ( .A(n1094), .ZN(n1079) );
AND3_X1 U782 ( .A1(n1082), .A2(n1090), .A3(n1095), .ZN(n1059) );
AND4_X1 U783 ( .A1(n1083), .A2(n1090), .A3(n1096), .A4(n1082), .ZN(n1055) );
NOR3_X1 U784 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1050) );
NOR3_X1 U786 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NAND3_X1 U787 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1101) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U789 ( .A(KEYINPUT7), .B(KEYINPUT39), .Z(n1108) );
XOR2_X1 U790 ( .A(n1109), .B(n1110), .Z(n1107) );
NAND3_X1 U791 ( .A1(KEYINPUT12), .A2(n1111), .A3(n1112), .ZN(n1105) );
INV_X1 U792 ( .A(n1113), .ZN(n1111) );
OR2_X1 U793 ( .A1(n1112), .A2(KEYINPUT12), .ZN(n1104) );
NOR3_X1 U794 ( .A1(n1114), .A2(n1078), .A3(n1087), .ZN(n1099) );
INV_X1 U795 ( .A(n1115), .ZN(n1078) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1114) );
XOR2_X1 U797 ( .A(KEYINPUT33), .B(KEYINPUT21), .Z(n1117) );
XOR2_X1 U798 ( .A(n1118), .B(G469), .Z(n1116) );
XNOR2_X1 U799 ( .A(KEYINPUT47), .B(n1119), .ZN(n1098) );
NAND2_X1 U800 ( .A1(n1120), .A2(n1113), .ZN(n1097) );
NAND2_X1 U801 ( .A1(KEYINPUT12), .A2(n1121), .ZN(n1120) );
XNOR2_X1 U802 ( .A(KEYINPUT8), .B(n1112), .ZN(n1121) );
XOR2_X1 U803 ( .A(n1122), .B(n1123), .Z(G72) );
XOR2_X1 U804 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U805 ( .A1(G953), .A2(n1126), .ZN(n1125) );
NAND2_X1 U806 ( .A1(G900), .A2(G227), .ZN(n1126) );
NAND3_X1 U807 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1124) );
XOR2_X1 U808 ( .A(KEYINPUT56), .B(n1130), .Z(n1129) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
AND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
INV_X1 U813 ( .A(KEYINPUT16), .ZN(n1136) );
XNOR2_X1 U814 ( .A(G125), .B(n1137), .ZN(n1135) );
NAND2_X1 U815 ( .A1(KEYINPUT16), .A2(n1138), .ZN(n1133) );
XOR2_X1 U816 ( .A(n1137), .B(G125), .Z(n1138) );
NAND2_X1 U817 ( .A1(KEYINPUT55), .A2(n1139), .ZN(n1137) );
XOR2_X1 U818 ( .A(n1140), .B(n1141), .Z(n1131) );
XNOR2_X1 U819 ( .A(KEYINPUT14), .B(n1142), .ZN(n1141) );
XNOR2_X1 U820 ( .A(n1143), .B(n1144), .ZN(n1140) );
NAND2_X1 U821 ( .A1(G953), .A2(n1145), .ZN(n1127) );
AND2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(n1122) );
XOR2_X1 U823 ( .A(n1148), .B(n1149), .Z(G69) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1147), .ZN(n1149) );
AND2_X1 U825 ( .A1(G224), .A2(G898), .ZN(n1150) );
NAND2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NAND2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1151) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1156) );
INV_X1 U830 ( .A(KEYINPUT41), .ZN(n1154) );
NAND2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1153) );
NAND2_X1 U832 ( .A1(G953), .A2(n1159), .ZN(n1158) );
XNOR2_X1 U833 ( .A(n1160), .B(n1161), .ZN(n1157) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1160) );
NAND2_X1 U835 ( .A1(n1147), .A2(n1164), .ZN(n1155) );
NOR3_X1 U836 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(G66) );
AND3_X1 U837 ( .A1(KEYINPUT60), .A2(G953), .A3(G952), .ZN(n1167) );
NOR2_X1 U838 ( .A1(KEYINPUT60), .A2(n1168), .ZN(n1166) );
INV_X1 U839 ( .A(n1169), .ZN(n1168) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1165) );
NAND2_X1 U841 ( .A1(n1172), .A2(n1110), .ZN(n1170) );
NOR2_X1 U842 ( .A1(n1169), .A2(n1173), .ZN(G63) );
XOR2_X1 U843 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U844 ( .A(KEYINPUT15), .B(n1176), .ZN(n1174) );
NOR3_X1 U845 ( .A1(n1177), .A2(KEYINPUT51), .A3(n1178), .ZN(n1176) );
NOR2_X1 U846 ( .A1(n1169), .A2(n1179), .ZN(G60) );
NOR2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U848 ( .A(KEYINPUT50), .B(n1182), .Z(n1181) );
NOR2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
AND2_X1 U850 ( .A1(n1184), .A2(n1183), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1172), .A2(G475), .ZN(n1184) );
XOR2_X1 U852 ( .A(G104), .B(n1185), .Z(G6) );
NOR2_X1 U853 ( .A1(n1186), .A2(n1187), .ZN(G57) );
XOR2_X1 U854 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U855 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND4_X1 U856 ( .A1(KEYINPUT18), .A2(G472), .A3(G902), .A4(n1192), .ZN(n1190) );
XNOR2_X1 U857 ( .A(KEYINPUT58), .B(n1052), .ZN(n1192) );
INV_X1 U858 ( .A(n1193), .ZN(n1052) );
XNOR2_X1 U859 ( .A(n1194), .B(n1195), .ZN(n1188) );
NOR2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NOR2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
INV_X1 U862 ( .A(n1200), .ZN(n1199) );
NOR2_X1 U863 ( .A1(KEYINPUT49), .A2(n1201), .ZN(n1198) );
NOR2_X1 U864 ( .A1(KEYINPUT57), .A2(n1202), .ZN(n1201) );
NOR2_X1 U865 ( .A1(G101), .A2(n1203), .ZN(n1196) );
NOR2_X1 U866 ( .A1(n1204), .A2(KEYINPUT57), .ZN(n1203) );
NOR2_X1 U867 ( .A1(KEYINPUT49), .A2(n1200), .ZN(n1204) );
NOR2_X1 U868 ( .A1(G952), .A2(n1205), .ZN(n1186) );
XNOR2_X1 U869 ( .A(G953), .B(KEYINPUT35), .ZN(n1205) );
NOR2_X1 U870 ( .A1(n1169), .A2(n1206), .ZN(G54) );
XOR2_X1 U871 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U872 ( .A(n1209), .B(n1210), .Z(n1208) );
AND2_X1 U873 ( .A1(G469), .A2(n1172), .ZN(n1210) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
XOR2_X1 U875 ( .A(n1213), .B(KEYINPUT9), .Z(n1212) );
NAND2_X1 U876 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
NOR2_X1 U878 ( .A1(n1169), .A2(n1216), .ZN(G51) );
XOR2_X1 U879 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U880 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U881 ( .A(n1221), .B(KEYINPUT29), .Z(n1220) );
NAND2_X1 U882 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U883 ( .A(KEYINPUT3), .B(n1224), .ZN(n1222) );
XOR2_X1 U884 ( .A(n1225), .B(n1226), .Z(n1217) );
NOR2_X1 U885 ( .A1(KEYINPUT40), .A2(n1227), .ZN(n1226) );
NAND3_X1 U886 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1225) );
NAND2_X1 U887 ( .A1(KEYINPUT0), .A2(n1177), .ZN(n1229) );
INV_X1 U888 ( .A(n1172), .ZN(n1177) );
NOR2_X1 U889 ( .A1(n1231), .A2(n1193), .ZN(n1172) );
NAND2_X1 U890 ( .A1(n1232), .A2(n1233), .ZN(n1228) );
INV_X1 U891 ( .A(KEYINPUT0), .ZN(n1233) );
NAND2_X1 U892 ( .A1(n1193), .A2(G902), .ZN(n1232) );
NOR2_X1 U893 ( .A1(n1164), .A2(n1146), .ZN(n1193) );
NAND4_X1 U894 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1146) );
NOR4_X1 U895 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
NOR2_X1 U896 ( .A1(n1242), .A2(n1243), .ZN(n1236) );
NOR3_X1 U897 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
AND2_X1 U898 ( .A1(n1244), .A2(n1247), .ZN(n1242) );
INV_X1 U899 ( .A(KEYINPUT30), .ZN(n1244) );
NAND2_X1 U900 ( .A1(n1248), .A2(n1249), .ZN(n1234) );
NAND2_X1 U901 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U902 ( .A1(n1252), .A2(n1253), .ZN(n1164) );
NOR4_X1 U903 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1185), .ZN(n1253) );
AND3_X1 U904 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1185) );
NOR4_X1 U905 ( .A1(n1047), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1252) );
NOR2_X1 U906 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NOR2_X1 U907 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
NOR2_X1 U908 ( .A1(n1251), .A2(n1267), .ZN(n1265) );
NOR3_X1 U909 ( .A1(n1268), .A2(n1068), .A3(n1251), .ZN(n1261) );
NAND3_X1 U910 ( .A1(n1269), .A2(n1267), .A3(n1075), .ZN(n1268) );
INV_X1 U911 ( .A(KEYINPUT53), .ZN(n1267) );
INV_X1 U912 ( .A(n1270), .ZN(n1260) );
AND3_X1 U913 ( .A1(n1257), .A2(n1258), .A3(n1094), .ZN(n1047) );
NOR2_X1 U914 ( .A1(n1147), .A2(G952), .ZN(n1169) );
XNOR2_X1 U915 ( .A(n1271), .B(n1241), .ZN(G48) );
AND2_X1 U916 ( .A1(n1272), .A2(n1259), .ZN(n1241) );
XOR2_X1 U917 ( .A(G143), .B(n1247), .Z(G45) );
NOR2_X1 U918 ( .A1(n1246), .A2(n1273), .ZN(n1247) );
NAND4_X1 U919 ( .A1(n1274), .A2(n1096), .A3(n1275), .A4(n1276), .ZN(n1246) );
NOR2_X1 U920 ( .A1(n1277), .A2(n1075), .ZN(n1275) );
XNOR2_X1 U921 ( .A(G140), .B(n1235), .ZN(G42) );
NAND4_X1 U922 ( .A1(n1248), .A2(n1259), .A3(n1119), .A4(n1062), .ZN(n1235) );
XNOR2_X1 U923 ( .A(G137), .B(n1278), .ZN(G39) );
NAND4_X1 U924 ( .A1(n1266), .A2(n1082), .A3(n1279), .A4(n1245), .ZN(n1278) );
XNOR2_X1 U925 ( .A(KEYINPUT10), .B(n1086), .ZN(n1279) );
INV_X1 U926 ( .A(n1066), .ZN(n1082) );
XOR2_X1 U927 ( .A(G134), .B(n1240), .Z(G36) );
AND3_X1 U928 ( .A1(n1096), .A2(n1094), .A3(n1248), .ZN(n1240) );
XNOR2_X1 U929 ( .A(G131), .B(n1280), .ZN(G33) );
NAND3_X1 U930 ( .A1(n1248), .A2(n1281), .A3(KEYINPUT25), .ZN(n1280) );
INV_X1 U931 ( .A(n1251), .ZN(n1281) );
NOR3_X1 U932 ( .A1(n1086), .A2(n1273), .A3(n1066), .ZN(n1248) );
NAND2_X1 U933 ( .A1(n1282), .A2(n1115), .ZN(n1066) );
XOR2_X1 U934 ( .A(KEYINPUT42), .B(n1077), .Z(n1282) );
XNOR2_X1 U935 ( .A(n1239), .B(n1283), .ZN(G30) );
NAND2_X1 U936 ( .A1(KEYINPUT19), .A2(G128), .ZN(n1283) );
AND2_X1 U937 ( .A1(n1272), .A2(n1094), .ZN(n1239) );
AND3_X1 U938 ( .A1(n1276), .A2(n1058), .A3(n1284), .ZN(n1272) );
XNOR2_X1 U939 ( .A(G101), .B(n1270), .ZN(G3) );
NAND3_X1 U940 ( .A1(n1096), .A2(n1276), .A3(n1285), .ZN(n1270) );
NOR3_X1 U941 ( .A1(n1075), .A2(n1286), .A3(n1072), .ZN(n1285) );
XOR2_X1 U942 ( .A(G125), .B(n1238), .Z(G27) );
AND4_X1 U943 ( .A1(n1284), .A2(n1259), .A3(n1119), .A4(n1090), .ZN(n1238) );
NOR3_X1 U944 ( .A1(n1257), .A2(n1273), .A3(n1075), .ZN(n1284) );
INV_X1 U945 ( .A(n1245), .ZN(n1273) );
NAND2_X1 U946 ( .A1(n1287), .A2(n1054), .ZN(n1245) );
XOR2_X1 U947 ( .A(KEYINPUT45), .B(n1288), .Z(n1287) );
AND4_X1 U948 ( .A1(n1145), .A2(n1289), .A3(G953), .A4(G902), .ZN(n1288) );
INV_X1 U949 ( .A(G900), .ZN(n1145) );
XNOR2_X1 U950 ( .A(n1290), .B(n1256), .ZN(G24) );
AND4_X1 U951 ( .A1(n1119), .A2(n1291), .A3(n1257), .A4(n1292), .ZN(n1256) );
NOR2_X1 U952 ( .A1(n1264), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U953 ( .A(G119), .B(n1294), .ZN(G21) );
NAND3_X1 U954 ( .A1(n1266), .A2(n1295), .A3(KEYINPUT23), .ZN(n1294) );
INV_X1 U955 ( .A(n1250), .ZN(n1266) );
NAND2_X1 U956 ( .A1(n1095), .A2(n1058), .ZN(n1250) );
XOR2_X1 U957 ( .A(G116), .B(n1255), .Z(G18) );
AND3_X1 U958 ( .A1(n1295), .A2(n1094), .A3(n1096), .ZN(n1255) );
XNOR2_X1 U959 ( .A(n1296), .B(n1297), .ZN(G15) );
NOR2_X1 U960 ( .A1(n1264), .A2(n1251), .ZN(n1297) );
NAND2_X1 U961 ( .A1(n1259), .A2(n1096), .ZN(n1251) );
NOR2_X1 U962 ( .A1(n1062), .A2(n1119), .ZN(n1096) );
INV_X1 U963 ( .A(n1058), .ZN(n1119) );
INV_X1 U964 ( .A(n1093), .ZN(n1259) );
NAND2_X1 U965 ( .A1(n1298), .A2(n1274), .ZN(n1093) );
XNOR2_X1 U966 ( .A(KEYINPUT22), .B(n1291), .ZN(n1298) );
INV_X1 U967 ( .A(n1295), .ZN(n1264) );
NOR3_X1 U968 ( .A1(n1068), .A2(n1286), .A3(n1075), .ZN(n1295) );
INV_X1 U969 ( .A(n1090), .ZN(n1068) );
NAND2_X1 U970 ( .A1(n1299), .A2(n1300), .ZN(n1090) );
OR2_X1 U971 ( .A1(n1086), .A2(KEYINPUT26), .ZN(n1300) );
NAND3_X1 U972 ( .A1(n1089), .A2(n1301), .A3(KEYINPUT26), .ZN(n1299) );
XOR2_X1 U973 ( .A(G110), .B(n1254), .Z(G12) );
AND2_X1 U974 ( .A1(n1095), .A2(n1258), .ZN(n1254) );
NOR4_X1 U975 ( .A1(n1086), .A2(n1075), .A3(n1058), .A4(n1286), .ZN(n1258) );
INV_X1 U976 ( .A(n1269), .ZN(n1286) );
NAND2_X1 U977 ( .A1(n1054), .A2(n1302), .ZN(n1269) );
NAND4_X1 U978 ( .A1(G902), .A2(G953), .A3(n1289), .A4(n1159), .ZN(n1302) );
INV_X1 U979 ( .A(G898), .ZN(n1159) );
NAND3_X1 U980 ( .A1(n1289), .A2(n1147), .A3(G952), .ZN(n1054) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n1289) );
XNOR2_X1 U982 ( .A(n1303), .B(G472), .ZN(n1058) );
NAND2_X1 U983 ( .A1(n1304), .A2(n1231), .ZN(n1303) );
XOR2_X1 U984 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U985 ( .A(G101), .B(n1307), .ZN(n1306) );
NAND2_X1 U986 ( .A1(KEYINPUT54), .A2(n1195), .ZN(n1307) );
NAND2_X1 U987 ( .A1(n1308), .A2(n1309), .ZN(n1195) );
NAND2_X1 U988 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U989 ( .A1(G116), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U990 ( .A(G113), .B(G119), .ZN(n1310) );
NAND2_X1 U991 ( .A1(n1313), .A2(n1312), .ZN(n1308) );
INV_X1 U992 ( .A(KEYINPUT48), .ZN(n1312) );
NAND2_X1 U993 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND3_X1 U994 ( .A1(G113), .A2(n1316), .A3(G116), .ZN(n1315) );
XNOR2_X1 U995 ( .A(n1191), .B(n1200), .ZN(n1305) );
NAND2_X1 U996 ( .A1(G210), .A2(n1317), .ZN(n1200) );
XOR2_X1 U997 ( .A(n1318), .B(n1319), .Z(n1191) );
NAND2_X1 U998 ( .A1(n1077), .A2(n1115), .ZN(n1075) );
NAND2_X1 U999 ( .A1(G214), .A2(n1320), .ZN(n1115) );
XNOR2_X1 U1000 ( .A(n1113), .B(n1230), .ZN(n1077) );
INV_X1 U1001 ( .A(n1112), .ZN(n1230) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1320), .ZN(n1112) );
NAND2_X1 U1003 ( .A1(n1321), .A2(n1231), .ZN(n1320) );
INV_X1 U1004 ( .A(G237), .ZN(n1321) );
NAND2_X1 U1005 ( .A1(n1322), .A2(n1323), .ZN(n1113) );
XOR2_X1 U1006 ( .A(n1227), .B(n1324), .Z(n1323) );
XNOR2_X1 U1007 ( .A(n1325), .B(n1221), .ZN(n1324) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1147), .ZN(n1221) );
NAND2_X1 U1009 ( .A1(n1326), .A2(n1224), .ZN(n1325) );
OR2_X1 U1010 ( .A1(n1327), .A2(G125), .ZN(n1224) );
XNOR2_X1 U1011 ( .A(KEYINPUT31), .B(n1223), .ZN(n1326) );
NAND2_X1 U1012 ( .A1(G125), .A2(n1327), .ZN(n1223) );
XOR2_X1 U1013 ( .A(G128), .B(n1319), .Z(n1327) );
NOR2_X1 U1014 ( .A1(KEYINPUT37), .A2(n1144), .ZN(n1319) );
XOR2_X1 U1015 ( .A(n1328), .B(n1163), .Z(n1227) );
XNOR2_X1 U1016 ( .A(n1290), .B(n1329), .ZN(n1163) );
NAND3_X1 U1017 ( .A1(n1330), .A2(n1331), .A3(KEYINPUT2), .ZN(n1328) );
NAND2_X1 U1018 ( .A1(n1162), .A2(n1161), .ZN(n1331) );
XOR2_X1 U1019 ( .A(KEYINPUT34), .B(n1332), .Z(n1330) );
NOR2_X1 U1020 ( .A1(n1162), .A2(n1161), .ZN(n1332) );
XNOR2_X1 U1021 ( .A(n1333), .B(n1334), .ZN(n1161) );
NOR2_X1 U1022 ( .A1(G104), .A2(KEYINPUT6), .ZN(n1334) );
AND3_X1 U1023 ( .A1(n1335), .A2(n1336), .A3(n1314), .ZN(n1162) );
NAND3_X1 U1024 ( .A1(G116), .A2(n1296), .A3(G119), .ZN(n1314) );
NAND2_X1 U1025 ( .A1(n1337), .A2(n1316), .ZN(n1336) );
XNOR2_X1 U1026 ( .A(G113), .B(G116), .ZN(n1337) );
OR3_X1 U1027 ( .A1(n1296), .A2(G116), .A3(n1316), .ZN(n1335) );
INV_X1 U1028 ( .A(G119), .ZN(n1316) );
XNOR2_X1 U1029 ( .A(KEYINPUT63), .B(n1231), .ZN(n1322) );
INV_X1 U1030 ( .A(n1276), .ZN(n1086) );
NOR2_X1 U1031 ( .A1(n1089), .A2(n1087), .ZN(n1276) );
INV_X1 U1032 ( .A(n1301), .ZN(n1087) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1338), .ZN(n1301) );
XOR2_X1 U1034 ( .A(n1339), .B(n1340), .Z(n1089) );
NOR2_X1 U1035 ( .A1(G469), .A2(KEYINPUT46), .ZN(n1340) );
XOR2_X1 U1036 ( .A(n1118), .B(KEYINPUT20), .Z(n1339) );
NAND2_X1 U1037 ( .A1(n1341), .A2(n1231), .ZN(n1118) );
XOR2_X1 U1038 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1039 ( .A(KEYINPUT17), .B(n1215), .ZN(n1343) );
NAND2_X1 U1040 ( .A1(n1344), .A2(G227), .ZN(n1215) );
XNOR2_X1 U1041 ( .A(G953), .B(KEYINPUT61), .ZN(n1344) );
XNOR2_X1 U1042 ( .A(n1207), .B(n1214), .ZN(n1342) );
XOR2_X1 U1043 ( .A(n1139), .B(n1329), .Z(n1214) );
INV_X1 U1044 ( .A(G140), .ZN(n1139) );
XOR2_X1 U1045 ( .A(n1345), .B(n1346), .Z(n1207) );
XOR2_X1 U1046 ( .A(n1144), .B(n1333), .Z(n1346) );
XNOR2_X1 U1047 ( .A(G107), .B(n1202), .ZN(n1333) );
INV_X1 U1048 ( .A(G101), .ZN(n1202) );
XOR2_X1 U1049 ( .A(G143), .B(G146), .Z(n1144) );
XOR2_X1 U1050 ( .A(n1318), .B(G104), .Z(n1345) );
XNOR2_X1 U1051 ( .A(n1347), .B(n1348), .ZN(n1318) );
INV_X1 U1052 ( .A(n1143), .ZN(n1348) );
XOR2_X1 U1053 ( .A(G137), .B(n1349), .Z(n1143) );
NAND2_X1 U1054 ( .A1(KEYINPUT24), .A2(n1142), .ZN(n1347) );
INV_X1 U1055 ( .A(G131), .ZN(n1142) );
NOR2_X1 U1056 ( .A1(n1072), .A2(n1257), .ZN(n1095) );
INV_X1 U1057 ( .A(n1062), .ZN(n1257) );
XNOR2_X1 U1058 ( .A(n1350), .B(n1351), .ZN(n1062) );
XOR2_X1 U1059 ( .A(KEYINPUT27), .B(n1110), .Z(n1351) );
AND2_X1 U1060 ( .A1(G217), .A2(n1338), .ZN(n1110) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1231), .ZN(n1338) );
NAND2_X1 U1062 ( .A1(KEYINPUT59), .A2(n1109), .ZN(n1350) );
NAND2_X1 U1063 ( .A1(n1171), .A2(n1231), .ZN(n1109) );
XOR2_X1 U1064 ( .A(n1352), .B(n1353), .Z(n1171) );
AND2_X1 U1065 ( .A1(n1354), .A2(G221), .ZN(n1353) );
XOR2_X1 U1066 ( .A(n1355), .B(G137), .Z(n1352) );
NAND2_X1 U1067 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1068 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1069 ( .A(KEYINPUT5), .B(n1360), .Z(n1356) );
NOR2_X1 U1070 ( .A1(n1359), .A2(n1358), .ZN(n1360) );
XNOR2_X1 U1071 ( .A(n1361), .B(n1329), .ZN(n1358) );
XOR2_X1 U1072 ( .A(G110), .B(KEYINPUT32), .Z(n1329) );
NAND2_X1 U1073 ( .A1(n1362), .A2(KEYINPUT11), .ZN(n1361) );
XNOR2_X1 U1074 ( .A(G128), .B(G119), .ZN(n1362) );
NAND2_X1 U1075 ( .A1(n1363), .A2(n1364), .ZN(n1359) );
NAND2_X1 U1076 ( .A1(n1365), .A2(n1271), .ZN(n1364) );
XOR2_X1 U1077 ( .A(KEYINPUT43), .B(n1366), .Z(n1363) );
NOR2_X1 U1078 ( .A1(n1365), .A2(n1271), .ZN(n1366) );
XNOR2_X1 U1079 ( .A(G140), .B(G125), .ZN(n1365) );
INV_X1 U1080 ( .A(n1083), .ZN(n1072) );
NAND2_X1 U1081 ( .A1(n1367), .A2(n1368), .ZN(n1083) );
OR3_X1 U1082 ( .A1(n1274), .A2(n1291), .A3(KEYINPUT22), .ZN(n1368) );
NAND2_X1 U1083 ( .A1(KEYINPUT22), .A2(n1094), .ZN(n1367) );
NOR2_X1 U1084 ( .A1(n1277), .A2(n1274), .ZN(n1094) );
INV_X1 U1085 ( .A(n1293), .ZN(n1274) );
XNOR2_X1 U1086 ( .A(n1369), .B(n1102), .ZN(n1293) );
XNOR2_X1 U1087 ( .A(n1370), .B(G475), .ZN(n1102) );
NAND2_X1 U1088 ( .A1(n1183), .A2(n1231), .ZN(n1370) );
XNOR2_X1 U1089 ( .A(n1371), .B(n1372), .ZN(n1183) );
XOR2_X1 U1090 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1091 ( .A(n1296), .B(G104), .ZN(n1374) );
INV_X1 U1092 ( .A(G113), .ZN(n1296) );
XNOR2_X1 U1093 ( .A(n1271), .B(G143), .ZN(n1373) );
INV_X1 U1094 ( .A(G146), .ZN(n1271) );
XOR2_X1 U1095 ( .A(n1375), .B(n1376), .Z(n1371) );
XOR2_X1 U1096 ( .A(n1377), .B(n1378), .Z(n1376) );
AND2_X1 U1097 ( .A1(n1317), .A2(G214), .ZN(n1378) );
NOR2_X1 U1098 ( .A1(G953), .A2(G237), .ZN(n1317) );
NOR2_X1 U1099 ( .A1(KEYINPUT38), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1100 ( .A(G125), .B(n1380), .Z(n1379) );
NOR2_X1 U1101 ( .A1(G140), .A2(KEYINPUT4), .ZN(n1380) );
XOR2_X1 U1102 ( .A(n1381), .B(n1382), .Z(n1375) );
NOR2_X1 U1103 ( .A1(G131), .A2(KEYINPUT52), .ZN(n1382) );
NAND2_X1 U1104 ( .A1(KEYINPUT1), .A2(n1290), .ZN(n1381) );
XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(KEYINPUT28), .ZN(n1369) );
INV_X1 U1106 ( .A(n1291), .ZN(n1277) );
XOR2_X1 U1107 ( .A(n1103), .B(KEYINPUT36), .Z(n1291) );
XOR2_X1 U1108 ( .A(n1383), .B(n1178), .Z(n1103) );
INV_X1 U1109 ( .A(G478), .ZN(n1178) );
NAND2_X1 U1110 ( .A1(n1175), .A2(n1231), .ZN(n1383) );
INV_X1 U1111 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1112 ( .A(n1384), .B(n1385), .ZN(n1175) );
XOR2_X1 U1113 ( .A(G116), .B(n1386), .Z(n1385) );
XNOR2_X1 U1114 ( .A(G143), .B(n1290), .ZN(n1386) );
INV_X1 U1115 ( .A(G122), .ZN(n1290) );
XOR2_X1 U1116 ( .A(n1387), .B(n1349), .Z(n1384) );
XOR2_X1 U1117 ( .A(G134), .B(G128), .Z(n1349) );
XOR2_X1 U1118 ( .A(n1388), .B(G107), .Z(n1387) );
NAND2_X1 U1119 ( .A1(G217), .A2(n1354), .ZN(n1388) );
AND2_X1 U1120 ( .A1(G234), .A2(n1147), .ZN(n1354) );
INV_X1 U1121 ( .A(G953), .ZN(n1147) );
endmodule


