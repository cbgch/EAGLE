//Key = 0100010010001100010010010101010001010100010111000101100101010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343;

XOR2_X1 U716 ( .A(n1005), .B(n1006), .Z(G9) );
NAND2_X1 U717 ( .A1(KEYINPUT1), .A2(G107), .ZN(n1006) );
NOR2_X1 U718 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U719 ( .A1(n1009), .A2(n1010), .A3(G953), .A4(n1011), .ZN(n1008) );
NOR2_X1 U720 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U721 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U722 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U723 ( .A(n1018), .ZN(n1017) );
NOR2_X1 U724 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NOR2_X1 U725 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U726 ( .A1(n1023), .A2(n1024), .ZN(n1019) );
NOR2_X1 U727 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
AND2_X1 U728 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U729 ( .A1(n1029), .A2(n1030), .ZN(n1025) );
NOR3_X1 U730 ( .A1(n1022), .A2(n1024), .A3(n1031), .ZN(n1014) );
NAND3_X1 U731 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1009) );
XOR2_X1 U732 ( .A(n1035), .B(KEYINPUT35), .Z(n1034) );
NAND2_X1 U733 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U734 ( .A1(n1018), .A2(n1038), .A3(n1039), .ZN(n1037) );
NAND2_X1 U735 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND3_X1 U736 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NAND2_X1 U737 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
NAND2_X1 U738 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U739 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND3_X1 U740 ( .A1(n1052), .A2(n1028), .A3(n1053), .ZN(n1047) );
NAND4_X1 U741 ( .A1(n1039), .A2(n1043), .A3(n1045), .A4(n1054), .ZN(n1036) );
INV_X1 U742 ( .A(n1022), .ZN(n1043) );
NAND2_X1 U743 ( .A1(n1051), .A2(n1028), .ZN(n1022) );
INV_X1 U744 ( .A(n1013), .ZN(n1039) );
NOR3_X1 U745 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U746 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1011) );
NOR4_X1 U747 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
XOR2_X1 U748 ( .A(n1063), .B(n1064), .Z(n1062) );
XOR2_X1 U749 ( .A(n1065), .B(n1066), .Z(n1061) );
XNOR2_X1 U750 ( .A(KEYINPUT51), .B(n1067), .ZN(n1066) );
NOR2_X1 U751 ( .A1(n1068), .A2(KEYINPUT32), .ZN(n1065) );
XOR2_X1 U752 ( .A(n1069), .B(KEYINPUT59), .Z(n1060) );
XOR2_X1 U753 ( .A(n1070), .B(KEYINPUT17), .Z(n1059) );
NOR3_X1 U754 ( .A1(n1053), .A2(n1071), .A3(n1044), .ZN(n1057) );
XOR2_X1 U755 ( .A(n1072), .B(n1073), .Z(n1056) );
XOR2_X1 U756 ( .A(n1074), .B(KEYINPUT28), .Z(n1073) );
NAND2_X1 U757 ( .A1(KEYINPUT5), .A2(n1075), .ZN(n1072) );
XOR2_X1 U758 ( .A(n1076), .B(n1077), .Z(n1055) );
NAND2_X1 U759 ( .A1(KEYINPUT44), .A2(n1078), .ZN(n1077) );
XOR2_X1 U760 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U761 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U762 ( .A(n1083), .ZN(n1082) );
NOR2_X1 U763 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U764 ( .A1(n1086), .A2(n1087), .ZN(n1079) );
NAND2_X1 U765 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U766 ( .A(n1032), .B(n1090), .Z(n1088) );
OR3_X1 U767 ( .A1(n1085), .A2(n1090), .A3(n1089), .ZN(n1086) );
XNOR2_X1 U768 ( .A(n1091), .B(n1092), .ZN(n1090) );
XOR2_X1 U769 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U770 ( .A1(G131), .A2(KEYINPUT19), .ZN(n1093) );
XOR2_X1 U771 ( .A(n1095), .B(n1096), .Z(n1091) );
XNOR2_X1 U772 ( .A(n1097), .B(n1098), .ZN(n1096) );
NOR2_X1 U773 ( .A1(KEYINPUT60), .A2(n1099), .ZN(n1098) );
XNOR2_X1 U774 ( .A(G125), .B(KEYINPUT55), .ZN(n1099) );
NAND2_X1 U775 ( .A1(KEYINPUT12), .A2(n1100), .ZN(n1095) );
NAND3_X1 U776 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(G69) );
NAND2_X1 U777 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U778 ( .A1(KEYINPUT42), .A2(n1106), .ZN(n1102) );
NAND2_X1 U779 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U780 ( .A(KEYINPUT26), .B(n1105), .ZN(n1108) );
INV_X1 U781 ( .A(n1104), .ZN(n1107) );
NAND2_X1 U782 ( .A1(n1109), .A2(n1110), .ZN(n1101) );
INV_X1 U783 ( .A(KEYINPUT42), .ZN(n1110) );
NAND2_X1 U784 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
OR3_X1 U785 ( .A1(n1105), .A2(n1104), .A3(KEYINPUT26), .ZN(n1112) );
XNOR2_X1 U786 ( .A(n1113), .B(n1114), .ZN(n1104) );
NOR2_X1 U787 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U788 ( .A1(G898), .A2(n1089), .ZN(n1115) );
NAND3_X1 U789 ( .A1(n1117), .A2(n1089), .A3(KEYINPUT49), .ZN(n1113) );
NAND2_X1 U790 ( .A1(KEYINPUT26), .A2(n1105), .ZN(n1111) );
NAND2_X1 U791 ( .A1(n1083), .A2(n1118), .ZN(n1105) );
NAND2_X1 U792 ( .A1(G224), .A2(n1119), .ZN(n1118) );
XNOR2_X1 U793 ( .A(KEYINPUT34), .B(n1120), .ZN(n1119) );
XOR2_X1 U794 ( .A(G953), .B(KEYINPUT53), .Z(n1083) );
NOR3_X1 U795 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(G66) );
NOR2_X1 U796 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U797 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR3_X1 U798 ( .A1(n1128), .A2(KEYINPUT4), .A3(n1129), .ZN(n1127) );
INV_X1 U799 ( .A(KEYINPUT52), .ZN(n1128) );
NOR2_X1 U800 ( .A1(KEYINPUT52), .A2(n1130), .ZN(n1126) );
NOR2_X1 U801 ( .A1(n1131), .A2(n1132), .ZN(n1122) );
INV_X1 U802 ( .A(n1124), .ZN(n1132) );
NOR2_X1 U803 ( .A1(KEYINPUT4), .A2(n1129), .ZN(n1131) );
INV_X1 U804 ( .A(n1130), .ZN(n1129) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1064), .ZN(n1130) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1134), .ZN(G63) );
XOR2_X1 U807 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U808 ( .A1(KEYINPUT0), .A2(n1137), .ZN(n1136) );
NAND2_X1 U809 ( .A1(n1138), .A2(G478), .ZN(n1135) );
NOR2_X1 U810 ( .A1(n1121), .A2(n1139), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1140), .B(n1141), .ZN(n1139) );
AND2_X1 U812 ( .A1(G475), .A2(n1138), .ZN(n1141) );
INV_X1 U813 ( .A(n1133), .ZN(n1138) );
XNOR2_X1 U814 ( .A(G104), .B(n1142), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1143), .A2(n1144), .ZN(G57) );
XOR2_X1 U816 ( .A(n1145), .B(KEYINPUT46), .Z(n1144) );
NAND2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U818 ( .A1(n1121), .A2(n1148), .ZN(n1147) );
OR3_X1 U819 ( .A1(G952), .A2(G953), .A3(n1148), .ZN(n1146) );
INV_X1 U820 ( .A(KEYINPUT31), .ZN(n1148) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1143) );
XOR2_X1 U822 ( .A(n1151), .B(n1152), .Z(n1149) );
NOR2_X1 U823 ( .A1(n1075), .A2(n1133), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1153), .A2(KEYINPUT29), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U826 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
NAND2_X1 U827 ( .A1(KEYINPUT13), .A2(n1159), .ZN(n1157) );
OR2_X1 U828 ( .A1(n1160), .A2(KEYINPUT13), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1121), .A2(n1161), .ZN(G54) );
XOR2_X1 U830 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U831 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U832 ( .A1(n1078), .A2(n1133), .ZN(n1164) );
XNOR2_X1 U833 ( .A(G140), .B(G110), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1121), .A2(n1166), .ZN(G51) );
XOR2_X1 U835 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U836 ( .A1(n1067), .A2(n1133), .ZN(n1168) );
NAND2_X1 U837 ( .A1(G902), .A2(n1169), .ZN(n1133) );
NAND2_X1 U838 ( .A1(n1032), .A2(n1033), .ZN(n1169) );
INV_X1 U839 ( .A(n1117), .ZN(n1033) );
NAND4_X1 U840 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1117) );
AND4_X1 U841 ( .A1(n1005), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1173) );
NAND3_X1 U842 ( .A1(n1054), .A2(n1177), .A3(n1028), .ZN(n1005) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U845 ( .A(KEYINPUT43), .B(n1182), .Z(n1181) );
INV_X1 U846 ( .A(n1142), .ZN(n1178) );
NAND3_X1 U847 ( .A1(n1028), .A2(n1177), .A3(n1183), .ZN(n1142) );
NAND2_X1 U848 ( .A1(n1184), .A2(n1185), .ZN(n1171) );
NAND2_X1 U849 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND4_X1 U850 ( .A1(n1028), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
NOR3_X1 U851 ( .A1(n1191), .A2(KEYINPUT63), .A3(n1051), .ZN(n1190) );
XNOR2_X1 U852 ( .A(n1192), .B(KEYINPUT14), .ZN(n1186) );
NAND2_X1 U853 ( .A1(KEYINPUT63), .A2(n1193), .ZN(n1170) );
AND4_X1 U854 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1032) );
AND4_X1 U855 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NOR3_X1 U856 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1196) );
NOR2_X1 U857 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
INV_X1 U858 ( .A(KEYINPUT62), .ZN(n1205) );
NOR3_X1 U859 ( .A1(KEYINPUT62), .A2(n1207), .A3(n1021), .ZN(n1203) );
NOR3_X1 U860 ( .A1(n1031), .A2(n1029), .A3(n1208), .ZN(n1202) );
INV_X1 U861 ( .A(n1183), .ZN(n1031) );
NAND2_X1 U862 ( .A1(KEYINPUT23), .A2(n1209), .ZN(n1167) );
XOR2_X1 U863 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U864 ( .A1(KEYINPUT3), .A2(n1212), .ZN(n1210) );
XNOR2_X1 U865 ( .A(n1213), .B(n1214), .ZN(n1212) );
NOR2_X1 U866 ( .A1(G125), .A2(KEYINPUT56), .ZN(n1213) );
NOR2_X1 U867 ( .A1(n1089), .A2(G952), .ZN(n1121) );
XNOR2_X1 U868 ( .A(G146), .B(n1194), .ZN(G48) );
NAND4_X1 U869 ( .A1(n1183), .A2(n1215), .A3(n1027), .A4(n1216), .ZN(n1194) );
XNOR2_X1 U870 ( .A(G143), .B(n1217), .ZN(G45) );
NOR2_X1 U871 ( .A1(n1218), .A2(KEYINPUT40), .ZN(n1217) );
INV_X1 U872 ( .A(n1199), .ZN(n1218) );
NAND4_X1 U873 ( .A1(n1216), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1199) );
NOR3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(n1021), .ZN(n1221) );
XNOR2_X1 U875 ( .A(G140), .B(n1195), .ZN(G42) );
NAND2_X1 U876 ( .A1(n1224), .A2(n1225), .ZN(n1195) );
XNOR2_X1 U877 ( .A(G137), .B(n1198), .ZN(G39) );
NAND4_X1 U878 ( .A1(n1018), .A2(n1225), .A3(n1050), .A4(n1226), .ZN(n1198) );
XNOR2_X1 U879 ( .A(G134), .B(n1201), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1054), .A2(n1220), .A3(n1225), .ZN(n1201) );
INV_X1 U881 ( .A(n1208), .ZN(n1225) );
NAND3_X1 U882 ( .A1(n1027), .A2(n1216), .A3(n1045), .ZN(n1208) );
XNOR2_X1 U883 ( .A(G131), .B(n1227), .ZN(G33) );
NAND4_X1 U884 ( .A1(n1228), .A2(n1183), .A3(n1229), .A4(n1045), .ZN(n1227) );
INV_X1 U885 ( .A(n1024), .ZN(n1045) );
NAND2_X1 U886 ( .A1(n1042), .A2(n1230), .ZN(n1024) );
NOR2_X1 U887 ( .A1(n1029), .A2(n1223), .ZN(n1229) );
INV_X1 U888 ( .A(n1027), .ZN(n1223) );
INV_X1 U889 ( .A(n1220), .ZN(n1029) );
XOR2_X1 U890 ( .A(n1216), .B(KEYINPUT11), .Z(n1228) );
XOR2_X1 U891 ( .A(n1200), .B(n1231), .Z(G30) );
NAND2_X1 U892 ( .A1(KEYINPUT8), .A2(G128), .ZN(n1231) );
NAND4_X1 U893 ( .A1(n1215), .A2(n1054), .A3(n1232), .A4(n1216), .ZN(n1200) );
XNOR2_X1 U894 ( .A(G101), .B(n1176), .ZN(G3) );
NAND3_X1 U895 ( .A1(n1177), .A2(n1220), .A3(n1018), .ZN(n1176) );
NOR3_X1 U896 ( .A1(n1233), .A2(n1234), .A3(n1180), .ZN(n1177) );
INV_X1 U897 ( .A(n1235), .ZN(n1180) );
XOR2_X1 U898 ( .A(n1206), .B(n1236), .Z(G27) );
XOR2_X1 U899 ( .A(KEYINPUT25), .B(G125), .Z(n1236) );
NAND2_X1 U900 ( .A1(n1207), .A2(n1184), .ZN(n1206) );
AND3_X1 U901 ( .A1(n1224), .A2(n1216), .A3(n1051), .ZN(n1207) );
INV_X1 U902 ( .A(n1030), .ZN(n1051) );
NAND2_X1 U903 ( .A1(n1013), .A2(n1237), .ZN(n1216) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1238), .A4(n1085), .ZN(n1237) );
INV_X1 U905 ( .A(G900), .ZN(n1085) );
AND3_X1 U906 ( .A1(n1049), .A2(n1050), .A3(n1183), .ZN(n1224) );
XOR2_X1 U907 ( .A(G122), .B(n1193), .Z(G24) );
AND4_X1 U908 ( .A1(n1189), .A2(n1239), .A3(n1240), .A4(n1028), .ZN(n1193) );
NOR2_X1 U909 ( .A1(n1191), .A2(n1021), .ZN(n1240) );
INV_X1 U910 ( .A(n1184), .ZN(n1021) );
XNOR2_X1 U911 ( .A(G119), .B(n1175), .ZN(G21) );
NAND3_X1 U912 ( .A1(n1215), .A2(n1018), .A3(n1239), .ZN(n1175) );
AND3_X1 U913 ( .A1(n1050), .A2(n1226), .A3(n1184), .ZN(n1215) );
XNOR2_X1 U914 ( .A(G116), .B(n1241), .ZN(G18) );
NAND2_X1 U915 ( .A1(n1192), .A2(n1184), .ZN(n1241) );
AND3_X1 U916 ( .A1(n1054), .A2(n1220), .A3(n1239), .ZN(n1192) );
NOR2_X1 U917 ( .A1(n1189), .A2(n1191), .ZN(n1054) );
INV_X1 U918 ( .A(n1219), .ZN(n1191) );
XNOR2_X1 U919 ( .A(G113), .B(n1174), .ZN(G15) );
NAND4_X1 U920 ( .A1(n1239), .A2(n1183), .A3(n1220), .A4(n1235), .ZN(n1174) );
NAND2_X1 U921 ( .A1(n1242), .A2(n1243), .ZN(n1220) );
OR3_X1 U922 ( .A1(n1244), .A2(n1049), .A3(KEYINPUT47), .ZN(n1243) );
NAND2_X1 U923 ( .A1(KEYINPUT47), .A2(n1028), .ZN(n1242) );
NOR2_X1 U924 ( .A1(n1226), .A2(n1244), .ZN(n1028) );
NOR2_X1 U925 ( .A1(n1222), .A2(n1219), .ZN(n1183) );
NOR2_X1 U926 ( .A1(n1030), .A2(n1234), .ZN(n1239) );
NAND2_X1 U927 ( .A1(n1052), .A2(n1245), .ZN(n1030) );
XNOR2_X1 U928 ( .A(G110), .B(n1246), .ZN(G12) );
NAND3_X1 U929 ( .A1(n1182), .A2(n1235), .A3(KEYINPUT61), .ZN(n1246) );
XOR2_X1 U930 ( .A(n1184), .B(KEYINPUT6), .Z(n1235) );
NOR2_X1 U931 ( .A1(n1042), .A2(n1044), .ZN(n1184) );
INV_X1 U932 ( .A(n1230), .ZN(n1044) );
NAND2_X1 U933 ( .A1(G214), .A2(n1247), .ZN(n1230) );
XOR2_X1 U934 ( .A(n1068), .B(n1067), .Z(n1042) );
NAND2_X1 U935 ( .A1(G210), .A2(n1247), .ZN(n1067) );
NAND2_X1 U936 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U937 ( .A(G237), .ZN(n1249) );
AND2_X1 U938 ( .A1(n1250), .A2(n1248), .ZN(n1068) );
XNOR2_X1 U939 ( .A(n1211), .B(n1251), .ZN(n1250) );
XNOR2_X1 U940 ( .A(G125), .B(n1252), .ZN(n1251) );
NAND2_X1 U941 ( .A1(KEYINPUT57), .A2(n1214), .ZN(n1252) );
XOR2_X1 U942 ( .A(n1116), .B(n1253), .Z(n1211) );
AND2_X1 U943 ( .A1(n1089), .A2(G224), .ZN(n1253) );
XNOR2_X1 U944 ( .A(n1254), .B(n1255), .ZN(n1116) );
XOR2_X1 U945 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U946 ( .A(n1258), .B(n1259), .Z(n1254) );
XOR2_X1 U947 ( .A(KEYINPUT39), .B(G110), .Z(n1259) );
NAND2_X1 U948 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NAND2_X1 U949 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
INV_X1 U950 ( .A(G113), .ZN(n1263) );
XOR2_X1 U951 ( .A(KEYINPUT41), .B(n1264), .Z(n1260) );
NOR2_X1 U952 ( .A1(n1262), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U953 ( .A(G113), .B(KEYINPUT2), .ZN(n1265) );
AND4_X1 U954 ( .A1(n1049), .A2(n1018), .A3(n1266), .A4(n1050), .ZN(n1182) );
XNOR2_X1 U955 ( .A(n1244), .B(KEYINPUT27), .ZN(n1050) );
XNOR2_X1 U956 ( .A(n1267), .B(n1063), .ZN(n1244) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1248), .ZN(n1063) );
XNOR2_X1 U958 ( .A(n1124), .B(KEYINPUT48), .ZN(n1268) );
XNOR2_X1 U959 ( .A(n1269), .B(n1270), .ZN(n1124) );
XOR2_X1 U960 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U961 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
INV_X1 U962 ( .A(G221), .ZN(n1274) );
XOR2_X1 U963 ( .A(n1275), .B(n1276), .Z(n1269) );
XOR2_X1 U964 ( .A(G146), .B(G137), .Z(n1276) );
NAND2_X1 U965 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
OR2_X1 U966 ( .A1(n1279), .A2(G110), .ZN(n1278) );
XOR2_X1 U967 ( .A(n1280), .B(KEYINPUT36), .Z(n1277) );
NAND2_X1 U968 ( .A1(G110), .A2(n1279), .ZN(n1280) );
XOR2_X1 U969 ( .A(G119), .B(G128), .Z(n1279) );
NAND2_X1 U970 ( .A1(KEYINPUT20), .A2(n1064), .ZN(n1267) );
NAND2_X1 U971 ( .A1(G217), .A2(n1281), .ZN(n1064) );
NOR2_X1 U972 ( .A1(n1234), .A2(n1233), .ZN(n1266) );
INV_X1 U973 ( .A(n1232), .ZN(n1233) );
XOR2_X1 U974 ( .A(n1027), .B(KEYINPUT18), .Z(n1232) );
NOR2_X1 U975 ( .A1(n1052), .A2(n1053), .ZN(n1027) );
INV_X1 U976 ( .A(n1245), .ZN(n1053) );
NAND2_X1 U977 ( .A1(G221), .A2(n1281), .ZN(n1245) );
NAND2_X1 U978 ( .A1(G234), .A2(n1248), .ZN(n1281) );
XNOR2_X1 U979 ( .A(n1076), .B(n1078), .ZN(n1052) );
INV_X1 U980 ( .A(G469), .ZN(n1078) );
NAND2_X1 U981 ( .A1(n1282), .A2(n1248), .ZN(n1076) );
XNOR2_X1 U982 ( .A(n1283), .B(n1165), .ZN(n1282) );
XNOR2_X1 U983 ( .A(n1284), .B(n1285), .ZN(n1165) );
XOR2_X1 U984 ( .A(n1286), .B(n1256), .Z(n1285) );
XOR2_X1 U985 ( .A(G101), .B(n1287), .Z(n1256) );
XNOR2_X1 U986 ( .A(KEYINPUT58), .B(n1288), .ZN(n1287) );
INV_X1 U987 ( .A(G104), .ZN(n1288) );
NOR2_X1 U988 ( .A1(G953), .A2(n1084), .ZN(n1286) );
INV_X1 U989 ( .A(G227), .ZN(n1084) );
NAND2_X1 U990 ( .A1(n1289), .A2(n1290), .ZN(n1284) );
NAND2_X1 U991 ( .A1(G107), .A2(n1291), .ZN(n1290) );
NAND2_X1 U992 ( .A1(n1158), .A2(n1292), .ZN(n1291) );
NAND2_X1 U993 ( .A1(n1293), .A2(n1294), .ZN(n1289) );
XNOR2_X1 U994 ( .A(n1160), .B(n1100), .ZN(n1293) );
NAND2_X1 U995 ( .A1(n1295), .A2(n1296), .ZN(n1283) );
OR4_X1 U996 ( .A1(G110), .A2(G140), .A3(KEYINPUT22), .A4(KEYINPUT38), .ZN(n1296) );
NAND2_X1 U997 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND2_X1 U998 ( .A1(n1299), .A2(n1097), .ZN(n1298) );
NAND2_X1 U999 ( .A1(KEYINPUT38), .A2(G110), .ZN(n1299) );
OR2_X1 U1000 ( .A1(G110), .A2(KEYINPUT22), .ZN(n1297) );
INV_X1 U1001 ( .A(n1188), .ZN(n1234) );
NAND2_X1 U1002 ( .A1(n1013), .A2(n1300), .ZN(n1188) );
NAND4_X1 U1003 ( .A1(G953), .A2(G902), .A3(n1238), .A4(n1120), .ZN(n1300) );
INV_X1 U1004 ( .A(G898), .ZN(n1120) );
NAND3_X1 U1005 ( .A1(n1238), .A2(n1089), .A3(G952), .ZN(n1013) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1238) );
NOR2_X1 U1007 ( .A1(n1219), .A2(n1189), .ZN(n1018) );
INV_X1 U1008 ( .A(n1222), .ZN(n1189) );
XNOR2_X1 U1009 ( .A(n1070), .B(KEYINPUT33), .ZN(n1222) );
XOR2_X1 U1010 ( .A(n1301), .B(n1302), .Z(n1070) );
XOR2_X1 U1011 ( .A(KEYINPUT21), .B(G475), .Z(n1302) );
NAND2_X1 U1012 ( .A1(n1140), .A2(n1248), .ZN(n1301) );
XNOR2_X1 U1013 ( .A(n1303), .B(n1304), .ZN(n1140) );
XOR2_X1 U1014 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1015 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U1016 ( .A1(G113), .A2(KEYINPUT30), .ZN(n1308) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U1018 ( .A(G104), .B(G122), .ZN(n1305) );
XNOR2_X1 U1019 ( .A(n1272), .B(n1310), .ZN(n1303) );
XOR2_X1 U1020 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1021 ( .A1(KEYINPUT50), .A2(n1313), .ZN(n1311) );
INV_X1 U1022 ( .A(G131), .ZN(n1313) );
XOR2_X1 U1023 ( .A(G125), .B(n1314), .Z(n1272) );
XNOR2_X1 U1024 ( .A(KEYINPUT45), .B(n1097), .ZN(n1314) );
INV_X1 U1025 ( .A(G140), .ZN(n1097) );
NAND2_X1 U1026 ( .A1(n1315), .A2(n1069), .ZN(n1219) );
NAND2_X1 U1027 ( .A1(G478), .A2(n1316), .ZN(n1069) );
OR2_X1 U1028 ( .A1(n1137), .A2(G902), .ZN(n1316) );
XNOR2_X1 U1029 ( .A(n1071), .B(KEYINPUT24), .ZN(n1315) );
NOR3_X1 U1030 ( .A1(G478), .A2(G902), .A3(n1137), .ZN(n1071) );
XNOR2_X1 U1031 ( .A(n1317), .B(n1318), .ZN(n1137) );
NOR2_X1 U1032 ( .A1(n1273), .A2(n1319), .ZN(n1318) );
INV_X1 U1033 ( .A(G217), .ZN(n1319) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1089), .ZN(n1273) );
INV_X1 U1035 ( .A(G953), .ZN(n1089) );
NAND3_X1 U1036 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1317) );
NAND2_X1 U1037 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1038 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1039 ( .A(KEYINPUT9), .B(n1327), .Z(n1325) );
NAND3_X1 U1040 ( .A1(n1327), .A2(n1328), .A3(n1326), .ZN(n1321) );
INV_X1 U1041 ( .A(n1323), .ZN(n1328) );
XNOR2_X1 U1042 ( .A(n1329), .B(n1330), .ZN(n1323) );
NOR2_X1 U1043 ( .A1(KEYINPUT7), .A2(G128), .ZN(n1330) );
XNOR2_X1 U1044 ( .A(G134), .B(G143), .ZN(n1329) );
OR2_X1 U1045 ( .A1(n1326), .A2(n1327), .ZN(n1320) );
XNOR2_X1 U1046 ( .A(n1331), .B(n1257), .ZN(n1327) );
XNOR2_X1 U1047 ( .A(G122), .B(n1294), .ZN(n1257) );
INV_X1 U1048 ( .A(G107), .ZN(n1294) );
NAND2_X1 U1049 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1050 ( .A(KEYINPUT16), .B(KEYINPUT15), .ZN(n1332) );
INV_X1 U1051 ( .A(KEYINPUT54), .ZN(n1326) );
INV_X1 U1052 ( .A(n1226), .ZN(n1049) );
XOR2_X1 U1053 ( .A(n1074), .B(n1075), .Z(n1226) );
INV_X1 U1054 ( .A(G472), .ZN(n1075) );
NAND2_X1 U1055 ( .A1(n1334), .A2(n1248), .ZN(n1074) );
INV_X1 U1056 ( .A(G902), .ZN(n1248) );
XOR2_X1 U1057 ( .A(n1335), .B(n1150), .Z(n1334) );
XNOR2_X1 U1058 ( .A(n1336), .B(G101), .ZN(n1150) );
NAND2_X1 U1059 ( .A1(G210), .A2(n1309), .ZN(n1336) );
NOR2_X1 U1060 ( .A1(G953), .A2(G237), .ZN(n1309) );
NOR2_X1 U1061 ( .A1(n1337), .A2(n1338), .ZN(n1335) );
XOR2_X1 U1062 ( .A(KEYINPUT10), .B(n1339), .Z(n1338) );
NOR2_X1 U1063 ( .A1(n1155), .A2(n1340), .ZN(n1339) );
AND2_X1 U1064 ( .A1(n1340), .A2(n1155), .ZN(n1337) );
XNOR2_X1 U1065 ( .A(G113), .B(n1262), .ZN(n1155) );
XOR2_X1 U1066 ( .A(n1333), .B(G119), .Z(n1262) );
INV_X1 U1067 ( .A(G116), .ZN(n1333) );
NAND3_X1 U1068 ( .A1(n1341), .A2(n1342), .A3(n1158), .ZN(n1340) );
OR2_X1 U1069 ( .A1(n1160), .A2(n1214), .ZN(n1158) );
OR2_X1 U1070 ( .A1(n1214), .A2(KEYINPUT37), .ZN(n1342) );
NAND2_X1 U1071 ( .A1(n1159), .A2(KEYINPUT37), .ZN(n1341) );
INV_X1 U1072 ( .A(n1292), .ZN(n1159) );
NAND2_X1 U1073 ( .A1(n1214), .A2(n1160), .ZN(n1292) );
XOR2_X1 U1074 ( .A(G131), .B(n1094), .Z(n1160) );
XNOR2_X1 U1075 ( .A(n1343), .B(G137), .ZN(n1094) );
INV_X1 U1076 ( .A(G134), .ZN(n1343) );
INV_X1 U1077 ( .A(n1100), .ZN(n1214) );
XOR2_X1 U1078 ( .A(G128), .B(n1312), .Z(n1100) );
XOR2_X1 U1079 ( .A(G143), .B(G146), .Z(n1312) );
endmodule


