//Key = 1101111110110011101101001111011000100100110110011110011111111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331;

XOR2_X1 U744 ( .A(n1020), .B(n1021), .Z(G9) );
XOR2_X1 U745 ( .A(KEYINPUT24), .B(G107), .Z(n1021) );
NAND4_X1 U746 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(G75) );
NAND4_X1 U747 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1024) );
NOR4_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
XOR2_X1 U749 ( .A(n1034), .B(n1035), .Z(n1033) );
XOR2_X1 U750 ( .A(KEYINPUT21), .B(n1036), .Z(n1032) );
XOR2_X1 U751 ( .A(KEYINPUT31), .B(n1037), .Z(n1031) );
NOR2_X1 U752 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U753 ( .A(n1040), .B(KEYINPUT57), .Z(n1038) );
XOR2_X1 U754 ( .A(n1041), .B(n1042), .Z(n1030) );
NOR2_X1 U755 ( .A1(n1043), .A2(KEYINPUT33), .ZN(n1041) );
AND3_X1 U756 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1028) );
XNOR2_X1 U757 ( .A(n1047), .B(n1048), .ZN(n1027) );
NOR2_X1 U758 ( .A1(n1049), .A2(KEYINPUT52), .ZN(n1048) );
XOR2_X1 U759 ( .A(KEYINPUT55), .B(n1050), .Z(n1026) );
NAND2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1023) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U762 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND3_X1 U764 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
OR3_X1 U765 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1065), .ZN(n1060) );
INV_X1 U767 ( .A(n1044), .ZN(n1065) );
XOR2_X1 U768 ( .A(KEYINPUT37), .B(n1067), .Z(n1066) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1058) );
NAND4_X1 U770 ( .A1(n1069), .A2(n1044), .A3(n1067), .A4(n1070), .ZN(n1053) );
NOR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR4_X1 U772 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
NOR2_X1 U773 ( .A1(n1055), .A2(n1046), .ZN(n1072) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1069) );
INV_X1 U775 ( .A(n1080), .ZN(n1051) );
XOR2_X1 U776 ( .A(n1081), .B(n1082), .Z(G72) );
NAND2_X1 U777 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U778 ( .A1(G900), .A2(G227), .ZN(n1083) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U781 ( .A1(n1025), .A2(n1088), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U783 ( .A(n1091), .B(KEYINPUT39), .Z(n1089) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1086) );
NAND2_X1 U785 ( .A1(n1094), .A2(G953), .ZN(n1093) );
XOR2_X1 U786 ( .A(n1095), .B(KEYINPUT38), .Z(n1094) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(n1092) );
NAND2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U790 ( .A(n1102), .B(KEYINPUT12), .Z(n1098) );
OR2_X1 U791 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
NAND2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1105), .A2(G137), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
XOR2_X1 U795 ( .A(n1108), .B(KEYINPUT51), .Z(n1106) );
XOR2_X1 U796 ( .A(KEYINPUT50), .B(KEYINPUT32), .Z(n1084) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
OR2_X1 U799 ( .A1(n1025), .A2(G224), .ZN(n1112) );
NAND3_X1 U800 ( .A1(G953), .A2(n1113), .A3(n1114), .ZN(n1109) );
XNOR2_X1 U801 ( .A(n1111), .B(KEYINPUT35), .ZN(n1114) );
XNOR2_X1 U802 ( .A(n1115), .B(n1116), .ZN(n1111) );
NOR2_X1 U803 ( .A1(n1117), .A2(G953), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U805 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1118) );
XOR2_X1 U807 ( .A(n1123), .B(KEYINPUT42), .Z(n1121) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1113) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U811 ( .A1(KEYINPUT3), .A2(n1128), .ZN(n1127) );
INV_X1 U812 ( .A(n1129), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1130), .A2(G217), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1131), .ZN(G63) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U816 ( .A1(n1039), .A2(n1134), .ZN(n1132) );
NOR2_X1 U817 ( .A1(n1124), .A2(n1135), .ZN(G60) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U819 ( .A(KEYINPUT11), .B(n1138), .Z(n1137) );
AND2_X1 U820 ( .A1(G475), .A2(n1130), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(G6) );
NOR2_X1 U822 ( .A1(n1124), .A2(n1141), .ZN(G57) );
XOR2_X1 U823 ( .A(n1142), .B(n1143), .Z(n1141) );
XNOR2_X1 U824 ( .A(n1144), .B(n1145), .ZN(n1143) );
NAND2_X1 U825 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NAND2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U827 ( .A(n1150), .B(n1151), .Z(n1146) );
AND2_X1 U828 ( .A1(G472), .A2(n1130), .ZN(n1151) );
OR2_X1 U829 ( .A1(n1149), .A2(n1148), .ZN(n1150) );
NAND3_X1 U830 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1148) );
NAND2_X1 U831 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR3_X1 U832 ( .A1(n1156), .A2(n1155), .A3(KEYINPUT17), .ZN(n1153) );
NAND2_X1 U833 ( .A1(KEYINPUT4), .A2(n1157), .ZN(n1156) );
NAND2_X1 U834 ( .A1(n1158), .A2(KEYINPUT17), .ZN(n1152) );
INV_X1 U835 ( .A(KEYINPUT44), .ZN(n1149) );
XOR2_X1 U836 ( .A(n1159), .B(KEYINPUT8), .Z(n1142) );
NOR2_X1 U837 ( .A1(n1124), .A2(n1160), .ZN(G54) );
XOR2_X1 U838 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U841 ( .A1(n1034), .A2(n1134), .ZN(n1166) );
INV_X1 U842 ( .A(G469), .ZN(n1034) );
XOR2_X1 U843 ( .A(n1167), .B(n1168), .Z(n1161) );
NOR2_X1 U844 ( .A1(G110), .A2(KEYINPUT13), .ZN(n1168) );
XNOR2_X1 U845 ( .A(G140), .B(n1169), .ZN(n1167) );
NOR2_X1 U846 ( .A1(n1124), .A2(n1170), .ZN(G51) );
XOR2_X1 U847 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U849 ( .A1(n1047), .A2(n1134), .ZN(n1174) );
INV_X1 U850 ( .A(n1130), .ZN(n1134) );
NOR2_X1 U851 ( .A1(n1175), .A2(n1022), .ZN(n1130) );
AND3_X1 U852 ( .A1(n1090), .A2(n1091), .A3(n1117), .ZN(n1022) );
AND4_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1117) );
AND4_X1 U854 ( .A1(n1020), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1179) );
NAND3_X1 U855 ( .A1(n1077), .A2(n1183), .A3(n1067), .ZN(n1020) );
NOR2_X1 U856 ( .A1(n1184), .A2(n1185), .ZN(n1178) );
NOR2_X1 U857 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
INV_X1 U858 ( .A(n1140), .ZN(n1184) );
NAND3_X1 U859 ( .A1(n1067), .A2(n1183), .A3(n1076), .ZN(n1140) );
AND4_X1 U860 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1090) );
NOR4_X1 U861 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
INV_X1 U862 ( .A(n1196), .ZN(n1195) );
NAND3_X1 U863 ( .A1(n1197), .A2(n1198), .A3(KEYINPUT0), .ZN(n1173) );
XNOR2_X1 U864 ( .A(KEYINPUT53), .B(n1199), .ZN(n1197) );
NOR2_X1 U865 ( .A1(n1025), .A2(G952), .ZN(n1124) );
XOR2_X1 U866 ( .A(n1200), .B(n1190), .Z(G48) );
NAND3_X1 U867 ( .A1(n1076), .A2(n1068), .A3(n1201), .ZN(n1190) );
XOR2_X1 U868 ( .A(G143), .B(n1202), .Z(G45) );
NOR2_X1 U869 ( .A1(KEYINPUT63), .A2(n1188), .ZN(n1202) );
NAND4_X1 U870 ( .A1(n1068), .A2(n1075), .A3(n1064), .A4(n1203), .ZN(n1188) );
AND3_X1 U871 ( .A1(n1050), .A2(n1204), .A3(n1205), .ZN(n1203) );
XNOR2_X1 U872 ( .A(G140), .B(n1189), .ZN(G42) );
NAND3_X1 U873 ( .A1(n1076), .A2(n1063), .A3(n1206), .ZN(n1189) );
XOR2_X1 U874 ( .A(n1107), .B(n1196), .Z(G39) );
NAND4_X1 U875 ( .A1(n1062), .A2(n1201), .A3(n1055), .A4(n1044), .ZN(n1196) );
XOR2_X1 U876 ( .A(G134), .B(n1194), .Z(G36) );
AND3_X1 U877 ( .A1(n1064), .A2(n1077), .A3(n1206), .ZN(n1194) );
XOR2_X1 U878 ( .A(G131), .B(n1193), .Z(G33) );
AND3_X1 U879 ( .A1(n1076), .A2(n1064), .A3(n1206), .ZN(n1193) );
AND4_X1 U880 ( .A1(n1062), .A2(n1075), .A3(n1205), .A4(n1044), .ZN(n1206) );
XNOR2_X1 U881 ( .A(G128), .B(n1091), .ZN(G30) );
NAND3_X1 U882 ( .A1(n1077), .A2(n1068), .A3(n1201), .ZN(n1091) );
AND4_X1 U883 ( .A1(n1207), .A2(n1075), .A3(n1205), .A4(n1208), .ZN(n1201) );
XOR2_X1 U884 ( .A(n1159), .B(n1209), .Z(G3) );
NAND2_X1 U885 ( .A1(n1210), .A2(n1068), .ZN(n1209) );
XOR2_X1 U886 ( .A(n1187), .B(KEYINPUT25), .Z(n1210) );
NAND3_X1 U887 ( .A1(n1064), .A2(n1211), .A3(n1212), .ZN(n1187) );
INV_X1 U888 ( .A(n1079), .ZN(n1212) );
NAND2_X1 U889 ( .A1(n1075), .A2(n1055), .ZN(n1079) );
XOR2_X1 U890 ( .A(G125), .B(n1192), .Z(G27) );
AND4_X1 U891 ( .A1(n1068), .A2(n1205), .A3(n1063), .A4(n1213), .ZN(n1192) );
AND2_X1 U892 ( .A1(n1057), .A2(n1076), .ZN(n1213) );
NAND2_X1 U893 ( .A1(n1080), .A2(n1214), .ZN(n1205) );
NAND4_X1 U894 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1095), .ZN(n1214) );
INV_X1 U895 ( .A(G900), .ZN(n1095) );
XNOR2_X1 U896 ( .A(G122), .B(n1176), .ZN(G24) );
NAND4_X1 U897 ( .A1(n1216), .A2(n1067), .A3(n1050), .A4(n1204), .ZN(n1176) );
NOR2_X1 U898 ( .A1(n1208), .A2(n1207), .ZN(n1067) );
XOR2_X1 U899 ( .A(n1177), .B(n1217), .Z(G21) );
XOR2_X1 U900 ( .A(KEYINPUT10), .B(G119), .Z(n1217) );
NAND4_X1 U901 ( .A1(n1207), .A2(n1216), .A3(n1055), .A4(n1208), .ZN(n1177) );
XNOR2_X1 U902 ( .A(n1182), .B(n1218), .ZN(G18) );
NOR2_X1 U903 ( .A1(KEYINPUT45), .A2(n1219), .ZN(n1218) );
NAND3_X1 U904 ( .A1(n1064), .A2(n1077), .A3(n1216), .ZN(n1182) );
XNOR2_X1 U905 ( .A(G113), .B(n1181), .ZN(G15) );
NAND3_X1 U906 ( .A1(n1076), .A2(n1064), .A3(n1216), .ZN(n1181) );
AND3_X1 U907 ( .A1(n1068), .A2(n1211), .A3(n1057), .ZN(n1216) );
NOR2_X1 U908 ( .A1(n1078), .A2(n1074), .ZN(n1057) );
AND2_X1 U909 ( .A1(n1207), .A2(n1220), .ZN(n1064) );
XOR2_X1 U910 ( .A(KEYINPUT22), .B(n1036), .Z(n1220) );
NOR2_X1 U911 ( .A1(n1204), .A2(n1221), .ZN(n1076) );
XOR2_X1 U912 ( .A(n1222), .B(n1180), .Z(G12) );
NAND3_X1 U913 ( .A1(n1183), .A2(n1055), .A3(n1063), .ZN(n1180) );
NOR2_X1 U914 ( .A1(n1207), .A2(n1036), .ZN(n1063) );
INV_X1 U915 ( .A(n1208), .ZN(n1036) );
NAND3_X1 U916 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1208) );
OR2_X1 U917 ( .A1(n1129), .A2(n1226), .ZN(n1225) );
NAND3_X1 U918 ( .A1(n1226), .A2(n1129), .A3(n1175), .ZN(n1224) );
NAND2_X1 U919 ( .A1(n1227), .A2(n1228), .ZN(n1129) );
NAND2_X1 U920 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XOR2_X1 U921 ( .A(KEYINPUT49), .B(n1231), .Z(n1227) );
NOR2_X1 U922 ( .A1(n1229), .A2(n1230), .ZN(n1231) );
XOR2_X1 U923 ( .A(n1232), .B(n1107), .Z(n1230) );
NAND2_X1 U924 ( .A1(G221), .A2(n1233), .ZN(n1232) );
XOR2_X1 U925 ( .A(n1234), .B(n1097), .Z(n1229) );
XOR2_X1 U926 ( .A(n1235), .B(G146), .Z(n1234) );
NAND2_X1 U927 ( .A1(n1236), .A2(KEYINPUT26), .ZN(n1235) );
XOR2_X1 U928 ( .A(n1222), .B(n1237), .Z(n1236) );
NOR2_X1 U929 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U930 ( .A(n1240), .B(KEYINPUT27), .Z(n1239) );
NAND2_X1 U931 ( .A1(G119), .A2(n1241), .ZN(n1240) );
NOR2_X1 U932 ( .A1(G119), .A2(n1241), .ZN(n1238) );
XOR2_X1 U933 ( .A(KEYINPUT48), .B(G128), .Z(n1241) );
NAND2_X1 U934 ( .A1(G217), .A2(n1242), .ZN(n1226) );
NAND2_X1 U935 ( .A1(G902), .A2(G217), .ZN(n1223) );
XOR2_X1 U936 ( .A(n1243), .B(n1042), .Z(n1207) );
XOR2_X1 U937 ( .A(G472), .B(KEYINPUT43), .Z(n1042) );
XNOR2_X1 U938 ( .A(KEYINPUT7), .B(n1244), .ZN(n1243) );
NOR2_X1 U939 ( .A1(n1043), .A2(KEYINPUT2), .ZN(n1244) );
AND2_X1 U940 ( .A1(n1245), .A2(n1175), .ZN(n1043) );
XNOR2_X1 U941 ( .A(n1155), .B(n1246), .ZN(n1245) );
XOR2_X1 U942 ( .A(n1247), .B(n1158), .Z(n1246) );
INV_X1 U943 ( .A(n1157), .ZN(n1158) );
XOR2_X1 U944 ( .A(n1248), .B(n1249), .Z(n1157) );
XOR2_X1 U945 ( .A(KEYINPUT40), .B(G116), .Z(n1249) );
XOR2_X1 U946 ( .A(n1250), .B(G113), .Z(n1248) );
NAND2_X1 U947 ( .A1(KEYINPUT6), .A2(n1251), .ZN(n1250) );
INV_X1 U948 ( .A(G119), .ZN(n1251) );
NOR2_X1 U949 ( .A1(n1252), .A2(n1253), .ZN(n1247) );
XOR2_X1 U950 ( .A(n1254), .B(KEYINPUT1), .Z(n1253) );
NAND2_X1 U951 ( .A1(n1159), .A2(n1145), .ZN(n1254) );
NOR2_X1 U952 ( .A1(n1145), .A2(n1159), .ZN(n1252) );
INV_X1 U953 ( .A(G101), .ZN(n1159) );
NAND3_X1 U954 ( .A1(n1255), .A2(n1025), .A3(G210), .ZN(n1145) );
XOR2_X1 U955 ( .A(KEYINPUT16), .B(G237), .Z(n1255) );
XNOR2_X1 U956 ( .A(n1256), .B(n1257), .ZN(n1155) );
NAND2_X1 U957 ( .A1(n1258), .A2(n1259), .ZN(n1055) );
OR3_X1 U958 ( .A1(n1204), .A2(n1050), .A3(KEYINPUT9), .ZN(n1259) );
INV_X1 U959 ( .A(n1221), .ZN(n1050) );
NAND2_X1 U960 ( .A1(KEYINPUT9), .A2(n1077), .ZN(n1258) );
AND2_X1 U961 ( .A1(n1221), .A2(n1204), .ZN(n1077) );
NAND3_X1 U962 ( .A1(n1260), .A2(n1261), .A3(n1045), .ZN(n1204) );
NAND2_X1 U963 ( .A1(n1262), .A2(n1039), .ZN(n1045) );
INV_X1 U964 ( .A(G478), .ZN(n1039) );
OR2_X1 U965 ( .A1(G478), .A2(KEYINPUT14), .ZN(n1261) );
NAND3_X1 U966 ( .A1(G478), .A2(n1040), .A3(KEYINPUT14), .ZN(n1260) );
INV_X1 U967 ( .A(n1262), .ZN(n1040) );
NOR2_X1 U968 ( .A1(n1133), .A2(G902), .ZN(n1262) );
XNOR2_X1 U969 ( .A(n1263), .B(n1264), .ZN(n1133) );
XOR2_X1 U970 ( .A(G107), .B(n1265), .Z(n1264) );
XOR2_X1 U971 ( .A(G134), .B(G122), .Z(n1265) );
XOR2_X1 U972 ( .A(n1266), .B(n1267), .Z(n1263) );
AND2_X1 U973 ( .A1(G217), .A2(n1233), .ZN(n1267) );
NOR2_X1 U974 ( .A1(n1242), .A2(G953), .ZN(n1233) );
INV_X1 U975 ( .A(G234), .ZN(n1242) );
XNOR2_X1 U976 ( .A(n1268), .B(n1269), .ZN(n1266) );
NAND2_X1 U977 ( .A1(KEYINPUT61), .A2(n1219), .ZN(n1269) );
INV_X1 U978 ( .A(G116), .ZN(n1219) );
NAND2_X1 U979 ( .A1(n1270), .A2(KEYINPUT5), .ZN(n1268) );
XNOR2_X1 U980 ( .A(n1271), .B(KEYINPUT60), .ZN(n1270) );
XOR2_X1 U981 ( .A(n1272), .B(G475), .Z(n1221) );
NAND2_X1 U982 ( .A1(n1136), .A2(n1175), .ZN(n1272) );
XNOR2_X1 U983 ( .A(n1273), .B(n1274), .ZN(n1136) );
XNOR2_X1 U984 ( .A(n1097), .B(n1275), .ZN(n1274) );
XNOR2_X1 U985 ( .A(n1276), .B(n1277), .ZN(n1275) );
NAND2_X1 U986 ( .A1(KEYINPUT47), .A2(G113), .ZN(n1277) );
NAND2_X1 U987 ( .A1(KEYINPUT18), .A2(n1139), .ZN(n1276) );
XOR2_X1 U988 ( .A(G125), .B(G140), .Z(n1097) );
XOR2_X1 U989 ( .A(n1278), .B(n1279), .Z(n1273) );
XOR2_X1 U990 ( .A(G122), .B(n1280), .Z(n1279) );
NOR2_X1 U991 ( .A1(KEYINPUT20), .A2(n1281), .ZN(n1280) );
XOR2_X1 U992 ( .A(n1282), .B(n1283), .Z(n1281) );
NOR2_X1 U993 ( .A1(KEYINPUT36), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U994 ( .A(G143), .B(n1285), .ZN(n1282) );
AND3_X1 U995 ( .A1(G214), .A2(n1025), .A3(n1286), .ZN(n1285) );
NAND2_X1 U996 ( .A1(KEYINPUT34), .A2(n1200), .ZN(n1278) );
AND3_X1 U997 ( .A1(n1075), .A2(n1211), .A3(n1068), .ZN(n1183) );
INV_X1 U998 ( .A(n1186), .ZN(n1068) );
NAND2_X1 U999 ( .A1(n1071), .A2(n1044), .ZN(n1186) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1287), .ZN(n1044) );
INV_X1 U1001 ( .A(n1062), .ZN(n1071) );
XOR2_X1 U1002 ( .A(n1049), .B(n1047), .Z(n1062) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1287), .ZN(n1047) );
NAND2_X1 U1004 ( .A1(n1286), .A2(n1175), .ZN(n1287) );
INV_X1 U1005 ( .A(G237), .ZN(n1286) );
AND2_X1 U1006 ( .A1(n1288), .A2(n1175), .ZN(n1049) );
XOR2_X1 U1007 ( .A(n1289), .B(n1290), .Z(n1288) );
INV_X1 U1008 ( .A(n1171), .ZN(n1290) );
XOR2_X1 U1009 ( .A(n1291), .B(n1292), .Z(n1171) );
INV_X1 U1010 ( .A(n1123), .ZN(n1292) );
XOR2_X1 U1011 ( .A(n1293), .B(n1294), .Z(n1123) );
XOR2_X1 U1012 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1013 ( .A(G116), .B(G113), .Z(n1296) );
XOR2_X1 U1014 ( .A(KEYINPUT41), .B(G119), .Z(n1295) );
XOR2_X1 U1015 ( .A(n1297), .B(n1298), .Z(n1293) );
XOR2_X1 U1016 ( .A(G104), .B(G101), .Z(n1298) );
NAND2_X1 U1017 ( .A1(KEYINPUT59), .A2(n1299), .ZN(n1297) );
INV_X1 U1018 ( .A(G107), .ZN(n1299) );
NAND2_X1 U1019 ( .A1(KEYINPUT54), .A2(n1122), .ZN(n1291) );
XOR2_X1 U1020 ( .A(G110), .B(G122), .Z(n1122) );
NAND2_X1 U1021 ( .A1(n1199), .A2(n1198), .ZN(n1289) );
NAND2_X1 U1022 ( .A1(n1300), .A2(n1301), .ZN(n1198) );
NAND2_X1 U1023 ( .A1(G224), .A2(n1025), .ZN(n1301) );
XOR2_X1 U1024 ( .A(n1256), .B(G125), .Z(n1300) );
NAND3_X1 U1025 ( .A1(n1302), .A2(n1025), .A3(G224), .ZN(n1199) );
XNOR2_X1 U1026 ( .A(G125), .B(n1256), .ZN(n1302) );
XOR2_X1 U1027 ( .A(n1303), .B(G128), .Z(n1256) );
NAND2_X1 U1028 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1029 ( .A1(G143), .A2(n1200), .ZN(n1305) );
XOR2_X1 U1030 ( .A(KEYINPUT19), .B(n1306), .Z(n1304) );
NOR2_X1 U1031 ( .A1(G143), .A2(n1200), .ZN(n1306) );
INV_X1 U1032 ( .A(G146), .ZN(n1200) );
NAND2_X1 U1033 ( .A1(n1307), .A2(n1080), .ZN(n1211) );
NAND3_X1 U1034 ( .A1(n1215), .A2(n1025), .A3(G952), .ZN(n1080) );
NAND4_X1 U1035 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1120), .ZN(n1307) );
INV_X1 U1036 ( .A(G898), .ZN(n1120) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1215) );
AND2_X1 U1038 ( .A1(n1308), .A2(n1078), .ZN(n1075) );
XNOR2_X1 U1039 ( .A(n1309), .B(G469), .ZN(n1078) );
NAND2_X1 U1040 ( .A1(KEYINPUT62), .A2(n1310), .ZN(n1309) );
INV_X1 U1041 ( .A(n1035), .ZN(n1310) );
NAND2_X1 U1042 ( .A1(n1311), .A2(n1175), .ZN(n1035) );
XOR2_X1 U1043 ( .A(n1312), .B(n1169), .Z(n1311) );
AND2_X1 U1044 ( .A1(G227), .A2(n1025), .ZN(n1169) );
INV_X1 U1045 ( .A(G953), .ZN(n1025) );
XOR2_X1 U1046 ( .A(n1313), .B(n1314), .Z(n1312) );
NOR2_X1 U1047 ( .A1(KEYINPUT23), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1048 ( .A(n1222), .B(n1316), .Z(n1315) );
XOR2_X1 U1049 ( .A(KEYINPUT30), .B(G140), .Z(n1316) );
NAND3_X1 U1050 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1313) );
OR2_X1 U1051 ( .A1(n1320), .A2(n1257), .ZN(n1319) );
NAND2_X1 U1052 ( .A1(KEYINPUT46), .A2(n1321), .ZN(n1318) );
NAND2_X1 U1053 ( .A1(n1322), .A2(n1320), .ZN(n1321) );
XOR2_X1 U1054 ( .A(KEYINPUT58), .B(n1165), .Z(n1322) );
INV_X1 U1055 ( .A(n1257), .ZN(n1165) );
NAND2_X1 U1056 ( .A1(n1323), .A2(n1324), .ZN(n1317) );
INV_X1 U1057 ( .A(KEYINPUT46), .ZN(n1324) );
NAND2_X1 U1058 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
OR2_X1 U1059 ( .A1(n1257), .A2(KEYINPUT58), .ZN(n1326) );
NAND3_X1 U1060 ( .A1(n1320), .A2(n1257), .A3(KEYINPUT58), .ZN(n1325) );
XNOR2_X1 U1061 ( .A(n1107), .B(n1105), .ZN(n1257) );
INV_X1 U1062 ( .A(n1108), .ZN(n1105) );
XOR2_X1 U1063 ( .A(n1284), .B(G134), .Z(n1108) );
INV_X1 U1064 ( .A(G131), .ZN(n1284) );
INV_X1 U1065 ( .A(G137), .ZN(n1107) );
XNOR2_X1 U1066 ( .A(n1163), .B(KEYINPUT56), .ZN(n1320) );
XOR2_X1 U1067 ( .A(n1327), .B(n1328), .Z(n1163) );
XOR2_X1 U1068 ( .A(KEYINPUT28), .B(G101), .Z(n1328) );
XNOR2_X1 U1069 ( .A(n1329), .B(n1100), .ZN(n1327) );
XNOR2_X1 U1070 ( .A(G146), .B(n1271), .ZN(n1100) );
XOR2_X1 U1071 ( .A(G128), .B(G143), .Z(n1271) );
NAND2_X1 U1072 ( .A1(n1330), .A2(KEYINPUT15), .ZN(n1329) );
XOR2_X1 U1073 ( .A(n1139), .B(G107), .Z(n1330) );
INV_X1 U1074 ( .A(G104), .ZN(n1139) );
XOR2_X1 U1075 ( .A(KEYINPUT29), .B(n1074), .Z(n1308) );
INV_X1 U1076 ( .A(n1046), .ZN(n1074) );
NAND2_X1 U1077 ( .A1(G221), .A2(n1331), .ZN(n1046) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1175), .ZN(n1331) );
INV_X1 U1079 ( .A(G902), .ZN(n1175) );
INV_X1 U1080 ( .A(G110), .ZN(n1222) );
endmodule


