//Key = 0110011000010001101000010110001001011101000011011011110111010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343;

XNOR2_X1 U736 ( .A(G107), .B(n1019), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1022), .A2(n1023), .A3(G953), .A4(n1024), .ZN(n1021) );
NOR4_X1 U739 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1023) );
NOR3_X1 U740 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1025) );
NOR2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1030) );
XNOR2_X1 U745 ( .A(KEYINPUT33), .B(n1040), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1041), .A2(n1040), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1022) );
NAND3_X1 U748 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND3_X1 U750 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
XNOR2_X1 U751 ( .A(KEYINPUT46), .B(n1028), .ZN(n1050) );
NAND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1047) );
NAND3_X1 U753 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND3_X1 U755 ( .A1(n1059), .A2(n1051), .A3(n1060), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1054) );
XNOR2_X1 U757 ( .A(n1058), .B(KEYINPUT5), .ZN(n1061) );
INV_X1 U758 ( .A(n1027), .ZN(n1058) );
INV_X1 U759 ( .A(n1028), .ZN(n1052) );
NOR3_X1 U760 ( .A1(n1024), .A2(G953), .A3(G952), .ZN(n1020) );
AND2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1024) );
NOR4_X1 U762 ( .A1(n1065), .A2(n1060), .A3(n1066), .A4(n1067), .ZN(n1064) );
XNOR2_X1 U763 ( .A(G469), .B(n1068), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1069), .A2(KEYINPUT7), .ZN(n1068) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
XNOR2_X1 U766 ( .A(KEYINPUT63), .B(G472), .ZN(n1071) );
NOR4_X1 U767 ( .A1(n1033), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1063) );
XOR2_X1 U768 ( .A(KEYINPUT9), .B(n1075), .Z(n1074) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U770 ( .A(KEYINPUT63), .B(G472), .Z(n1077) );
XNOR2_X1 U771 ( .A(n1078), .B(n1079), .ZN(n1073) );
NAND2_X1 U772 ( .A1(KEYINPUT55), .A2(n1080), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1081), .B(n1082), .Z(G72) );
NAND2_X1 U774 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U775 ( .A1(G900), .A2(G227), .ZN(n1083) );
NAND4_X1 U776 ( .A1(KEYINPUT48), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1081) );
NAND3_X1 U777 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND2_X1 U778 ( .A1(G953), .A2(n1090), .ZN(n1085) );
NAND2_X1 U779 ( .A1(G900), .A2(n1087), .ZN(n1090) );
OR2_X1 U780 ( .A1(n1088), .A2(n1087), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1087) );
XNOR2_X1 U782 ( .A(n1093), .B(n1094), .ZN(n1092) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(n1091) );
NOR2_X1 U784 ( .A1(KEYINPUT58), .A2(n1097), .ZN(n1096) );
XOR2_X1 U785 ( .A(n1098), .B(KEYINPUT51), .Z(n1097) );
NAND2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U788 ( .A(KEYINPUT3), .B(n1103), .ZN(n1102) );
XNOR2_X1 U789 ( .A(KEYINPUT4), .B(G134), .ZN(n1101) );
XOR2_X1 U790 ( .A(n1104), .B(KEYINPUT8), .Z(n1099) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U792 ( .A(KEYINPUT3), .B(n1103), .Z(n1106) );
XOR2_X1 U793 ( .A(KEYINPUT4), .B(G134), .Z(n1105) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U796 ( .A(n1111), .B(n1112), .ZN(n1110) );
NOR2_X1 U797 ( .A1(KEYINPUT29), .A2(n1113), .ZN(n1111) );
NOR2_X1 U798 ( .A1(G898), .A2(n1089), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1107) );
NAND3_X1 U800 ( .A1(KEYINPUT35), .A2(n1116), .A3(n1089), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U802 ( .A1(G953), .A2(n1119), .ZN(n1114) );
NAND2_X1 U803 ( .A1(G224), .A2(n1120), .ZN(n1119) );
XNOR2_X1 U804 ( .A(KEYINPUT28), .B(n1121), .ZN(n1120) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND3_X1 U807 ( .A1(G902), .A2(n1126), .A3(n1127), .ZN(n1124) );
XNOR2_X1 U808 ( .A(KEYINPUT6), .B(n1128), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1129), .ZN(G63) );
NOR2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U811 ( .A(KEYINPUT34), .B(n1132), .Z(n1131) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
AND2_X1 U813 ( .A1(n1134), .A2(n1133), .ZN(n1130) );
NAND2_X1 U814 ( .A1(n1135), .A2(G478), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1136), .ZN(G60) );
XNOR2_X1 U816 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR3_X1 U817 ( .A1(n1139), .A2(KEYINPUT17), .A3(n1140), .ZN(n1138) );
INV_X1 U818 ( .A(n1135), .ZN(n1139) );
XNOR2_X1 U819 ( .A(G104), .B(n1141), .ZN(G6) );
NAND3_X1 U820 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
XNOR2_X1 U821 ( .A(n1051), .B(KEYINPUT50), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1122), .A2(n1145), .ZN(G57) );
XOR2_X1 U823 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U824 ( .A(KEYINPUT57), .B(n1148), .Z(n1147) );
NOR4_X1 U825 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NOR3_X1 U826 ( .A1(n1153), .A2(n1093), .A3(n1154), .ZN(n1150) );
NOR3_X1 U827 ( .A1(n1155), .A2(n1093), .A3(n1156), .ZN(n1149) );
XOR2_X1 U828 ( .A(n1157), .B(n1158), .Z(n1146) );
NAND2_X1 U829 ( .A1(KEYINPUT36), .A2(n1159), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1135), .A2(G472), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1122), .A2(n1160), .ZN(G54) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U833 ( .A1(KEYINPUT14), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U834 ( .A(n1164), .B(n1165), .ZN(n1163) );
XOR2_X1 U835 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U837 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U838 ( .A(KEYINPUT52), .B(n1172), .Z(n1168) );
NOR2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1172) );
XNOR2_X1 U840 ( .A(KEYINPUT25), .B(n1153), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1135), .A2(G469), .ZN(n1161) );
NOR2_X1 U842 ( .A1(n1122), .A2(n1173), .ZN(G51) );
NOR3_X1 U843 ( .A1(n1078), .A2(n1174), .A3(n1175), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U845 ( .A1(n1042), .A2(n1178), .ZN(n1176) );
AND3_X1 U846 ( .A1(n1177), .A2(n1080), .A3(n1135), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1179), .A2(n1042), .ZN(n1135) );
INV_X1 U848 ( .A(n1128), .ZN(n1042) );
NAND3_X1 U849 ( .A1(n1117), .A2(n1180), .A3(n1181), .ZN(n1128) );
INV_X1 U850 ( .A(n1088), .ZN(n1181) );
NAND4_X1 U851 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1088) );
AND3_X1 U852 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
NAND2_X1 U853 ( .A1(n1142), .A2(n1189), .ZN(n1184) );
NAND2_X1 U854 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND3_X1 U855 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NAND2_X1 U856 ( .A1(n1195), .A2(n1196), .ZN(n1190) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U858 ( .A1(n1199), .A2(n1049), .ZN(n1182) );
XOR2_X1 U859 ( .A(n1200), .B(KEYINPUT45), .Z(n1199) );
XNOR2_X1 U860 ( .A(KEYINPUT44), .B(n1118), .ZN(n1180) );
AND4_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1117) );
AND3_X1 U862 ( .A1(n1205), .A2(n1019), .A3(n1206), .ZN(n1204) );
NAND3_X1 U863 ( .A1(n1051), .A2(n1143), .A3(n1207), .ZN(n1019) );
NAND2_X1 U864 ( .A1(n1143), .A2(n1208), .ZN(n1203) );
NAND2_X1 U865 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U866 ( .A1(n1142), .A2(n1051), .ZN(n1210) );
NAND2_X1 U867 ( .A1(n1057), .A2(n1044), .ZN(n1209) );
NOR2_X1 U868 ( .A1(n1089), .A2(G952), .ZN(n1122) );
XNOR2_X1 U869 ( .A(G146), .B(n1211), .ZN(G48) );
NAND4_X1 U870 ( .A1(n1142), .A2(n1194), .A3(n1192), .A4(n1212), .ZN(n1211) );
XNOR2_X1 U871 ( .A(KEYINPUT2), .B(n1193), .ZN(n1212) );
XNOR2_X1 U872 ( .A(G143), .B(n1183), .ZN(G45) );
NAND3_X1 U873 ( .A1(n1062), .A2(n1192), .A3(n1213), .ZN(n1183) );
NOR3_X1 U874 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
XOR2_X1 U875 ( .A(G140), .B(n1217), .Z(G42) );
NOR3_X1 U876 ( .A1(n1218), .A2(n1219), .A3(n1038), .ZN(n1217) );
INV_X1 U877 ( .A(n1195), .ZN(n1219) );
XNOR2_X1 U878 ( .A(KEYINPUT59), .B(n1197), .ZN(n1218) );
XNOR2_X1 U879 ( .A(G137), .B(n1186), .ZN(G39) );
NAND3_X1 U880 ( .A1(n1194), .A2(n1044), .A3(n1195), .ZN(n1186) );
XNOR2_X1 U881 ( .A(G134), .B(n1188), .ZN(G36) );
NAND3_X1 U882 ( .A1(n1195), .A2(n1207), .A3(n1062), .ZN(n1188) );
XNOR2_X1 U883 ( .A(G131), .B(n1220), .ZN(G33) );
NAND3_X1 U884 ( .A1(n1195), .A2(n1221), .A3(n1062), .ZN(n1220) );
XNOR2_X1 U885 ( .A(KEYINPUT54), .B(n1038), .ZN(n1221) );
INV_X1 U886 ( .A(n1142), .ZN(n1038) );
NOR3_X1 U887 ( .A1(n1222), .A2(n1215), .A3(n1027), .ZN(n1195) );
NAND2_X1 U888 ( .A1(n1223), .A2(n1224), .ZN(n1027) );
XNOR2_X1 U889 ( .A(KEYINPUT61), .B(n1059), .ZN(n1223) );
INV_X1 U890 ( .A(n1193), .ZN(n1215) );
XOR2_X1 U891 ( .A(n1187), .B(n1225), .Z(G30) );
XNOR2_X1 U892 ( .A(G128), .B(KEYINPUT19), .ZN(n1225) );
NAND4_X1 U893 ( .A1(n1194), .A2(n1207), .A3(n1192), .A4(n1193), .ZN(n1187) );
XNOR2_X1 U894 ( .A(G101), .B(n1201), .ZN(G3) );
NAND3_X1 U895 ( .A1(n1044), .A2(n1143), .A3(n1062), .ZN(n1201) );
NOR2_X1 U896 ( .A1(n1226), .A2(n1227), .ZN(n1143) );
INV_X1 U897 ( .A(n1192), .ZN(n1226) );
XOR2_X1 U898 ( .A(G125), .B(n1228), .Z(G27) );
NOR2_X1 U899 ( .A1(n1229), .A2(n1200), .ZN(n1228) );
NAND4_X1 U900 ( .A1(n1142), .A2(n1046), .A3(n1057), .A4(n1193), .ZN(n1200) );
NAND2_X1 U901 ( .A1(n1028), .A2(n1230), .ZN(n1193) );
NAND4_X1 U902 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1232), .ZN(n1230) );
INV_X1 U903 ( .A(G900), .ZN(n1232) );
XNOR2_X1 U904 ( .A(G122), .B(n1118), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1233), .A2(n1051), .A3(n1234), .A4(n1235), .ZN(n1118) );
INV_X1 U906 ( .A(n1026), .ZN(n1051) );
NAND2_X1 U907 ( .A1(n1236), .A2(n1237), .ZN(n1026) );
XOR2_X1 U908 ( .A(n1238), .B(KEYINPUT49), .Z(n1236) );
XNOR2_X1 U909 ( .A(G119), .B(n1202), .ZN(G21) );
NAND3_X1 U910 ( .A1(n1194), .A2(n1044), .A3(n1233), .ZN(n1202) );
NOR2_X1 U911 ( .A1(n1238), .A2(n1237), .ZN(n1194) );
XOR2_X1 U912 ( .A(n1239), .B(G116), .Z(G18) );
NAND2_X1 U913 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
OR2_X1 U914 ( .A1(n1205), .A2(KEYINPUT21), .ZN(n1241) );
OR2_X1 U915 ( .A1(n1242), .A2(n1229), .ZN(n1205) );
NAND3_X1 U916 ( .A1(n1049), .A2(n1242), .A3(KEYINPUT21), .ZN(n1240) );
OR4_X1 U917 ( .A1(n1040), .A2(n1198), .A3(n1041), .A4(n1227), .ZN(n1242) );
INV_X1 U918 ( .A(n1207), .ZN(n1041) );
NOR2_X1 U919 ( .A1(n1235), .A2(n1214), .ZN(n1207) );
INV_X1 U920 ( .A(n1234), .ZN(n1214) );
INV_X1 U921 ( .A(n1062), .ZN(n1198) );
XNOR2_X1 U922 ( .A(G113), .B(n1206), .ZN(G15) );
NAND3_X1 U923 ( .A1(n1142), .A2(n1062), .A3(n1233), .ZN(n1206) );
NOR3_X1 U924 ( .A1(n1229), .A2(n1227), .A3(n1040), .ZN(n1233) );
INV_X1 U925 ( .A(n1046), .ZN(n1040) );
NOR2_X1 U926 ( .A1(n1037), .A2(n1243), .ZN(n1046) );
NOR2_X1 U927 ( .A1(n1072), .A2(n1237), .ZN(n1062) );
NOR2_X1 U928 ( .A1(n1234), .A2(n1216), .ZN(n1142) );
INV_X1 U929 ( .A(n1235), .ZN(n1216) );
XNOR2_X1 U930 ( .A(G110), .B(n1244), .ZN(G12) );
NAND4_X1 U931 ( .A1(n1245), .A2(n1246), .A3(n1057), .A4(n1247), .ZN(n1244) );
NOR2_X1 U932 ( .A1(n1227), .A2(n1033), .ZN(n1247) );
INV_X1 U933 ( .A(n1044), .ZN(n1033) );
NOR2_X1 U934 ( .A1(n1234), .A2(n1235), .ZN(n1044) );
XOR2_X1 U935 ( .A(n1248), .B(n1140), .Z(n1235) );
INV_X1 U936 ( .A(G475), .ZN(n1140) );
NAND2_X1 U937 ( .A1(n1179), .A2(n1137), .ZN(n1248) );
NAND2_X1 U938 ( .A1(n1249), .A2(n1250), .ZN(n1137) );
NAND2_X1 U939 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U940 ( .A(KEYINPUT39), .B(n1253), .Z(n1249) );
NOR2_X1 U941 ( .A1(n1251), .A2(n1252), .ZN(n1253) );
XNOR2_X1 U942 ( .A(n1254), .B(n1255), .ZN(n1252) );
XNOR2_X1 U943 ( .A(KEYINPUT16), .B(n1256), .ZN(n1255) );
XNOR2_X1 U944 ( .A(G104), .B(G113), .ZN(n1254) );
XOR2_X1 U945 ( .A(n1257), .B(n1258), .Z(n1251) );
NOR2_X1 U946 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
AND2_X1 U947 ( .A1(n1261), .A2(G146), .ZN(n1259) );
XOR2_X1 U948 ( .A(n1098), .B(KEYINPUT20), .Z(n1261) );
NAND3_X1 U949 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1257) );
NAND2_X1 U950 ( .A1(KEYINPUT24), .A2(n1265), .ZN(n1264) );
NAND3_X1 U951 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1263) );
INV_X1 U952 ( .A(KEYINPUT24), .ZN(n1267) );
OR2_X1 U953 ( .A1(n1268), .A2(n1266), .ZN(n1262) );
NOR2_X1 U954 ( .A1(n1269), .A2(n1265), .ZN(n1266) );
XNOR2_X1 U955 ( .A(n1270), .B(G143), .ZN(n1265) );
NAND3_X1 U956 ( .A1(n1271), .A2(n1272), .A3(G214), .ZN(n1270) );
XNOR2_X1 U957 ( .A(KEYINPUT37), .B(n1089), .ZN(n1271) );
INV_X1 U958 ( .A(KEYINPUT15), .ZN(n1269) );
INV_X1 U959 ( .A(G131), .ZN(n1268) );
XNOR2_X1 U960 ( .A(n1273), .B(G478), .ZN(n1234) );
NAND2_X1 U961 ( .A1(n1133), .A2(n1179), .ZN(n1273) );
XOR2_X1 U962 ( .A(n1274), .B(n1275), .Z(n1133) );
AND2_X1 U963 ( .A1(n1276), .A2(G217), .ZN(n1275) );
NAND2_X1 U964 ( .A1(n1277), .A2(KEYINPUT26), .ZN(n1274) );
XOR2_X1 U965 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U966 ( .A(G134), .B(n1280), .ZN(n1279) );
XNOR2_X1 U967 ( .A(KEYINPUT22), .B(KEYINPUT13), .ZN(n1280) );
XOR2_X1 U968 ( .A(n1281), .B(n1282), .Z(n1278) );
XNOR2_X1 U969 ( .A(n1283), .B(n1284), .ZN(n1282) );
NAND2_X1 U970 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
OR2_X1 U971 ( .A1(n1256), .A2(G116), .ZN(n1286) );
XOR2_X1 U972 ( .A(n1287), .B(KEYINPUT41), .Z(n1285) );
NAND2_X1 U973 ( .A1(G116), .A2(n1256), .ZN(n1287) );
AND2_X1 U974 ( .A1(n1028), .A2(n1288), .ZN(n1227) );
NAND4_X1 U975 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1121), .ZN(n1288) );
INV_X1 U976 ( .A(G898), .ZN(n1121) );
NAND3_X1 U977 ( .A1(n1231), .A2(n1089), .A3(G952), .ZN(n1028) );
NAND2_X1 U978 ( .A1(G237), .A2(G234), .ZN(n1231) );
INV_X1 U979 ( .A(n1197), .ZN(n1057) );
NAND2_X1 U980 ( .A1(n1237), .A2(n1072), .ZN(n1197) );
INV_X1 U981 ( .A(n1238), .ZN(n1072) );
XOR2_X1 U982 ( .A(n1289), .B(n1127), .Z(n1238) );
AND2_X1 U983 ( .A1(G217), .A2(n1290), .ZN(n1127) );
NAND2_X1 U984 ( .A1(n1125), .A2(n1179), .ZN(n1289) );
XNOR2_X1 U985 ( .A(n1291), .B(n1292), .ZN(n1125) );
XNOR2_X1 U986 ( .A(n1293), .B(n1103), .ZN(n1292) );
NAND2_X1 U987 ( .A1(G221), .A2(n1276), .ZN(n1293) );
AND2_X1 U988 ( .A1(G234), .A2(n1089), .ZN(n1276) );
XOR2_X1 U989 ( .A(n1294), .B(n1295), .Z(n1291) );
NOR2_X1 U990 ( .A1(n1296), .A2(n1260), .ZN(n1295) );
NOR2_X1 U991 ( .A1(n1098), .A2(G146), .ZN(n1260) );
AND2_X1 U992 ( .A1(n1098), .A2(G146), .ZN(n1296) );
XNOR2_X1 U993 ( .A(G125), .B(G140), .ZN(n1098) );
NAND2_X1 U994 ( .A1(KEYINPUT53), .A2(n1297), .ZN(n1294) );
XNOR2_X1 U995 ( .A(n1298), .B(n1299), .ZN(n1297) );
NOR2_X1 U996 ( .A1(KEYINPUT42), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U997 ( .A(G119), .B(G128), .ZN(n1300) );
XNOR2_X1 U998 ( .A(n1070), .B(G472), .ZN(n1237) );
INV_X1 U999 ( .A(n1076), .ZN(n1070) );
NAND2_X1 U1000 ( .A1(n1301), .A2(n1179), .ZN(n1076) );
XNOR2_X1 U1001 ( .A(n1158), .B(n1302), .ZN(n1301) );
XOR2_X1 U1002 ( .A(n1303), .B(KEYINPUT43), .Z(n1302) );
NAND2_X1 U1003 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1004 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1005 ( .A1(KEYINPUT18), .A2(n1093), .ZN(n1307) );
XNOR2_X1 U1006 ( .A(n1155), .B(n1156), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(KEYINPUT18), .A2(n1308), .ZN(n1304) );
OR2_X1 U1008 ( .A1(n1151), .A2(n1152), .ZN(n1308) );
NOR3_X1 U1009 ( .A1(n1153), .A2(n1309), .A3(n1156), .ZN(n1152) );
NOR3_X1 U1010 ( .A1(n1154), .A2(n1309), .A3(n1155), .ZN(n1151) );
INV_X1 U1011 ( .A(n1156), .ZN(n1154) );
XNOR2_X1 U1012 ( .A(n1310), .B(KEYINPUT12), .ZN(n1156) );
XNOR2_X1 U1013 ( .A(n1311), .B(G101), .ZN(n1158) );
NAND3_X1 U1014 ( .A1(n1272), .A2(n1089), .A3(G210), .ZN(n1311) );
OR2_X1 U1015 ( .A1(n1192), .A2(KEYINPUT10), .ZN(n1246) );
NOR2_X1 U1016 ( .A1(n1229), .A2(n1222), .ZN(n1192) );
INV_X1 U1017 ( .A(n1049), .ZN(n1229) );
NAND2_X1 U1018 ( .A1(KEYINPUT10), .A2(n1312), .ZN(n1245) );
NAND2_X1 U1019 ( .A1(n1049), .A2(n1222), .ZN(n1312) );
INV_X1 U1020 ( .A(n1035), .ZN(n1222) );
NOR2_X1 U1021 ( .A1(n1243), .A2(n1313), .ZN(n1035) );
INV_X1 U1022 ( .A(n1037), .ZN(n1313) );
XOR2_X1 U1023 ( .A(n1069), .B(G469), .Z(n1037) );
AND2_X1 U1024 ( .A1(n1314), .A2(n1179), .ZN(n1069) );
XOR2_X1 U1025 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1026 ( .A(n1317), .B(n1166), .ZN(n1316) );
NAND2_X1 U1027 ( .A1(G227), .A2(n1089), .ZN(n1166) );
NOR2_X1 U1028 ( .A1(KEYINPUT31), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1029 ( .A(KEYINPUT23), .B(n1164), .Z(n1318) );
XOR2_X1 U1030 ( .A(G140), .B(G110), .Z(n1164) );
XNOR2_X1 U1031 ( .A(n1319), .B(n1170), .ZN(n1315) );
XOR2_X1 U1032 ( .A(n1320), .B(n1321), .Z(n1170) );
XNOR2_X1 U1033 ( .A(KEYINPUT62), .B(n1322), .ZN(n1320) );
NOR2_X1 U1034 ( .A1(G101), .A2(KEYINPUT60), .ZN(n1322) );
NAND2_X1 U1035 ( .A1(KEYINPUT1), .A2(n1153), .ZN(n1319) );
INV_X1 U1036 ( .A(n1155), .ZN(n1153) );
XNOR2_X1 U1037 ( .A(n1094), .B(n1323), .ZN(n1155) );
NOR3_X1 U1038 ( .A1(KEYINPUT0), .A2(n1324), .A3(n1325), .ZN(n1323) );
NOR2_X1 U1039 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
XNOR2_X1 U1040 ( .A(G134), .B(n1103), .ZN(n1327) );
INV_X1 U1041 ( .A(KEYINPUT47), .ZN(n1326) );
NOR3_X1 U1042 ( .A1(KEYINPUT47), .A2(G134), .A3(n1103), .ZN(n1324) );
XOR2_X1 U1043 ( .A(G137), .B(KEYINPUT56), .Z(n1103) );
XNOR2_X1 U1044 ( .A(G131), .B(KEYINPUT32), .ZN(n1094) );
XOR2_X1 U1045 ( .A(n1065), .B(KEYINPUT40), .Z(n1243) );
INV_X1 U1046 ( .A(n1036), .ZN(n1065) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1290), .ZN(n1036) );
NAND2_X1 U1048 ( .A1(n1328), .A2(G234), .ZN(n1290) );
XNOR2_X1 U1049 ( .A(G902), .B(KEYINPUT27), .ZN(n1328) );
NOR2_X1 U1050 ( .A1(n1059), .A2(n1060), .ZN(n1049) );
INV_X1 U1051 ( .A(n1224), .ZN(n1060) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1329), .ZN(n1224) );
XNOR2_X1 U1053 ( .A(n1078), .B(n1080), .ZN(n1059) );
INV_X1 U1054 ( .A(n1178), .ZN(n1080) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1329), .ZN(n1178) );
NAND2_X1 U1056 ( .A1(n1272), .A2(n1179), .ZN(n1329) );
INV_X1 U1057 ( .A(G902), .ZN(n1179) );
INV_X1 U1058 ( .A(G237), .ZN(n1272) );
NOR2_X1 U1059 ( .A1(n1177), .A2(G902), .ZN(n1078) );
XOR2_X1 U1060 ( .A(n1330), .B(n1331), .Z(n1177) );
XOR2_X1 U1061 ( .A(KEYINPUT38), .B(G125), .Z(n1331) );
XOR2_X1 U1062 ( .A(n1332), .B(n1333), .Z(n1330) );
AND2_X1 U1063 ( .A1(n1089), .A2(G224), .ZN(n1333) );
INV_X1 U1064 ( .A(G953), .ZN(n1089) );
NAND2_X1 U1065 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
NAND2_X1 U1066 ( .A1(n1336), .A2(n1112), .ZN(n1335) );
INV_X1 U1067 ( .A(n1337), .ZN(n1112) );
XOR2_X1 U1068 ( .A(n1338), .B(n1321), .Z(n1336) );
XNOR2_X1 U1069 ( .A(n1339), .B(n1093), .ZN(n1321) );
NAND2_X1 U1070 ( .A1(n1340), .A2(n1337), .ZN(n1334) );
XOR2_X1 U1071 ( .A(n1341), .B(n1256), .Z(n1337) );
INV_X1 U1072 ( .A(G122), .ZN(n1256) );
NAND2_X1 U1073 ( .A1(KEYINPUT30), .A2(n1298), .ZN(n1341) );
INV_X1 U1074 ( .A(G110), .ZN(n1298) );
XNOR2_X1 U1075 ( .A(n1093), .B(n1113), .ZN(n1340) );
XNOR2_X1 U1076 ( .A(n1338), .B(n1339), .ZN(n1113) );
XOR2_X1 U1077 ( .A(G104), .B(n1281), .Z(n1339) );
XNOR2_X1 U1078 ( .A(G107), .B(KEYINPUT11), .ZN(n1281) );
XOR2_X1 U1079 ( .A(n1310), .B(G101), .Z(n1338) );
XNOR2_X1 U1080 ( .A(G113), .B(n1342), .ZN(n1310) );
XNOR2_X1 U1081 ( .A(n1343), .B(G116), .ZN(n1342) );
INV_X1 U1082 ( .A(G119), .ZN(n1343) );
INV_X1 U1083 ( .A(n1309), .ZN(n1093) );
XNOR2_X1 U1084 ( .A(G146), .B(n1284), .ZN(n1309) );
XOR2_X1 U1085 ( .A(G128), .B(G143), .Z(n1284) );
endmodule


