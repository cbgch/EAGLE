//Key = 0110000011000100110100100101101111100111110101001010100010010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U749 ( .A(n1047), .B(n1048), .Z(G9) );
NAND4_X1 U750 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NOR2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
XOR2_X1 U752 ( .A(n1055), .B(KEYINPUT52), .Z(n1049) );
NOR2_X1 U753 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR3_X1 U754 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NOR2_X1 U755 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
INV_X1 U756 ( .A(n1050), .ZN(n1062) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U758 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR4_X1 U759 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U761 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U762 ( .A1(KEYINPUT7), .A2(n1076), .ZN(n1074) );
NOR3_X1 U763 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1070) );
XOR2_X1 U764 ( .A(KEYINPUT39), .B(n1080), .Z(n1077) );
NOR2_X1 U765 ( .A1(n1053), .A2(n1081), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1082), .A2(n1083), .ZN(n1066) );
AND3_X1 U767 ( .A1(KEYINPUT7), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR4_X1 U768 ( .A1(n1068), .A2(n1086), .A3(n1073), .A4(n1081), .ZN(n1063) );
NOR2_X1 U769 ( .A1(n1087), .A2(n1052), .ZN(n1086) );
NOR2_X1 U770 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U771 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1058) );
NAND4_X1 U772 ( .A1(n1080), .A2(n1093), .A3(n1094), .A4(n1084), .ZN(n1092) );
NOR2_X1 U773 ( .A1(n1068), .A2(n1095), .ZN(n1094) );
NOR2_X1 U774 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
INV_X1 U775 ( .A(n1083), .ZN(n1068) );
NOR3_X1 U776 ( .A1(n1098), .A2(G953), .A3(G952), .ZN(n1056) );
INV_X1 U777 ( .A(n1090), .ZN(n1098) );
NAND4_X1 U778 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1090) );
NOR4_X1 U779 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
XNOR2_X1 U780 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U781 ( .A1(n1109), .A2(KEYINPUT4), .ZN(n1108) );
XOR2_X1 U782 ( .A(n1110), .B(n1111), .Z(n1105) );
NOR2_X1 U783 ( .A1(G469), .A2(KEYINPUT20), .ZN(n1111) );
NOR2_X1 U784 ( .A1(n1112), .A2(n1113), .ZN(n1104) );
INV_X1 U785 ( .A(G472), .ZN(n1113) );
NOR2_X1 U786 ( .A1(G902), .A2(n1114), .ZN(n1112) );
NOR2_X1 U787 ( .A1(n1065), .A2(n1115), .ZN(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT49), .B(n1116), .Z(n1115) );
XOR2_X1 U789 ( .A(KEYINPUT17), .B(n1117), .Z(n1100) );
XOR2_X1 U790 ( .A(n1118), .B(n1119), .Z(G72) );
XOR2_X1 U791 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U792 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U793 ( .A(n1124), .B(n1125), .Z(n1122) );
XNOR2_X1 U794 ( .A(n1126), .B(n1127), .ZN(n1125) );
XOR2_X1 U795 ( .A(KEYINPUT61), .B(n1128), .Z(n1124) );
NAND2_X1 U796 ( .A1(n1129), .A2(n1091), .ZN(n1120) );
NOR2_X1 U797 ( .A1(n1130), .A2(n1091), .ZN(n1118) );
NOR2_X1 U798 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U799 ( .A(n1133), .B(n1134), .Z(G69) );
NOR2_X1 U800 ( .A1(n1135), .A2(n1091), .ZN(n1134) );
AND2_X1 U801 ( .A1(G224), .A2(G898), .ZN(n1135) );
NOR2_X1 U802 ( .A1(KEYINPUT26), .A2(n1136), .ZN(n1133) );
XOR2_X1 U803 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U804 ( .A1(n1139), .A2(G953), .ZN(n1138) );
NOR2_X1 U805 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U806 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
XOR2_X1 U807 ( .A(n1144), .B(n1145), .Z(n1142) );
XOR2_X1 U808 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U809 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
XNOR2_X1 U810 ( .A(KEYINPUT40), .B(n1150), .ZN(n1148) );
XOR2_X1 U811 ( .A(KEYINPUT41), .B(KEYINPUT22), .Z(n1144) );
NOR2_X1 U812 ( .A1(n1151), .A2(n1152), .ZN(G66) );
NOR3_X1 U813 ( .A1(n1107), .A2(n1153), .A3(n1154), .ZN(n1152) );
AND3_X1 U814 ( .A1(n1155), .A2(n1109), .A3(n1156), .ZN(n1154) );
NOR2_X1 U815 ( .A1(n1157), .A2(n1155), .ZN(n1153) );
NOR2_X1 U816 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U817 ( .A1(n1151), .A2(n1160), .ZN(G63) );
XOR2_X1 U818 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U819 ( .A1(n1156), .A2(G478), .ZN(n1161) );
NOR2_X1 U820 ( .A1(n1151), .A2(n1163), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
NOR4_X1 U822 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U823 ( .A1(n1171), .A2(n1172), .ZN(n1164) );
NOR2_X1 U824 ( .A1(n1167), .A2(n1168), .ZN(n1172) );
NOR2_X1 U825 ( .A1(n1158), .A2(n1169), .ZN(n1171) );
INV_X1 U826 ( .A(G475), .ZN(n1169) );
XOR2_X1 U827 ( .A(G104), .B(n1173), .Z(G6) );
AND3_X1 U828 ( .A1(n1174), .A2(n1050), .A3(n1085), .ZN(n1173) );
NOR2_X1 U829 ( .A1(n1151), .A2(n1175), .ZN(G57) );
XOR2_X1 U830 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U831 ( .A1(n1156), .A2(G472), .ZN(n1176) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1178), .ZN(G54) );
XOR2_X1 U833 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U834 ( .A(n1181), .B(n1182), .Z(n1179) );
NOR2_X1 U835 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND3_X1 U836 ( .A1(G469), .A2(n1060), .A3(n1185), .ZN(n1181) );
XOR2_X1 U837 ( .A(n1186), .B(KEYINPUT30), .Z(n1185) );
NOR2_X1 U838 ( .A1(n1151), .A2(n1187), .ZN(G51) );
XOR2_X1 U839 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U840 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U841 ( .A1(n1156), .A2(n1192), .ZN(n1191) );
INV_X1 U842 ( .A(n1170), .ZN(n1156) );
NAND2_X1 U843 ( .A1(G902), .A2(n1060), .ZN(n1170) );
INV_X1 U844 ( .A(n1158), .ZN(n1060) );
NOR3_X1 U845 ( .A1(n1141), .A2(n1193), .A3(n1129), .ZN(n1158) );
NAND4_X1 U846 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1129) );
NOR4_X1 U847 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NOR2_X1 U848 ( .A1(KEYINPUT57), .A2(n1202), .ZN(n1201) );
NOR3_X1 U849 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1196) );
NOR4_X1 U850 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1076), .ZN(n1205) );
NAND2_X1 U851 ( .A1(n1209), .A2(n1097), .ZN(n1207) );
INV_X1 U852 ( .A(KEYINPUT11), .ZN(n1206) );
NOR2_X1 U853 ( .A1(KEYINPUT11), .A2(n1210), .ZN(n1204) );
INV_X1 U854 ( .A(n1211), .ZN(n1203) );
NAND2_X1 U855 ( .A1(n1075), .A2(n1212), .ZN(n1194) );
NAND2_X1 U856 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND4_X1 U857 ( .A1(n1215), .A2(n1216), .A3(n1093), .A4(n1217), .ZN(n1213) );
AND2_X1 U858 ( .A1(n1096), .A2(KEYINPUT57), .ZN(n1217) );
XOR2_X1 U859 ( .A(KEYINPUT59), .B(n1218), .Z(n1193) );
NAND4_X1 U860 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1141) );
NOR4_X1 U861 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222) );
INV_X1 U862 ( .A(n1227), .ZN(n1226) );
INV_X1 U863 ( .A(n1228), .ZN(n1225) );
OR2_X1 U864 ( .A1(n1229), .A2(KEYINPUT0), .ZN(n1221) );
NAND3_X1 U865 ( .A1(n1050), .A2(n1230), .A3(n1174), .ZN(n1220) );
NAND2_X1 U866 ( .A1(n1054), .A2(n1231), .ZN(n1230) );
OR2_X1 U867 ( .A1(n1076), .A2(KEYINPUT3), .ZN(n1231) );
NAND3_X1 U868 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1219) );
NAND2_X1 U869 ( .A1(n1052), .A2(n1235), .ZN(n1233) );
NAND4_X1 U870 ( .A1(n1053), .A2(KEYINPUT3), .A3(n1085), .A4(n1050), .ZN(n1235) );
NAND2_X1 U871 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
NAND3_X1 U872 ( .A1(n1238), .A2(n1084), .A3(KEYINPUT0), .ZN(n1236) );
NAND2_X1 U873 ( .A1(n1239), .A2(KEYINPUT9), .ZN(n1190) );
XOR2_X1 U874 ( .A(n1240), .B(n1241), .Z(n1239) );
NOR3_X1 U875 ( .A1(n1242), .A2(KEYINPUT62), .A3(n1243), .ZN(n1241) );
NOR2_X1 U876 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
XNOR2_X1 U877 ( .A(KEYINPUT56), .B(n1246), .ZN(n1245) );
NOR2_X1 U878 ( .A1(n1091), .A2(G952), .ZN(n1151) );
XOR2_X1 U879 ( .A(n1247), .B(G146), .Z(G48) );
NAND2_X1 U880 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR3_X1 U881 ( .A1(n1214), .A2(n1085), .A3(KEYINPUT28), .ZN(n1249) );
NAND2_X1 U882 ( .A1(n1200), .A2(KEYINPUT28), .ZN(n1248) );
NOR2_X1 U883 ( .A1(n1214), .A2(n1076), .ZN(n1200) );
XOR2_X1 U884 ( .A(n1250), .B(n1195), .Z(G45) );
NAND3_X1 U885 ( .A1(n1096), .A2(n1251), .A3(n1252), .ZN(n1195) );
NOR3_X1 U886 ( .A1(n1237), .A2(n1253), .A3(n1099), .ZN(n1252) );
XOR2_X1 U887 ( .A(n1254), .B(n1255), .Z(G42) );
NOR2_X1 U888 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NOR3_X1 U889 ( .A1(n1258), .A2(n1259), .A3(n1065), .ZN(n1257) );
INV_X1 U890 ( .A(KEYINPUT5), .ZN(n1258) );
NOR2_X1 U891 ( .A1(KEYINPUT5), .A2(n1211), .ZN(n1256) );
NAND2_X1 U892 ( .A1(n1259), .A2(n1093), .ZN(n1211) );
AND3_X1 U893 ( .A1(n1251), .A2(n1085), .A3(n1097), .ZN(n1259) );
XNOR2_X1 U894 ( .A(n1199), .B(n1260), .ZN(G39) );
XOR2_X1 U895 ( .A(KEYINPUT8), .B(G137), .Z(n1260) );
AND3_X1 U896 ( .A1(n1251), .A2(n1093), .A3(n1238), .ZN(n1199) );
XNOR2_X1 U897 ( .A(G134), .B(n1202), .ZN(G36) );
NAND4_X1 U898 ( .A1(n1096), .A2(n1251), .A3(n1093), .A4(n1075), .ZN(n1202) );
XOR2_X1 U899 ( .A(n1198), .B(n1261), .Z(G33) );
NOR2_X1 U900 ( .A1(KEYINPUT24), .A2(n1262), .ZN(n1261) );
AND4_X1 U901 ( .A1(n1096), .A2(n1251), .A3(n1085), .A4(n1093), .ZN(n1198) );
INV_X1 U902 ( .A(n1065), .ZN(n1093) );
NAND2_X1 U903 ( .A1(n1263), .A2(n1089), .ZN(n1065) );
XOR2_X1 U904 ( .A(G128), .B(n1264), .Z(G30) );
NOR2_X1 U905 ( .A1(n1054), .A2(n1214), .ZN(n1264) );
NAND4_X1 U906 ( .A1(n1251), .A2(n1052), .A3(n1265), .A4(n1266), .ZN(n1214) );
INV_X1 U907 ( .A(n1237), .ZN(n1052) );
NOR2_X1 U908 ( .A1(n1216), .A2(n1053), .ZN(n1251) );
XOR2_X1 U909 ( .A(G101), .B(n1140), .Z(G3) );
INV_X1 U910 ( .A(n1218), .ZN(n1140) );
NAND3_X1 U911 ( .A1(n1080), .A2(n1096), .A3(n1174), .ZN(n1218) );
XNOR2_X1 U912 ( .A(G125), .B(n1210), .ZN(G27) );
NAND4_X1 U913 ( .A1(n1209), .A2(n1097), .A3(n1085), .A4(n1208), .ZN(n1210) );
INV_X1 U914 ( .A(n1216), .ZN(n1208) );
NAND2_X1 U915 ( .A1(n1267), .A2(n1268), .ZN(n1216) );
NAND2_X1 U916 ( .A1(n1123), .A2(n1269), .ZN(n1268) );
NAND2_X1 U917 ( .A1(n1270), .A2(n1132), .ZN(n1123) );
INV_X1 U918 ( .A(G900), .ZN(n1132) );
XOR2_X1 U919 ( .A(n1271), .B(G122), .Z(G24) );
NAND2_X1 U920 ( .A1(KEYINPUT2), .A2(n1227), .ZN(n1271) );
NAND4_X1 U921 ( .A1(n1272), .A2(n1050), .A3(n1273), .A4(n1117), .ZN(n1227) );
NOR2_X1 U922 ( .A1(n1266), .A2(n1265), .ZN(n1050) );
XOR2_X1 U923 ( .A(n1229), .B(n1274), .Z(G21) );
NAND2_X1 U924 ( .A1(KEYINPUT16), .A2(G119), .ZN(n1274) );
NAND2_X1 U925 ( .A1(n1272), .A2(n1238), .ZN(n1229) );
AND3_X1 U926 ( .A1(n1265), .A2(n1266), .A3(n1080), .ZN(n1238) );
INV_X1 U927 ( .A(n1275), .ZN(n1266) );
XOR2_X1 U928 ( .A(n1224), .B(n1276), .Z(G18) );
NOR2_X1 U929 ( .A1(KEYINPUT46), .A2(n1277), .ZN(n1276) );
XOR2_X1 U930 ( .A(KEYINPUT34), .B(G116), .Z(n1277) );
AND3_X1 U931 ( .A1(n1096), .A2(n1075), .A3(n1272), .ZN(n1224) );
INV_X1 U932 ( .A(n1054), .ZN(n1075) );
NAND2_X1 U933 ( .A1(n1278), .A2(n1273), .ZN(n1054) );
INV_X1 U934 ( .A(n1099), .ZN(n1273) );
XOR2_X1 U935 ( .A(G113), .B(n1223), .Z(G15) );
AND3_X1 U936 ( .A1(n1096), .A2(n1085), .A3(n1272), .ZN(n1223) );
AND2_X1 U937 ( .A1(n1209), .A2(n1234), .ZN(n1272) );
INV_X1 U938 ( .A(n1055), .ZN(n1234) );
NOR2_X1 U939 ( .A1(n1237), .A2(n1073), .ZN(n1209) );
INV_X1 U940 ( .A(n1076), .ZN(n1085) );
NAND2_X1 U941 ( .A1(n1099), .A2(n1279), .ZN(n1076) );
XOR2_X1 U942 ( .A(KEYINPUT60), .B(n1117), .Z(n1279) );
NOR2_X1 U943 ( .A1(n1265), .A2(n1275), .ZN(n1096) );
XOR2_X1 U944 ( .A(n1280), .B(n1228), .Z(G12) );
NAND3_X1 U945 ( .A1(n1097), .A2(n1080), .A3(n1174), .ZN(n1228) );
NOR3_X1 U946 ( .A1(n1055), .A2(n1053), .A3(n1237), .ZN(n1174) );
NAND2_X1 U947 ( .A1(n1088), .A2(n1089), .ZN(n1237) );
NAND2_X1 U948 ( .A1(G214), .A2(n1281), .ZN(n1089) );
INV_X1 U949 ( .A(n1263), .ZN(n1088) );
XOR2_X1 U950 ( .A(n1282), .B(n1192), .Z(n1263) );
AND2_X1 U951 ( .A1(G210), .A2(n1281), .ZN(n1192) );
NAND2_X1 U952 ( .A1(n1283), .A2(n1186), .ZN(n1281) );
NAND2_X1 U953 ( .A1(n1284), .A2(n1186), .ZN(n1282) );
XOR2_X1 U954 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U955 ( .A(n1240), .B(n1188), .ZN(n1286) );
XNOR2_X1 U956 ( .A(n1287), .B(n1288), .ZN(n1188) );
INV_X1 U957 ( .A(n1147), .ZN(n1288) );
XOR2_X1 U958 ( .A(n1289), .B(G122), .Z(n1147) );
NAND2_X1 U959 ( .A1(KEYINPUT32), .A2(n1280), .ZN(n1289) );
NAND2_X1 U960 ( .A1(n1149), .A2(n1150), .ZN(n1287) );
NAND2_X1 U961 ( .A1(n1290), .A2(n1291), .ZN(n1150) );
XNOR2_X1 U962 ( .A(n1292), .B(n1293), .ZN(n1291) );
XOR2_X1 U963 ( .A(G113), .B(n1294), .Z(n1290) );
NAND2_X1 U964 ( .A1(n1295), .A2(n1296), .ZN(n1149) );
XOR2_X1 U965 ( .A(n1293), .B(n1292), .Z(n1296) );
NOR2_X1 U966 ( .A1(KEYINPUT35), .A2(G101), .ZN(n1292) );
NAND2_X1 U967 ( .A1(n1297), .A2(n1298), .ZN(n1293) );
NAND2_X1 U968 ( .A1(G104), .A2(n1047), .ZN(n1298) );
XOR2_X1 U969 ( .A(n1299), .B(KEYINPUT12), .Z(n1297) );
NAND2_X1 U970 ( .A1(G107), .A2(n1300), .ZN(n1299) );
XOR2_X1 U971 ( .A(n1301), .B(n1294), .Z(n1295) );
NAND2_X1 U972 ( .A1(G224), .A2(n1091), .ZN(n1240) );
XOR2_X1 U973 ( .A(KEYINPUT42), .B(n1302), .Z(n1285) );
NOR2_X1 U974 ( .A1(n1303), .A2(n1243), .ZN(n1302) );
AND2_X1 U975 ( .A1(n1246), .A2(n1244), .ZN(n1243) );
NOR2_X1 U976 ( .A1(n1246), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U977 ( .A(KEYINPUT31), .B(n1244), .ZN(n1304) );
XNOR2_X1 U978 ( .A(G125), .B(KEYINPUT15), .ZN(n1244) );
XOR2_X1 U979 ( .A(n1305), .B(n1306), .Z(n1246) );
INV_X1 U980 ( .A(n1215), .ZN(n1053) );
NAND2_X1 U981 ( .A1(n1307), .A2(n1308), .ZN(n1215) );
OR2_X1 U982 ( .A1(n1073), .A2(KEYINPUT43), .ZN(n1308) );
INV_X1 U983 ( .A(n1084), .ZN(n1073) );
NOR2_X1 U984 ( .A1(n1079), .A2(n1103), .ZN(n1084) );
INV_X1 U985 ( .A(n1078), .ZN(n1103) );
NAND3_X1 U986 ( .A1(n1079), .A2(n1078), .A3(KEYINPUT43), .ZN(n1307) );
NAND2_X1 U987 ( .A1(G221), .A2(n1309), .ZN(n1078) );
XNOR2_X1 U988 ( .A(n1110), .B(G469), .ZN(n1079) );
NAND2_X1 U989 ( .A1(n1310), .A2(n1186), .ZN(n1110) );
XOR2_X1 U990 ( .A(n1311), .B(n1180), .Z(n1310) );
XNOR2_X1 U991 ( .A(n1312), .B(n1313), .ZN(n1180) );
XNOR2_X1 U992 ( .A(n1314), .B(n1128), .ZN(n1313) );
XNOR2_X1 U993 ( .A(n1315), .B(G143), .ZN(n1128) );
XNOR2_X1 U994 ( .A(KEYINPUT38), .B(KEYINPUT10), .ZN(n1315) );
NAND2_X1 U995 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
OR2_X1 U996 ( .A1(n1318), .A2(G107), .ZN(n1317) );
XOR2_X1 U997 ( .A(n1319), .B(KEYINPUT63), .Z(n1316) );
NAND2_X1 U998 ( .A1(G107), .A2(n1318), .ZN(n1319) );
XNOR2_X1 U999 ( .A(n1300), .B(KEYINPUT27), .ZN(n1318) );
INV_X1 U1000 ( .A(G104), .ZN(n1300) );
NOR3_X1 U1001 ( .A1(n1184), .A2(n1320), .A3(n1321), .ZN(n1311) );
AND2_X1 U1002 ( .A1(KEYINPUT1), .A2(n1183), .ZN(n1321) );
AND2_X1 U1003 ( .A1(n1322), .A2(n1323), .ZN(n1183) );
NOR2_X1 U1004 ( .A1(KEYINPUT1), .A2(n1323), .ZN(n1320) );
NOR2_X1 U1005 ( .A1(n1323), .A2(n1322), .ZN(n1184) );
NOR2_X1 U1006 ( .A1(n1131), .A2(G953), .ZN(n1322) );
INV_X1 U1007 ( .A(G227), .ZN(n1131) );
XOR2_X1 U1008 ( .A(G110), .B(n1254), .Z(n1323) );
NAND2_X1 U1009 ( .A1(n1267), .A2(n1324), .ZN(n1055) );
NAND2_X1 U1010 ( .A1(n1143), .A2(n1269), .ZN(n1324) );
NAND2_X1 U1011 ( .A1(n1270), .A2(n1325), .ZN(n1143) );
INV_X1 U1012 ( .A(G898), .ZN(n1325) );
XOR2_X1 U1013 ( .A(G953), .B(KEYINPUT53), .Z(n1270) );
AND2_X1 U1014 ( .A1(n1083), .A2(n1326), .ZN(n1267) );
NAND2_X1 U1015 ( .A1(n1269), .A2(n1186), .ZN(n1326) );
NAND2_X1 U1016 ( .A1(n1327), .A2(n1091), .ZN(n1269) );
XNOR2_X1 U1017 ( .A(G952), .B(KEYINPUT37), .ZN(n1327) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1083) );
INV_X1 U1019 ( .A(n1081), .ZN(n1080) );
NAND2_X1 U1020 ( .A1(n1099), .A2(n1278), .ZN(n1081) );
XOR2_X1 U1021 ( .A(n1253), .B(KEYINPUT14), .Z(n1278) );
INV_X1 U1022 ( .A(n1117), .ZN(n1253) );
XOR2_X1 U1023 ( .A(n1165), .B(G475), .Z(n1117) );
AND2_X1 U1024 ( .A1(n1328), .A2(n1186), .ZN(n1165) );
OR2_X1 U1025 ( .A1(n1168), .A2(n1167), .ZN(n1328) );
AND2_X1 U1026 ( .A1(n1329), .A2(n1330), .ZN(n1167) );
XNOR2_X1 U1027 ( .A(n1331), .B(KEYINPUT36), .ZN(n1168) );
OR2_X1 U1028 ( .A1(n1330), .A2(n1329), .ZN(n1331) );
XNOR2_X1 U1029 ( .A(n1332), .B(G104), .ZN(n1329) );
NAND2_X1 U1030 ( .A1(KEYINPUT50), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1031 ( .A(G122), .B(G113), .Z(n1333) );
XNOR2_X1 U1032 ( .A(n1334), .B(n1127), .ZN(n1330) );
XOR2_X1 U1033 ( .A(G125), .B(G140), .Z(n1127) );
XNOR2_X1 U1034 ( .A(n1335), .B(n1336), .ZN(n1334) );
NOR2_X1 U1035 ( .A1(G146), .A2(KEYINPUT29), .ZN(n1336) );
NOR2_X1 U1036 ( .A1(KEYINPUT6), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1037 ( .A(n1338), .B(G131), .Z(n1337) );
NAND2_X1 U1038 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND4_X1 U1039 ( .A1(G143), .A2(G214), .A3(n1283), .A4(n1091), .ZN(n1340) );
XOR2_X1 U1040 ( .A(n1341), .B(KEYINPUT55), .Z(n1339) );
NAND2_X1 U1041 ( .A1(n1250), .A2(n1342), .ZN(n1341) );
NAND3_X1 U1042 ( .A1(n1283), .A2(n1091), .A3(G214), .ZN(n1342) );
XOR2_X1 U1043 ( .A(n1343), .B(G478), .Z(n1099) );
NAND2_X1 U1044 ( .A1(n1162), .A2(n1186), .ZN(n1343) );
INV_X1 U1045 ( .A(G902), .ZN(n1186) );
XOR2_X1 U1046 ( .A(n1344), .B(n1345), .Z(n1162) );
AND2_X1 U1047 ( .A1(n1346), .A2(G217), .ZN(n1345) );
NAND3_X1 U1048 ( .A1(KEYINPUT25), .A2(n1347), .A3(n1348), .ZN(n1344) );
XOR2_X1 U1049 ( .A(n1349), .B(KEYINPUT58), .Z(n1348) );
OR2_X1 U1050 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1051 ( .A1(n1351), .A2(n1350), .ZN(n1347) );
XOR2_X1 U1052 ( .A(G134), .B(n1352), .Z(n1350) );
NOR2_X1 U1053 ( .A1(KEYINPUT23), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1054 ( .A(G143), .B(G128), .Z(n1353) );
XNOR2_X1 U1055 ( .A(n1047), .B(n1354), .ZN(n1351) );
XOR2_X1 U1056 ( .A(G122), .B(G116), .Z(n1354) );
INV_X1 U1057 ( .A(G107), .ZN(n1047) );
AND2_X1 U1058 ( .A1(n1275), .A2(n1265), .ZN(n1097) );
XOR2_X1 U1059 ( .A(n1107), .B(n1109), .Z(n1265) );
INV_X1 U1060 ( .A(n1159), .ZN(n1109) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1309), .ZN(n1159) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1355), .ZN(n1309) );
XOR2_X1 U1063 ( .A(KEYINPUT48), .B(G902), .Z(n1355) );
NOR2_X1 U1064 ( .A1(n1155), .A2(G902), .ZN(n1107) );
XNOR2_X1 U1065 ( .A(n1356), .B(n1357), .ZN(n1155) );
XOR2_X1 U1066 ( .A(n1358), .B(n1359), .Z(n1357) );
NAND2_X1 U1067 ( .A1(G221), .A2(n1346), .ZN(n1359) );
AND2_X1 U1068 ( .A1(G234), .A2(n1091), .ZN(n1346) );
NAND2_X1 U1069 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
OR2_X1 U1070 ( .A1(n1254), .A2(G125), .ZN(n1361) );
XOR2_X1 U1071 ( .A(n1362), .B(KEYINPUT47), .Z(n1360) );
NAND2_X1 U1072 ( .A1(G125), .A2(n1254), .ZN(n1362) );
INV_X1 U1073 ( .A(G140), .ZN(n1254) );
XOR2_X1 U1074 ( .A(n1363), .B(n1364), .Z(n1356) );
NOR2_X1 U1075 ( .A1(KEYINPUT51), .A2(n1365), .ZN(n1364) );
XOR2_X1 U1076 ( .A(n1366), .B(n1367), .Z(n1365) );
NOR2_X1 U1077 ( .A1(G110), .A2(KEYINPUT21), .ZN(n1367) );
XOR2_X1 U1078 ( .A(n1368), .B(n1369), .Z(n1366) );
NOR2_X1 U1079 ( .A1(G119), .A2(KEYINPUT44), .ZN(n1369) );
INV_X1 U1080 ( .A(G128), .ZN(n1368) );
XOR2_X1 U1081 ( .A(n1370), .B(G146), .Z(n1363) );
INV_X1 U1082 ( .A(G137), .ZN(n1370) );
NOR2_X1 U1083 ( .A1(n1371), .A2(n1116), .ZN(n1275) );
NOR3_X1 U1084 ( .A1(G472), .A2(G902), .A3(n1114), .ZN(n1116) );
AND2_X1 U1085 ( .A1(G472), .A2(n1372), .ZN(n1371) );
OR2_X1 U1086 ( .A1(n1114), .A2(G902), .ZN(n1372) );
XOR2_X1 U1087 ( .A(n1177), .B(n1373), .Z(n1114) );
XOR2_X1 U1088 ( .A(KEYINPUT45), .B(KEYINPUT18), .Z(n1373) );
XOR2_X1 U1089 ( .A(n1374), .B(n1375), .Z(n1177) );
XOR2_X1 U1090 ( .A(n1376), .B(n1377), .Z(n1375) );
XOR2_X1 U1091 ( .A(n1305), .B(n1378), .Z(n1377) );
NAND2_X1 U1092 ( .A1(KEYINPUT19), .A2(n1301), .ZN(n1378) );
INV_X1 U1093 ( .A(G113), .ZN(n1301) );
NAND2_X1 U1094 ( .A1(KEYINPUT13), .A2(n1250), .ZN(n1305) );
INV_X1 U1095 ( .A(G143), .ZN(n1250) );
AND3_X1 U1096 ( .A1(G210), .A2(n1091), .A3(n1283), .ZN(n1376) );
INV_X1 U1097 ( .A(G237), .ZN(n1283) );
INV_X1 U1098 ( .A(G953), .ZN(n1091) );
XOR2_X1 U1099 ( .A(n1312), .B(n1294), .Z(n1374) );
XOR2_X1 U1100 ( .A(G116), .B(G119), .Z(n1294) );
XOR2_X1 U1101 ( .A(n1126), .B(n1379), .Z(n1312) );
XOR2_X1 U1102 ( .A(KEYINPUT54), .B(G101), .Z(n1379) );
XOR2_X1 U1103 ( .A(n1380), .B(n1381), .Z(n1126) );
XOR2_X1 U1104 ( .A(G134), .B(n1382), .Z(n1381) );
XOR2_X1 U1105 ( .A(KEYINPUT33), .B(G137), .Z(n1382) );
XOR2_X1 U1106 ( .A(n1262), .B(n1306), .Z(n1380) );
XOR2_X1 U1107 ( .A(G128), .B(G146), .Z(n1306) );
INV_X1 U1108 ( .A(G131), .ZN(n1262) );
INV_X1 U1109 ( .A(G110), .ZN(n1280) );
endmodule


