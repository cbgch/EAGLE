//Key = 1111111111101001101101110100111001110100111110111001000010010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314;

XOR2_X1 U738 ( .A(n1008), .B(n1009), .Z(G9) );
NOR2_X1 U739 ( .A1(G107), .A2(KEYINPUT53), .ZN(n1009) );
NOR2_X1 U740 ( .A1(n1010), .A2(n1011), .ZN(G75) );
XOR2_X1 U741 ( .A(n1012), .B(KEYINPUT15), .Z(n1011) );
NAND3_X1 U742 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NAND2_X1 U743 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U744 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND3_X1 U745 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NAND2_X1 U746 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NAND2_X1 U747 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
OR2_X1 U748 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U749 ( .A1(n1029), .A2(n1030), .ZN(n1023) );
NAND2_X1 U750 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U751 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND3_X1 U752 ( .A1(n1025), .A2(n1035), .A3(n1029), .ZN(n1018) );
NAND2_X1 U753 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U754 ( .A1(n1022), .A2(n1038), .ZN(n1037) );
NAND2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U756 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U757 ( .A1(n1020), .A2(n1043), .ZN(n1036) );
NAND3_X1 U758 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U759 ( .A1(n1022), .A2(n1047), .ZN(n1045) );
OR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1047), .ZN(n1044) );
INV_X1 U761 ( .A(KEYINPUT43), .ZN(n1047) );
INV_X1 U762 ( .A(n1050), .ZN(n1016) );
INV_X1 U763 ( .A(n1051), .ZN(n1013) );
NOR2_X1 U764 ( .A1(G952), .A2(n1051), .ZN(n1010) );
NAND2_X1 U765 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND4_X1 U766 ( .A1(n1054), .A2(n1055), .A3(n1022), .A4(n1056), .ZN(n1053) );
NOR3_X1 U767 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
XNOR2_X1 U768 ( .A(G472), .B(n1060), .ZN(n1059) );
XOR2_X1 U769 ( .A(n1061), .B(n1062), .Z(n1057) );
XNOR2_X1 U770 ( .A(n1063), .B(KEYINPUT9), .ZN(n1062) );
NAND2_X1 U771 ( .A1(KEYINPUT4), .A2(n1064), .ZN(n1061) );
INV_X1 U772 ( .A(n1042), .ZN(n1055) );
XOR2_X1 U773 ( .A(n1065), .B(n1066), .Z(G72) );
XOR2_X1 U774 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U775 ( .A1(n1069), .A2(G953), .ZN(n1068) );
NOR2_X1 U776 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
XOR2_X1 U777 ( .A(n1072), .B(n1073), .Z(n1071) );
XNOR2_X1 U778 ( .A(KEYINPUT56), .B(n1074), .ZN(n1073) );
XOR2_X1 U779 ( .A(n1075), .B(n1076), .Z(n1072) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U781 ( .A(n1079), .B(KEYINPUT48), .Z(n1078) );
NAND2_X1 U782 ( .A1(G131), .A2(n1080), .ZN(n1079) );
NOR2_X1 U783 ( .A1(G131), .A2(n1080), .ZN(n1077) );
XOR2_X1 U784 ( .A(G137), .B(G134), .Z(n1080) );
NOR2_X1 U785 ( .A1(G900), .A2(n1081), .ZN(n1070) );
XNOR2_X1 U786 ( .A(KEYINPUT35), .B(n1052), .ZN(n1081) );
NOR2_X1 U787 ( .A1(n1082), .A2(n1052), .ZN(n1065) );
NOR2_X1 U788 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U789 ( .A(n1085), .B(n1086), .Z(G69) );
NOR2_X1 U790 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U791 ( .A1(G224), .A2(n1052), .ZN(n1087) );
NOR3_X1 U792 ( .A1(KEYINPUT50), .A2(n1089), .A3(n1090), .ZN(n1085) );
NOR3_X1 U793 ( .A1(n1091), .A2(n1088), .A3(n1092), .ZN(n1090) );
XOR2_X1 U794 ( .A(n1093), .B(KEYINPUT16), .Z(n1092) );
NOR2_X1 U795 ( .A1(n1094), .A2(n1093), .ZN(n1089) );
NAND2_X1 U796 ( .A1(n1052), .A2(n1095), .ZN(n1093) );
NAND2_X1 U797 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
INV_X1 U798 ( .A(n1091), .ZN(n1094) );
XOR2_X1 U799 ( .A(n1098), .B(n1099), .Z(n1091) );
NOR3_X1 U800 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(G66) );
NOR4_X1 U801 ( .A1(n1103), .A2(n1104), .A3(KEYINPUT58), .A4(n1105), .ZN(n1102) );
NOR2_X1 U802 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NOR3_X1 U803 ( .A1(n1104), .A2(n1108), .A3(n1105), .ZN(n1107) );
NOR2_X1 U804 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U805 ( .A(KEYINPUT58), .ZN(n1110) );
INV_X1 U806 ( .A(n1103), .ZN(n1106) );
NAND2_X1 U807 ( .A1(n1109), .A2(KEYINPUT3), .ZN(n1103) );
XNOR2_X1 U808 ( .A(n1111), .B(KEYINPUT30), .ZN(n1109) );
NOR2_X1 U809 ( .A1(n1100), .A2(n1112), .ZN(G63) );
NOR3_X1 U810 ( .A1(n1063), .A2(n1113), .A3(n1114), .ZN(n1112) );
AND3_X1 U811 ( .A1(n1115), .A2(G478), .A3(n1116), .ZN(n1114) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1115), .ZN(n1113) );
NOR2_X1 U813 ( .A1(n1015), .A2(n1064), .ZN(n1117) );
NOR2_X1 U814 ( .A1(n1100), .A2(n1118), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1119), .B(n1120), .ZN(n1118) );
AND2_X1 U816 ( .A1(G475), .A2(n1116), .ZN(n1120) );
XNOR2_X1 U817 ( .A(G104), .B(n1097), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1121), .A2(n1122), .ZN(G57) );
XOR2_X1 U819 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U820 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U821 ( .A1(KEYINPUT17), .A2(n1127), .ZN(n1126) );
NAND2_X1 U822 ( .A1(KEYINPUT1), .A2(n1128), .ZN(n1125) );
NAND2_X1 U823 ( .A1(n1116), .A2(G472), .ZN(n1128) );
XOR2_X1 U824 ( .A(n1129), .B(n1130), .Z(n1123) );
NOR2_X1 U825 ( .A1(G952), .A2(n1131), .ZN(n1121) );
XNOR2_X1 U826 ( .A(G953), .B(KEYINPUT24), .ZN(n1131) );
NOR2_X1 U827 ( .A1(n1100), .A2(n1132), .ZN(G54) );
XOR2_X1 U828 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U829 ( .A(KEYINPUT10), .B(n1135), .Z(n1134) );
AND2_X1 U830 ( .A1(G469), .A2(n1116), .ZN(n1135) );
NOR2_X1 U831 ( .A1(n1100), .A2(n1136), .ZN(G51) );
XOR2_X1 U832 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U833 ( .A1(n1139), .A2(n1104), .ZN(n1138) );
INV_X1 U834 ( .A(n1116), .ZN(n1104) );
NOR2_X1 U835 ( .A1(n1140), .A2(n1015), .ZN(n1116) );
AND3_X1 U836 ( .A1(n1096), .A2(n1141), .A3(n1069), .ZN(n1015) );
AND4_X1 U837 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1069) );
NOR4_X1 U838 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
AND2_X1 U839 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U840 ( .A1(n1152), .A2(n1153), .ZN(n1142) );
XNOR2_X1 U841 ( .A(KEYINPUT60), .B(n1154), .ZN(n1152) );
XNOR2_X1 U842 ( .A(KEYINPUT34), .B(n1097), .ZN(n1141) );
NAND3_X1 U843 ( .A1(n1155), .A2(n1020), .A3(n1027), .ZN(n1097) );
AND4_X1 U844 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1096) );
AND4_X1 U845 ( .A1(n1008), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1159) );
NAND3_X1 U846 ( .A1(n1028), .A2(n1020), .A3(n1155), .ZN(n1008) );
NAND3_X1 U847 ( .A1(n1163), .A2(n1028), .A3(n1164), .ZN(n1158) );
XOR2_X1 U848 ( .A(n1165), .B(n1166), .Z(n1137) );
NOR2_X1 U849 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U850 ( .A(n1169), .B(KEYINPUT46), .Z(n1168) );
INV_X1 U851 ( .A(n1170), .ZN(n1167) );
NOR2_X1 U852 ( .A1(n1052), .A2(G952), .ZN(n1100) );
XOR2_X1 U853 ( .A(n1171), .B(n1149), .Z(G48) );
AND4_X1 U854 ( .A1(n1027), .A2(n1172), .A3(n1153), .A4(n1173), .ZN(n1149) );
NAND2_X1 U855 ( .A1(KEYINPUT23), .A2(n1174), .ZN(n1171) );
XNOR2_X1 U856 ( .A(G143), .B(n1143), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1175), .A2(n1153), .A3(n1176), .A4(n1177), .ZN(n1143) );
XNOR2_X1 U858 ( .A(G140), .B(n1151), .ZN(G42) );
NAND4_X1 U859 ( .A1(n1027), .A2(n1172), .A3(n1022), .A4(n1041), .ZN(n1151) );
XNOR2_X1 U860 ( .A(G137), .B(n1150), .ZN(G39) );
NAND4_X1 U861 ( .A1(n1029), .A2(n1172), .A3(n1022), .A4(n1173), .ZN(n1150) );
XOR2_X1 U862 ( .A(n1148), .B(n1178), .Z(G36) );
NOR2_X1 U863 ( .A1(KEYINPUT55), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U864 ( .A(G134), .B(KEYINPUT45), .ZN(n1179) );
AND3_X1 U865 ( .A1(n1022), .A2(n1028), .A3(n1175), .ZN(n1148) );
XOR2_X1 U866 ( .A(G131), .B(n1147), .Z(G33) );
AND3_X1 U867 ( .A1(n1175), .A2(n1022), .A3(n1027), .ZN(n1147) );
NOR2_X1 U868 ( .A1(n1049), .A2(n1180), .ZN(n1022) );
AND3_X1 U869 ( .A1(n1181), .A2(n1182), .A3(n1163), .ZN(n1175) );
XNOR2_X1 U870 ( .A(n1146), .B(n1183), .ZN(G30) );
NOR2_X1 U871 ( .A1(G128), .A2(KEYINPUT27), .ZN(n1183) );
AND4_X1 U872 ( .A1(n1172), .A2(n1028), .A3(n1153), .A4(n1173), .ZN(n1146) );
AND3_X1 U873 ( .A1(n1042), .A2(n1182), .A3(n1181), .ZN(n1172) );
XNOR2_X1 U874 ( .A(G101), .B(n1156), .ZN(G3) );
NAND3_X1 U875 ( .A1(n1163), .A2(n1155), .A3(n1029), .ZN(n1156) );
XNOR2_X1 U876 ( .A(n1074), .B(n1184), .ZN(G27) );
NOR2_X1 U877 ( .A1(n1046), .A2(n1154), .ZN(n1184) );
NAND4_X1 U878 ( .A1(n1027), .A2(n1025), .A3(n1185), .A4(n1041), .ZN(n1154) );
AND2_X1 U879 ( .A1(n1182), .A2(n1042), .ZN(n1185) );
NAND2_X1 U880 ( .A1(n1050), .A2(n1186), .ZN(n1182) );
NAND4_X1 U881 ( .A1(G902), .A2(G953), .A3(n1187), .A4(n1084), .ZN(n1186) );
INV_X1 U882 ( .A(G900), .ZN(n1084) );
INV_X1 U883 ( .A(n1058), .ZN(n1025) );
XNOR2_X1 U884 ( .A(G122), .B(n1157), .ZN(G24) );
NAND4_X1 U885 ( .A1(n1164), .A2(n1020), .A3(n1176), .A4(n1177), .ZN(n1157) );
NOR2_X1 U886 ( .A1(n1173), .A2(n1042), .ZN(n1020) );
XNOR2_X1 U887 ( .A(G119), .B(n1162), .ZN(G21) );
NAND4_X1 U888 ( .A1(n1164), .A2(n1029), .A3(n1042), .A4(n1173), .ZN(n1162) );
XNOR2_X1 U889 ( .A(G116), .B(n1188), .ZN(G18) );
NOR2_X1 U890 ( .A1(KEYINPUT32), .A2(n1189), .ZN(n1188) );
NOR3_X1 U891 ( .A1(n1190), .A2(n1039), .A3(n1191), .ZN(n1189) );
INV_X1 U892 ( .A(n1164), .ZN(n1191) );
NOR3_X1 U893 ( .A1(n1046), .A2(n1192), .A3(n1058), .ZN(n1164) );
INV_X1 U894 ( .A(n1153), .ZN(n1046) );
XNOR2_X1 U895 ( .A(n1193), .B(KEYINPUT14), .ZN(n1153) );
INV_X1 U896 ( .A(n1163), .ZN(n1039) );
XOR2_X1 U897 ( .A(KEYINPUT18), .B(n1028), .Z(n1190) );
AND2_X1 U898 ( .A1(n1054), .A2(n1176), .ZN(n1028) );
XNOR2_X1 U899 ( .A(G113), .B(n1161), .ZN(G15) );
NAND3_X1 U900 ( .A1(n1027), .A2(n1163), .A3(n1194), .ZN(n1161) );
NOR3_X1 U901 ( .A1(n1058), .A2(n1192), .A3(n1193), .ZN(n1194) );
NAND2_X1 U902 ( .A1(n1034), .A2(n1195), .ZN(n1058) );
NOR2_X1 U903 ( .A1(n1042), .A2(n1041), .ZN(n1163) );
NOR2_X1 U904 ( .A1(n1176), .A2(n1054), .ZN(n1027) );
INV_X1 U905 ( .A(n1177), .ZN(n1054) );
NAND3_X1 U906 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(G12) );
OR2_X1 U907 ( .A1(n1199), .A2(KEYINPUT62), .ZN(n1198) );
NAND3_X1 U908 ( .A1(KEYINPUT62), .A2(n1199), .A3(n1200), .ZN(n1197) );
NAND2_X1 U909 ( .A1(G110), .A2(n1201), .ZN(n1196) );
NAND2_X1 U910 ( .A1(n1202), .A2(KEYINPUT62), .ZN(n1201) );
XNOR2_X1 U911 ( .A(n1199), .B(KEYINPUT51), .ZN(n1202) );
INV_X1 U912 ( .A(n1160), .ZN(n1199) );
NAND4_X1 U913 ( .A1(n1029), .A2(n1155), .A3(n1041), .A4(n1042), .ZN(n1160) );
XOR2_X1 U914 ( .A(n1203), .B(n1105), .Z(n1042) );
NAND2_X1 U915 ( .A1(G217), .A2(n1204), .ZN(n1105) );
NAND2_X1 U916 ( .A1(n1111), .A2(n1140), .ZN(n1203) );
XNOR2_X1 U917 ( .A(n1205), .B(n1206), .ZN(n1111) );
XOR2_X1 U918 ( .A(KEYINPUT7), .B(G137), .Z(n1206) );
XOR2_X1 U919 ( .A(n1207), .B(n1208), .Z(n1205) );
AND2_X1 U920 ( .A1(G221), .A2(n1209), .ZN(n1208) );
NAND2_X1 U921 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
NAND2_X1 U922 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U923 ( .A(KEYINPUT37), .B(n1214), .Z(n1210) );
NOR2_X1 U924 ( .A1(n1212), .A2(n1213), .ZN(n1214) );
NAND3_X1 U925 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1213) );
NAND2_X1 U926 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U927 ( .A(KEYINPUT0), .ZN(n1219) );
NAND3_X1 U928 ( .A1(KEYINPUT0), .A2(n1220), .A3(n1174), .ZN(n1216) );
OR2_X1 U929 ( .A1(n1174), .A2(n1220), .ZN(n1215) );
NOR2_X1 U930 ( .A1(KEYINPUT39), .A2(n1218), .ZN(n1220) );
XOR2_X1 U931 ( .A(n1221), .B(n1222), .Z(n1218) );
NAND2_X1 U932 ( .A1(KEYINPUT6), .A2(n1074), .ZN(n1221) );
XNOR2_X1 U933 ( .A(n1223), .B(n1224), .ZN(n1212) );
XOR2_X1 U934 ( .A(KEYINPUT38), .B(G128), .Z(n1224) );
XNOR2_X1 U935 ( .A(n1225), .B(n1226), .ZN(n1223) );
NOR2_X1 U936 ( .A1(KEYINPUT31), .A2(n1200), .ZN(n1226) );
INV_X1 U937 ( .A(G110), .ZN(n1200) );
NOR2_X1 U938 ( .A1(G119), .A2(KEYINPUT36), .ZN(n1225) );
INV_X1 U939 ( .A(n1173), .ZN(n1041) );
NAND2_X1 U940 ( .A1(n1227), .A2(n1228), .ZN(n1173) );
NAND2_X1 U941 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XOR2_X1 U942 ( .A(KEYINPUT25), .B(n1231), .Z(n1227) );
NOR2_X1 U943 ( .A1(n1229), .A2(n1230), .ZN(n1231) );
INV_X1 U944 ( .A(G472), .ZN(n1230) );
INV_X1 U945 ( .A(n1060), .ZN(n1229) );
NAND2_X1 U946 ( .A1(n1232), .A2(n1140), .ZN(n1060) );
XOR2_X1 U947 ( .A(n1233), .B(n1129), .Z(n1232) );
XOR2_X1 U948 ( .A(n1234), .B(G101), .Z(n1129) );
NAND3_X1 U949 ( .A1(n1235), .A2(n1052), .A3(G210), .ZN(n1234) );
XNOR2_X1 U950 ( .A(KEYINPUT12), .B(n1236), .ZN(n1235) );
NAND2_X1 U951 ( .A1(n1237), .A2(n1238), .ZN(n1233) );
NAND2_X1 U952 ( .A1(n1127), .A2(n1130), .ZN(n1238) );
XOR2_X1 U953 ( .A(KEYINPUT59), .B(n1239), .Z(n1237) );
NOR2_X1 U954 ( .A1(n1127), .A2(n1130), .ZN(n1239) );
XNOR2_X1 U955 ( .A(n1240), .B(n1241), .ZN(n1130) );
XNOR2_X1 U956 ( .A(n1242), .B(n1243), .ZN(n1127) );
NAND2_X1 U957 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
NAND2_X1 U958 ( .A1(G119), .A2(n1246), .ZN(n1245) );
XOR2_X1 U959 ( .A(KEYINPUT41), .B(n1247), .Z(n1244) );
NOR2_X1 U960 ( .A1(G119), .A2(n1246), .ZN(n1247) );
INV_X1 U961 ( .A(G116), .ZN(n1246) );
NOR3_X1 U962 ( .A1(n1193), .A2(n1192), .A3(n1031), .ZN(n1155) );
INV_X1 U963 ( .A(n1181), .ZN(n1031) );
NOR2_X1 U964 ( .A1(n1034), .A2(n1033), .ZN(n1181) );
INV_X1 U965 ( .A(n1195), .ZN(n1033) );
NAND2_X1 U966 ( .A1(G221), .A2(n1204), .ZN(n1195) );
NAND2_X1 U967 ( .A1(G234), .A2(n1140), .ZN(n1204) );
XOR2_X1 U968 ( .A(n1248), .B(G469), .Z(n1034) );
NAND2_X1 U969 ( .A1(n1133), .A2(n1140), .ZN(n1248) );
XOR2_X1 U970 ( .A(n1249), .B(n1250), .Z(n1133) );
XNOR2_X1 U971 ( .A(n1241), .B(n1251), .ZN(n1250) );
XNOR2_X1 U972 ( .A(G110), .B(n1252), .ZN(n1251) );
NOR2_X1 U973 ( .A1(G953), .A2(n1083), .ZN(n1252) );
INV_X1 U974 ( .A(G227), .ZN(n1083) );
XNOR2_X1 U975 ( .A(n1253), .B(n1254), .ZN(n1241) );
XOR2_X1 U976 ( .A(G134), .B(G131), .Z(n1254) );
NAND2_X1 U977 ( .A1(KEYINPUT21), .A2(n1255), .ZN(n1253) );
XOR2_X1 U978 ( .A(KEYINPUT5), .B(G137), .Z(n1255) );
XOR2_X1 U979 ( .A(n1075), .B(n1256), .Z(n1249) );
XOR2_X1 U980 ( .A(n1257), .B(n1258), .Z(n1075) );
XOR2_X1 U981 ( .A(G140), .B(G128), .Z(n1258) );
XNOR2_X1 U982 ( .A(G143), .B(n1259), .ZN(n1257) );
XNOR2_X1 U983 ( .A(KEYINPUT54), .B(n1174), .ZN(n1259) );
AND2_X1 U984 ( .A1(n1050), .A2(n1260), .ZN(n1192) );
NAND3_X1 U985 ( .A1(n1088), .A2(n1187), .A3(G902), .ZN(n1260) );
NOR2_X1 U986 ( .A1(G898), .A2(n1052), .ZN(n1088) );
NAND3_X1 U987 ( .A1(n1187), .A2(n1052), .A3(G952), .ZN(n1050) );
NAND2_X1 U988 ( .A1(G237), .A2(G234), .ZN(n1187) );
NAND2_X1 U989 ( .A1(n1261), .A2(n1049), .ZN(n1193) );
XNOR2_X1 U990 ( .A(n1139), .B(n1262), .ZN(n1049) );
NOR2_X1 U991 ( .A1(G902), .A2(n1263), .ZN(n1262) );
XOR2_X1 U992 ( .A(n1165), .B(n1264), .Z(n1263) );
NAND2_X1 U993 ( .A1(KEYINPUT33), .A2(n1265), .ZN(n1264) );
NAND2_X1 U994 ( .A1(n1169), .A2(n1170), .ZN(n1265) );
NAND3_X1 U995 ( .A1(n1266), .A2(n1052), .A3(G224), .ZN(n1170) );
XNOR2_X1 U996 ( .A(G125), .B(n1240), .ZN(n1266) );
NAND2_X1 U997 ( .A1(n1267), .A2(n1268), .ZN(n1169) );
NAND2_X1 U998 ( .A1(G224), .A2(n1052), .ZN(n1268) );
XNOR2_X1 U999 ( .A(n1240), .B(n1074), .ZN(n1267) );
INV_X1 U1000 ( .A(G125), .ZN(n1074) );
XNOR2_X1 U1001 ( .A(n1269), .B(n1270), .ZN(n1240) );
NAND2_X1 U1002 ( .A1(KEYINPUT44), .A2(n1174), .ZN(n1269) );
INV_X1 U1003 ( .A(G146), .ZN(n1174) );
NAND3_X1 U1004 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1165) );
OR2_X1 U1005 ( .A1(n1098), .A2(KEYINPUT42), .ZN(n1273) );
NAND3_X1 U1006 ( .A1(KEYINPUT42), .A2(n1098), .A3(n1274), .ZN(n1272) );
NAND2_X1 U1007 ( .A1(n1099), .A2(n1275), .ZN(n1271) );
NAND2_X1 U1008 ( .A1(n1276), .A2(KEYINPUT42), .ZN(n1275) );
XNOR2_X1 U1009 ( .A(n1098), .B(KEYINPUT29), .ZN(n1276) );
XNOR2_X1 U1010 ( .A(n1277), .B(n1278), .ZN(n1098) );
XNOR2_X1 U1011 ( .A(G119), .B(n1279), .ZN(n1278) );
XNOR2_X1 U1012 ( .A(KEYINPUT40), .B(KEYINPUT2), .ZN(n1279) );
XNOR2_X1 U1013 ( .A(n1256), .B(n1280), .ZN(n1277) );
XNOR2_X1 U1014 ( .A(G116), .B(n1281), .ZN(n1280) );
NAND2_X1 U1015 ( .A1(KEYINPUT28), .A2(n1243), .ZN(n1281) );
XOR2_X1 U1016 ( .A(G101), .B(n1282), .Z(n1256) );
XOR2_X1 U1017 ( .A(G107), .B(G104), .Z(n1282) );
INV_X1 U1018 ( .A(n1274), .ZN(n1099) );
XOR2_X1 U1019 ( .A(G110), .B(G122), .Z(n1274) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1283), .ZN(n1139) );
XNOR2_X1 U1021 ( .A(n1180), .B(KEYINPUT20), .ZN(n1261) );
INV_X1 U1022 ( .A(n1048), .ZN(n1180) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1283), .ZN(n1048) );
NAND2_X1 U1024 ( .A1(n1236), .A2(n1140), .ZN(n1283) );
NOR2_X1 U1025 ( .A1(n1176), .A2(n1177), .ZN(n1029) );
XNOR2_X1 U1026 ( .A(n1284), .B(G475), .ZN(n1177) );
NAND2_X1 U1027 ( .A1(n1119), .A2(n1140), .ZN(n1284) );
INV_X1 U1028 ( .A(G902), .ZN(n1140) );
XNOR2_X1 U1029 ( .A(n1285), .B(n1286), .ZN(n1119) );
XNOR2_X1 U1030 ( .A(n1287), .B(n1288), .ZN(n1286) );
NOR2_X1 U1031 ( .A1(KEYINPUT11), .A2(n1289), .ZN(n1288) );
NOR3_X1 U1032 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
NOR2_X1 U1033 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NOR2_X1 U1034 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
INV_X1 U1035 ( .A(KEYINPUT47), .ZN(n1296) );
XNOR2_X1 U1036 ( .A(n1297), .B(KEYINPUT61), .ZN(n1295) );
AND3_X1 U1037 ( .A1(n1294), .A2(n1297), .A3(KEYINPUT47), .ZN(n1291) );
XOR2_X1 U1038 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U1039 ( .A(G143), .B(G131), .Z(n1299) );
NAND3_X1 U1040 ( .A1(n1236), .A2(n1052), .A3(G214), .ZN(n1298) );
INV_X1 U1041 ( .A(G237), .ZN(n1236) );
NOR2_X1 U1042 ( .A1(KEYINPUT47), .A2(n1297), .ZN(n1290) );
XNOR2_X1 U1043 ( .A(n1300), .B(n1222), .ZN(n1297) );
XOR2_X1 U1044 ( .A(G140), .B(KEYINPUT8), .Z(n1222) );
XNOR2_X1 U1045 ( .A(G125), .B(G146), .ZN(n1300) );
NAND2_X1 U1046 ( .A1(KEYINPUT19), .A2(n1243), .ZN(n1287) );
INV_X1 U1047 ( .A(G113), .ZN(n1243) );
XNOR2_X1 U1048 ( .A(G104), .B(n1301), .ZN(n1285) );
XOR2_X1 U1049 ( .A(KEYINPUT49), .B(G122), .Z(n1301) );
XOR2_X1 U1050 ( .A(n1063), .B(n1302), .Z(n1176) );
XNOR2_X1 U1051 ( .A(KEYINPUT57), .B(n1064), .ZN(n1302) );
INV_X1 U1052 ( .A(G478), .ZN(n1064) );
NOR2_X1 U1053 ( .A1(n1115), .A2(G902), .ZN(n1063) );
XOR2_X1 U1054 ( .A(n1303), .B(n1304), .Z(n1115) );
XOR2_X1 U1055 ( .A(G134), .B(n1305), .Z(n1304) );
NOR2_X1 U1056 ( .A1(KEYINPUT26), .A2(n1270), .ZN(n1305) );
XNOR2_X1 U1057 ( .A(G128), .B(G143), .ZN(n1270) );
XOR2_X1 U1058 ( .A(n1306), .B(n1307), .Z(n1303) );
NOR2_X1 U1059 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1060 ( .A(n1310), .B(KEYINPUT63), .Z(n1309) );
NAND2_X1 U1061 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1062 ( .A(KEYINPUT52), .B(n1313), .Z(n1312) );
NOR2_X1 U1063 ( .A1(n1311), .A2(n1313), .ZN(n1308) );
XOR2_X1 U1064 ( .A(G107), .B(KEYINPUT13), .Z(n1313) );
XNOR2_X1 U1065 ( .A(G116), .B(n1314), .ZN(n1311) );
XOR2_X1 U1066 ( .A(KEYINPUT22), .B(G122), .Z(n1314) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1209), .ZN(n1306) );
AND2_X1 U1068 ( .A1(G234), .A2(n1052), .ZN(n1209) );
INV_X1 U1069 ( .A(G953), .ZN(n1052) );
endmodule


