//Key = 1111101110111100011010111110001110110010001111100101010011100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;

XOR2_X1 U727 ( .A(G107), .B(n1011), .Z(G9) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U729 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
XOR2_X1 U730 ( .A(n1018), .B(KEYINPUT59), .Z(n1017) );
NAND2_X1 U731 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U732 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NAND3_X1 U733 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1019) );
NAND2_X1 U734 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND2_X1 U735 ( .A1(n1022), .A2(n1029), .ZN(n1028) );
NAND2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
XNOR2_X1 U738 ( .A(n1034), .B(KEYINPUT63), .ZN(n1032) );
NAND2_X1 U739 ( .A1(n1035), .A2(n1036), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1037), .A2(n1035), .ZN(n1027) );
NAND3_X1 U741 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1014) );
NAND3_X1 U742 ( .A1(n1022), .A2(n1041), .A3(n1026), .ZN(n1040) );
NAND2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U744 ( .A1(n1035), .A2(n1044), .A3(n1045), .ZN(n1043) );
XOR2_X1 U745 ( .A(KEYINPUT29), .B(n1034), .Z(n1044) );
NAND2_X1 U746 ( .A1(n1024), .A2(n1046), .ZN(n1042) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U748 ( .A1(n1049), .A2(n1050), .A3(n1034), .ZN(n1048) );
NAND3_X1 U749 ( .A1(n1035), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND4_X1 U750 ( .A1(n1023), .A2(n1024), .A3(n1053), .A4(n1054), .ZN(n1038) );
AND3_X1 U751 ( .A1(n1034), .A2(n1035), .A3(n1026), .ZN(n1023) );
NOR3_X1 U752 ( .A1(n1016), .A2(G952), .A3(n1055), .ZN(n1012) );
INV_X1 U753 ( .A(n1039), .ZN(n1055) );
NAND4_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1039) );
NOR4_X1 U755 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
AND3_X1 U756 ( .A1(KEYINPUT45), .A2(n1064), .A3(n1065), .ZN(n1063) );
NOR2_X1 U757 ( .A1(KEYINPUT45), .A2(n1065), .ZN(n1062) );
XOR2_X1 U758 ( .A(KEYINPUT36), .B(n1066), .Z(n1061) );
NAND3_X1 U759 ( .A1(n1067), .A2(n1068), .A3(n1049), .ZN(n1060) );
XOR2_X1 U760 ( .A(KEYINPUT8), .B(n1069), .Z(n1068) );
NOR3_X1 U761 ( .A1(n1070), .A2(n1051), .A3(n1071), .ZN(n1058) );
NAND2_X1 U762 ( .A1(n1072), .A2(n1073), .ZN(G72) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
OR2_X1 U764 ( .A1(n1076), .A2(G227), .ZN(n1075) );
INV_X1 U765 ( .A(n1077), .ZN(n1074) );
NAND3_X1 U766 ( .A1(G953), .A2(n1078), .A3(n1077), .ZN(n1072) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1077) );
NOR2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U769 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U770 ( .A(G125), .B(n1085), .Z(n1084) );
NOR2_X1 U771 ( .A1(KEYINPUT50), .A2(n1086), .ZN(n1085) );
XOR2_X1 U772 ( .A(n1087), .B(G131), .Z(n1086) );
NOR2_X1 U773 ( .A1(G900), .A2(n1076), .ZN(n1081) );
NAND3_X1 U774 ( .A1(n1088), .A2(n1076), .A3(KEYINPUT23), .ZN(n1079) );
NAND2_X1 U775 ( .A1(G900), .A2(G227), .ZN(n1078) );
XOR2_X1 U776 ( .A(n1089), .B(n1090), .Z(G69) );
XOR2_X1 U777 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U779 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U780 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
XOR2_X1 U781 ( .A(n1099), .B(KEYINPUT0), .Z(n1098) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1100), .ZN(n1097) );
XNOR2_X1 U784 ( .A(KEYINPUT30), .B(n1102), .ZN(n1100) );
NOR2_X1 U785 ( .A1(G898), .A2(n1076), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1076), .A2(n1103), .ZN(n1091) );
XOR2_X1 U787 ( .A(KEYINPUT28), .B(n1104), .Z(n1103) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
AND2_X1 U789 ( .A1(n1107), .A2(n1076), .ZN(n1089) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(G66) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
AND2_X1 U795 ( .A1(n1117), .A2(n1116), .ZN(n1110) );
INV_X1 U796 ( .A(KEYINPUT6), .ZN(n1117) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1118), .ZN(G63) );
XOR2_X1 U798 ( .A(n1119), .B(n1120), .Z(n1118) );
AND2_X1 U799 ( .A1(G478), .A2(n1121), .ZN(n1120) );
NAND2_X1 U800 ( .A1(KEYINPUT20), .A2(n1122), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1108), .A2(n1123), .ZN(G60) );
XOR2_X1 U802 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND3_X1 U803 ( .A1(G902), .A2(n1126), .A3(G475), .ZN(n1125) );
XOR2_X1 U804 ( .A(KEYINPUT10), .B(n1127), .Z(n1126) );
XOR2_X1 U805 ( .A(G104), .B(n1128), .Z(G6) );
NOR2_X1 U806 ( .A1(n1108), .A2(n1129), .ZN(G57) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U810 ( .A1(KEYINPUT47), .A2(n1136), .ZN(n1135) );
AND2_X1 U811 ( .A1(G472), .A2(n1121), .ZN(n1134) );
XNOR2_X1 U812 ( .A(n1137), .B(n1138), .ZN(n1130) );
XOR2_X1 U813 ( .A(KEYINPUT48), .B(G101), .Z(n1138) );
NOR2_X1 U814 ( .A1(n1108), .A2(n1139), .ZN(G54) );
XOR2_X1 U815 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U816 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XNOR2_X1 U818 ( .A(KEYINPUT32), .B(n1146), .ZN(n1144) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
XOR2_X1 U820 ( .A(n1146), .B(KEYINPUT13), .Z(n1148) );
NAND2_X1 U821 ( .A1(n1121), .A2(G469), .ZN(n1146) );
INV_X1 U822 ( .A(n1115), .ZN(n1121) );
INV_X1 U823 ( .A(n1145), .ZN(n1147) );
NOR2_X1 U824 ( .A1(n1108), .A2(n1149), .ZN(G51) );
NOR2_X1 U825 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U827 ( .A1(n1154), .A2(n1115), .ZN(n1153) );
NAND2_X1 U828 ( .A1(G902), .A2(n1015), .ZN(n1115) );
INV_X1 U829 ( .A(n1127), .ZN(n1015) );
NOR2_X1 U830 ( .A1(n1107), .A2(n1088), .ZN(n1127) );
NAND4_X1 U831 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1088) );
NOR4_X1 U832 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
INV_X1 U833 ( .A(n1163), .ZN(n1162) );
NAND2_X1 U834 ( .A1(n1037), .A2(n1164), .ZN(n1157) );
NAND2_X1 U835 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND3_X1 U836 ( .A1(n1021), .A2(n1033), .A3(n1167), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1168), .B(KEYINPUT39), .Z(n1167) );
NAND2_X1 U838 ( .A1(n1169), .A2(n1168), .ZN(n1165) );
NAND4_X1 U839 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1107) );
NOR4_X1 U840 ( .A1(n1174), .A2(n1175), .A3(n1011), .A4(n1128), .ZN(n1173) );
AND3_X1 U841 ( .A1(n1176), .A2(n1035), .A3(n1021), .ZN(n1128) );
AND3_X1 U842 ( .A1(n1045), .A2(n1035), .A3(n1176), .ZN(n1011) );
NOR2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(n1172) );
NOR3_X1 U844 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
INV_X1 U846 ( .A(KEYINPUT16), .ZN(n1183) );
AND3_X1 U847 ( .A1(n1184), .A2(n1036), .A3(n1022), .ZN(n1182) );
INV_X1 U848 ( .A(n1185), .ZN(n1184) );
NOR2_X1 U849 ( .A1(KEYINPUT16), .A2(n1186), .ZN(n1180) );
INV_X1 U850 ( .A(n1187), .ZN(n1177) );
NOR2_X1 U851 ( .A1(n1188), .A2(n1189), .ZN(n1152) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(n1189) );
INV_X1 U853 ( .A(KEYINPUT44), .ZN(n1188) );
NOR2_X1 U854 ( .A1(KEYINPUT44), .A2(n1192), .ZN(n1150) );
XOR2_X1 U855 ( .A(n1191), .B(n1193), .Z(n1192) );
INV_X1 U856 ( .A(n1190), .ZN(n1193) );
XOR2_X1 U857 ( .A(n1194), .B(n1195), .Z(n1191) );
NAND3_X1 U858 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1194) );
NAND2_X1 U859 ( .A1(G125), .A2(n1199), .ZN(n1198) );
OR3_X1 U860 ( .A1(n1199), .A2(G125), .A3(KEYINPUT33), .ZN(n1197) );
NAND2_X1 U861 ( .A1(KEYINPUT12), .A2(n1200), .ZN(n1199) );
NAND2_X1 U862 ( .A1(KEYINPUT33), .A2(n1201), .ZN(n1196) );
INV_X1 U863 ( .A(n1200), .ZN(n1201) );
NOR2_X1 U864 ( .A1(n1076), .A2(G952), .ZN(n1108) );
XOR2_X1 U865 ( .A(n1160), .B(n1202), .Z(G48) );
NOR2_X1 U866 ( .A1(KEYINPUT9), .A2(n1203), .ZN(n1202) );
AND3_X1 U867 ( .A1(n1021), .A2(n1204), .A3(n1205), .ZN(n1160) );
XNOR2_X1 U868 ( .A(G143), .B(n1155), .ZN(G45) );
NAND4_X1 U869 ( .A1(n1036), .A2(n1204), .A3(n1033), .A4(n1206), .ZN(n1155) );
AND3_X1 U870 ( .A1(n1066), .A2(n1168), .A3(n1207), .ZN(n1206) );
XNOR2_X1 U871 ( .A(G140), .B(n1156), .ZN(G42) );
NAND2_X1 U872 ( .A1(n1208), .A2(n1037), .ZN(n1156) );
XOR2_X1 U873 ( .A(n1209), .B(n1210), .Z(G39) );
NAND3_X1 U874 ( .A1(n1037), .A2(n1169), .A3(n1211), .ZN(n1210) );
XOR2_X1 U875 ( .A(n1168), .B(KEYINPUT61), .Z(n1211) );
INV_X1 U876 ( .A(n1179), .ZN(n1169) );
XNOR2_X1 U877 ( .A(G134), .B(n1212), .ZN(G36) );
NAND2_X1 U878 ( .A1(KEYINPUT38), .A2(n1159), .ZN(n1212) );
AND4_X1 U879 ( .A1(n1037), .A2(n1033), .A3(n1045), .A4(n1168), .ZN(n1159) );
XOR2_X1 U880 ( .A(n1213), .B(n1214), .Z(G33) );
XNOR2_X1 U881 ( .A(G131), .B(KEYINPUT21), .ZN(n1214) );
NAND4_X1 U882 ( .A1(n1215), .A2(n1037), .A3(n1021), .A4(n1033), .ZN(n1213) );
AND2_X1 U883 ( .A1(n1034), .A2(n1204), .ZN(n1037) );
NOR2_X1 U884 ( .A1(n1069), .A2(n1216), .ZN(n1034) );
XOR2_X1 U885 ( .A(n1168), .B(KEYINPUT37), .Z(n1215) );
XOR2_X1 U886 ( .A(G128), .B(n1217), .Z(G30) );
NOR2_X1 U887 ( .A1(KEYINPUT15), .A2(n1163), .ZN(n1217) );
NAND3_X1 U888 ( .A1(n1045), .A2(n1218), .A3(n1205), .ZN(n1163) );
AND4_X1 U889 ( .A1(n1036), .A2(n1219), .A3(n1168), .A4(n1050), .ZN(n1205) );
XOR2_X1 U890 ( .A(G101), .B(n1175), .Z(G3) );
AND3_X1 U891 ( .A1(n1033), .A2(n1176), .A3(n1024), .ZN(n1175) );
XOR2_X1 U892 ( .A(G125), .B(n1161), .Z(G27) );
AND3_X1 U893 ( .A1(n1022), .A2(n1036), .A3(n1208), .ZN(n1161) );
AND4_X1 U894 ( .A1(n1049), .A2(n1021), .A3(n1168), .A4(n1050), .ZN(n1208) );
NAND2_X1 U895 ( .A1(n1220), .A2(n1221), .ZN(n1168) );
NAND4_X1 U896 ( .A1(n1222), .A2(G953), .A3(G902), .A4(n1223), .ZN(n1221) );
INV_X1 U897 ( .A(G900), .ZN(n1223) );
XOR2_X1 U898 ( .A(n1224), .B(KEYINPUT55), .Z(n1222) );
XOR2_X1 U899 ( .A(KEYINPUT2), .B(n1026), .Z(n1220) );
INV_X1 U900 ( .A(n1225), .ZN(n1026) );
XOR2_X1 U901 ( .A(n1226), .B(n1187), .Z(G24) );
NAND4_X1 U902 ( .A1(n1186), .A2(n1035), .A3(n1066), .A4(n1207), .ZN(n1187) );
NOR2_X1 U903 ( .A1(n1050), .A2(n1219), .ZN(n1035) );
XOR2_X1 U904 ( .A(G119), .B(n1227), .Z(G21) );
NOR2_X1 U905 ( .A1(n1228), .A2(n1179), .ZN(n1227) );
NAND3_X1 U906 ( .A1(n1219), .A2(n1050), .A3(n1024), .ZN(n1179) );
XOR2_X1 U907 ( .A(G116), .B(n1174), .Z(G18) );
AND3_X1 U908 ( .A1(n1186), .A2(n1045), .A3(n1033), .ZN(n1174) );
AND2_X1 U909 ( .A1(n1229), .A2(n1207), .ZN(n1045) );
XNOR2_X1 U910 ( .A(G113), .B(n1170), .ZN(G15) );
NAND3_X1 U911 ( .A1(n1033), .A2(n1186), .A3(n1021), .ZN(n1170) );
NOR2_X1 U912 ( .A1(n1207), .A2(n1229), .ZN(n1021) );
INV_X1 U913 ( .A(n1228), .ZN(n1186) );
NAND3_X1 U914 ( .A1(n1036), .A2(n1185), .A3(n1022), .ZN(n1228) );
NOR2_X1 U915 ( .A1(n1230), .A2(n1231), .ZN(n1022) );
INV_X1 U916 ( .A(n1053), .ZN(n1230) );
AND2_X1 U917 ( .A1(n1232), .A2(n1219), .ZN(n1033) );
INV_X1 U918 ( .A(n1049), .ZN(n1219) );
XOR2_X1 U919 ( .A(n1050), .B(KEYINPUT3), .Z(n1232) );
XOR2_X1 U920 ( .A(n1233), .B(n1171), .Z(G12) );
NAND4_X1 U921 ( .A1(n1024), .A2(n1176), .A3(n1049), .A4(n1050), .ZN(n1171) );
OR2_X1 U922 ( .A1(n1070), .A2(n1234), .ZN(n1050) );
AND2_X1 U923 ( .A1(n1065), .A2(n1064), .ZN(n1234) );
NOR2_X1 U924 ( .A1(n1064), .A2(n1065), .ZN(n1070) );
INV_X1 U925 ( .A(n1114), .ZN(n1065) );
NAND2_X1 U926 ( .A1(G217), .A2(n1235), .ZN(n1114) );
OR2_X1 U927 ( .A1(n1116), .A2(G902), .ZN(n1064) );
XNOR2_X1 U928 ( .A(n1236), .B(n1237), .ZN(n1116) );
XOR2_X1 U929 ( .A(n1233), .B(n1238), .Z(n1237) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U931 ( .A1(G119), .A2(n1241), .ZN(n1240) );
XOR2_X1 U932 ( .A(n1242), .B(KEYINPUT27), .Z(n1239) );
OR2_X1 U933 ( .A1(n1241), .A2(G119), .ZN(n1242) );
XOR2_X1 U934 ( .A(n1243), .B(n1244), .Z(n1236) );
NOR2_X1 U935 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U936 ( .A(KEYINPUT14), .B(n1247), .Z(n1246) );
NOR2_X1 U937 ( .A1(n1209), .A2(n1248), .ZN(n1247) );
AND2_X1 U938 ( .A1(n1209), .A2(n1248), .ZN(n1245) );
NAND3_X1 U939 ( .A1(G234), .A2(n1076), .A3(G221), .ZN(n1248) );
NAND2_X1 U940 ( .A1(KEYINPUT42), .A2(n1249), .ZN(n1243) );
XOR2_X1 U941 ( .A(n1250), .B(G472), .Z(n1049) );
NAND2_X1 U942 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U943 ( .A(n1253), .B(n1254), .Z(n1251) );
XNOR2_X1 U944 ( .A(n1255), .B(n1136), .ZN(n1254) );
XOR2_X1 U945 ( .A(n1256), .B(n1200), .Z(n1136) );
NAND2_X1 U946 ( .A1(KEYINPUT53), .A2(n1137), .ZN(n1255) );
AND3_X1 U947 ( .A1(n1257), .A2(n1076), .A3(G210), .ZN(n1137) );
XOR2_X1 U948 ( .A(G101), .B(n1258), .Z(n1253) );
NOR2_X1 U949 ( .A1(KEYINPUT41), .A2(n1132), .ZN(n1258) );
XNOR2_X1 U950 ( .A(n1102), .B(KEYINPUT57), .ZN(n1132) );
AND3_X1 U951 ( .A1(n1218), .A2(n1185), .A3(n1036), .ZN(n1176) );
NOR2_X1 U952 ( .A1(n1052), .A2(n1216), .ZN(n1036) );
XNOR2_X1 U953 ( .A(n1051), .B(KEYINPUT58), .ZN(n1216) );
AND2_X1 U954 ( .A1(n1259), .A2(n1260), .ZN(n1051) );
XOR2_X1 U955 ( .A(KEYINPUT62), .B(G214), .Z(n1259) );
INV_X1 U956 ( .A(n1069), .ZN(n1052) );
XNOR2_X1 U957 ( .A(n1154), .B(n1261), .ZN(n1069) );
NOR2_X1 U958 ( .A1(G902), .A2(n1262), .ZN(n1261) );
XOR2_X1 U959 ( .A(n1190), .B(n1263), .Z(n1262) );
NOR2_X1 U960 ( .A1(KEYINPUT54), .A2(n1264), .ZN(n1263) );
XOR2_X1 U961 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U962 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U963 ( .A1(KEYINPUT7), .A2(n1200), .ZN(n1268) );
NAND2_X1 U964 ( .A1(n1269), .A2(n1270), .ZN(n1200) );
NAND2_X1 U965 ( .A1(n1271), .A2(n1203), .ZN(n1270) );
XOR2_X1 U966 ( .A(KEYINPUT35), .B(n1272), .Z(n1271) );
NAND2_X1 U967 ( .A1(n1273), .A2(G146), .ZN(n1269) );
XNOR2_X1 U968 ( .A(G143), .B(n1274), .ZN(n1273) );
INV_X1 U969 ( .A(G125), .ZN(n1267) );
NAND2_X1 U970 ( .A1(KEYINPUT49), .A2(n1195), .ZN(n1265) );
NOR2_X1 U971 ( .A1(n1105), .A2(G953), .ZN(n1195) );
INV_X1 U972 ( .A(G224), .ZN(n1105) );
XOR2_X1 U973 ( .A(n1275), .B(n1096), .Z(n1190) );
XOR2_X1 U974 ( .A(G110), .B(G122), .Z(n1096) );
NAND2_X1 U975 ( .A1(KEYINPUT17), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U976 ( .A(n1102), .B(n1101), .ZN(n1276) );
XNOR2_X1 U977 ( .A(G101), .B(n1277), .ZN(n1101) );
XNOR2_X1 U978 ( .A(n1278), .B(n1279), .ZN(n1102) );
XOR2_X1 U979 ( .A(KEYINPUT26), .B(G119), .Z(n1279) );
XNOR2_X1 U980 ( .A(G113), .B(G116), .ZN(n1278) );
NAND2_X1 U981 ( .A1(G210), .A2(n1260), .ZN(n1154) );
NAND2_X1 U982 ( .A1(n1252), .A2(n1257), .ZN(n1260) );
NAND2_X1 U983 ( .A1(n1225), .A2(n1280), .ZN(n1185) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1106), .ZN(n1280) );
INV_X1 U985 ( .A(G898), .ZN(n1106) );
NAND3_X1 U986 ( .A1(n1281), .A2(n1224), .A3(G952), .ZN(n1225) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1224) );
INV_X1 U988 ( .A(n1016), .ZN(n1281) );
XOR2_X1 U989 ( .A(n1076), .B(KEYINPUT43), .Z(n1016) );
XOR2_X1 U990 ( .A(n1204), .B(KEYINPUT60), .Z(n1218) );
NOR2_X1 U991 ( .A1(n1231), .A2(n1053), .ZN(n1204) );
NOR2_X1 U992 ( .A1(n1282), .A2(n1071), .ZN(n1053) );
NOR3_X1 U993 ( .A1(G469), .A2(G902), .A3(n1283), .ZN(n1071) );
XOR2_X1 U994 ( .A(KEYINPUT34), .B(n1057), .Z(n1282) );
NAND2_X1 U995 ( .A1(G469), .A2(n1284), .ZN(n1057) );
OR2_X1 U996 ( .A1(n1283), .A2(G902), .ZN(n1284) );
XNOR2_X1 U997 ( .A(n1285), .B(n1141), .ZN(n1283) );
XNOR2_X1 U998 ( .A(n1286), .B(n1287), .ZN(n1141) );
XOR2_X1 U999 ( .A(n1288), .B(n1083), .Z(n1287) );
XOR2_X1 U1000 ( .A(n1289), .B(n1290), .Z(n1083) );
XOR2_X1 U1001 ( .A(n1291), .B(n1292), .Z(n1289) );
NOR2_X1 U1002 ( .A1(G143), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1003 ( .A(KEYINPUT52), .B(KEYINPUT22), .ZN(n1293) );
NAND2_X1 U1004 ( .A1(KEYINPUT46), .A2(n1274), .ZN(n1291) );
XNOR2_X1 U1005 ( .A(KEYINPUT35), .B(n1241), .ZN(n1274) );
INV_X1 U1006 ( .A(G128), .ZN(n1241) );
NAND2_X1 U1007 ( .A1(G227), .A2(n1076), .ZN(n1288) );
XOR2_X1 U1008 ( .A(n1256), .B(G110), .Z(n1286) );
NAND2_X1 U1009 ( .A1(n1294), .A2(n1295), .ZN(n1256) );
NAND2_X1 U1010 ( .A1(G131), .A2(n1087), .ZN(n1295) );
XOR2_X1 U1011 ( .A(n1296), .B(KEYINPUT5), .Z(n1294) );
OR2_X1 U1012 ( .A1(n1087), .A2(G131), .ZN(n1296) );
XOR2_X1 U1013 ( .A(n1209), .B(n1297), .Z(n1087) );
INV_X1 U1014 ( .A(G137), .ZN(n1209) );
XOR2_X1 U1015 ( .A(n1145), .B(KEYINPUT51), .Z(n1285) );
XOR2_X1 U1016 ( .A(n1298), .B(G101), .Z(n1145) );
NAND2_X1 U1017 ( .A1(KEYINPUT18), .A2(n1277), .ZN(n1298) );
XOR2_X1 U1018 ( .A(G104), .B(G107), .Z(n1277) );
XNOR2_X1 U1019 ( .A(n1054), .B(KEYINPUT56), .ZN(n1231) );
INV_X1 U1020 ( .A(n1056), .ZN(n1054) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1235), .ZN(n1056) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1252), .ZN(n1235) );
NOR2_X1 U1023 ( .A1(n1207), .A2(n1066), .ZN(n1024) );
INV_X1 U1024 ( .A(n1229), .ZN(n1066) );
XNOR2_X1 U1025 ( .A(G475), .B(n1299), .ZN(n1229) );
AND2_X1 U1026 ( .A1(n1124), .A2(n1252), .ZN(n1299) );
NAND2_X1 U1027 ( .A1(n1300), .A2(n1301), .ZN(n1124) );
NAND2_X1 U1028 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1029 ( .A(KEYINPUT31), .B(n1304), .Z(n1300) );
NOR2_X1 U1030 ( .A1(n1303), .A2(n1302), .ZN(n1304) );
XOR2_X1 U1031 ( .A(n1305), .B(n1306), .Z(n1302) );
XNOR2_X1 U1032 ( .A(n1307), .B(n1308), .ZN(n1306) );
XOR2_X1 U1033 ( .A(KEYINPUT4), .B(G143), .Z(n1308) );
NAND3_X1 U1034 ( .A1(n1257), .A2(n1076), .A3(G214), .ZN(n1307) );
INV_X1 U1035 ( .A(G237), .ZN(n1257) );
XNOR2_X1 U1036 ( .A(n1309), .B(n1249), .ZN(n1305) );
XOR2_X1 U1037 ( .A(G125), .B(n1290), .Z(n1249) );
XNOR2_X1 U1038 ( .A(G140), .B(n1203), .ZN(n1290) );
INV_X1 U1039 ( .A(G146), .ZN(n1203) );
NAND2_X1 U1040 ( .A1(KEYINPUT11), .A2(G131), .ZN(n1309) );
XOR2_X1 U1041 ( .A(G104), .B(n1310), .Z(n1303) );
XOR2_X1 U1042 ( .A(G122), .B(G113), .Z(n1310) );
XOR2_X1 U1043 ( .A(n1311), .B(n1067), .Z(n1207) );
XOR2_X1 U1044 ( .A(n1312), .B(G478), .Z(n1067) );
NAND2_X1 U1045 ( .A1(n1122), .A2(n1252), .ZN(n1312) );
INV_X1 U1046 ( .A(G902), .ZN(n1252) );
XNOR2_X1 U1047 ( .A(n1313), .B(n1314), .ZN(n1122) );
XOR2_X1 U1048 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1049 ( .A(G107), .B(G116), .ZN(n1316) );
NAND3_X1 U1050 ( .A1(G234), .A2(n1076), .A3(G217), .ZN(n1315) );
INV_X1 U1051 ( .A(G953), .ZN(n1076) );
XOR2_X1 U1052 ( .A(n1317), .B(n1297), .Z(n1313) );
XOR2_X1 U1053 ( .A(G134), .B(KEYINPUT24), .Z(n1297) );
XNOR2_X1 U1054 ( .A(n1318), .B(n1319), .ZN(n1317) );
NAND2_X1 U1055 ( .A1(KEYINPUT25), .A2(n1226), .ZN(n1319) );
INV_X1 U1056 ( .A(G122), .ZN(n1226) );
NAND2_X1 U1057 ( .A1(KEYINPUT1), .A2(n1272), .ZN(n1318) );
XOR2_X1 U1058 ( .A(G128), .B(G143), .Z(n1272) );
XNOR2_X1 U1059 ( .A(KEYINPUT40), .B(KEYINPUT19), .ZN(n1311) );
INV_X1 U1060 ( .A(G110), .ZN(n1233) );
endmodule


