//Key = 0110101011010110000100100001111100011000010011001100011111000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271;

XNOR2_X1 U705 ( .A(G107), .B(n973), .ZN(G9) );
NOR2_X1 U706 ( .A1(n974), .A2(n975), .ZN(G75) );
NOR4_X1 U707 ( .A1(G953), .A2(n976), .A3(n977), .A4(n978), .ZN(n975) );
NOR2_X1 U708 ( .A1(n979), .A2(n980), .ZN(n977) );
NOR2_X1 U709 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR3_X1 U710 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
NOR2_X1 U711 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U712 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR2_X1 U713 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR2_X1 U714 ( .A1(n992), .A2(n993), .ZN(n986) );
NOR3_X1 U715 ( .A1(n993), .A2(n994), .A3(n989), .ZN(n981) );
INV_X1 U716 ( .A(n995), .ZN(n989) );
NOR3_X1 U717 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n994) );
NOR2_X1 U718 ( .A1(n999), .A2(n983), .ZN(n998) );
NOR2_X1 U719 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR2_X1 U721 ( .A1(n1004), .A2(n1005), .ZN(n997) );
XOR2_X1 U722 ( .A(n985), .B(KEYINPUT40), .Z(n1005) );
XOR2_X1 U723 ( .A(n1006), .B(KEYINPUT39), .Z(n1004) );
NAND2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U725 ( .A1(n1009), .A2(n985), .ZN(n996) );
INV_X1 U726 ( .A(n1010), .ZN(n985) );
INV_X1 U727 ( .A(n1011), .ZN(n993) );
NOR3_X1 U728 ( .A1(n976), .A2(G953), .A3(G952), .ZN(n974) );
AND4_X1 U729 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n976) );
NOR4_X1 U730 ( .A1(n1008), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1015) );
XNOR2_X1 U731 ( .A(n1019), .B(n1020), .ZN(n1017) );
NOR2_X1 U732 ( .A1(G478), .A2(KEYINPUT24), .ZN(n1020) );
NOR2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1014) );
XOR2_X1 U734 ( .A(n1023), .B(n1024), .Z(n1022) );
XNOR2_X1 U735 ( .A(n1025), .B(n1026), .ZN(n1021) );
NAND2_X1 U736 ( .A1(KEYINPUT56), .A2(n1027), .ZN(n1026) );
XOR2_X1 U737 ( .A(n1028), .B(n1029), .Z(n1013) );
XOR2_X1 U738 ( .A(n1030), .B(n1031), .Z(n1012) );
XOR2_X1 U739 ( .A(n1032), .B(n1033), .Z(G72) );
NOR2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U741 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1032) );
NAND2_X1 U743 ( .A1(n1040), .A2(n1035), .ZN(n1039) );
XNOR2_X1 U744 ( .A(n1041), .B(n1042), .ZN(n1040) );
NOR3_X1 U745 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
XOR2_X1 U746 ( .A(n1046), .B(KEYINPUT32), .Z(n1045) );
OR2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U748 ( .A1(G900), .A2(n1041), .A3(G953), .ZN(n1038) );
XNOR2_X1 U749 ( .A(n1049), .B(n1050), .ZN(n1041) );
XOR2_X1 U750 ( .A(n1051), .B(n1052), .Z(G69) );
XOR2_X1 U751 ( .A(n1053), .B(n1054), .Z(n1052) );
NAND2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U753 ( .A1(G953), .A2(n1057), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1058), .B(n1059), .ZN(n1055) );
NAND2_X1 U755 ( .A1(n1035), .A2(n1060), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1035), .ZN(n1051) );
AND2_X1 U758 ( .A1(G224), .A2(G898), .ZN(n1063) );
NOR2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(G66) );
NOR3_X1 U760 ( .A1(n1025), .A2(n1066), .A3(n1067), .ZN(n1065) );
AND3_X1 U761 ( .A1(n1068), .A2(n1027), .A3(n1069), .ZN(n1067) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1068), .ZN(n1066) );
AND2_X1 U763 ( .A1(n978), .A2(n1027), .ZN(n1070) );
INV_X1 U764 ( .A(n1071), .ZN(n1027) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1072), .ZN(G63) );
NOR3_X1 U766 ( .A1(n1019), .A2(n1073), .A3(n1074), .ZN(n1072) );
AND3_X1 U767 ( .A1(n1075), .A2(n1069), .A3(G478), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1075), .ZN(n1073) );
AND2_X1 U769 ( .A1(n978), .A2(G478), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1064), .A2(n1077), .ZN(G60) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1077) );
XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n1080), .ZN(n1079) );
NOR3_X1 U773 ( .A1(n1081), .A2(KEYINPUT37), .A3(n1028), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(G6) );
OR2_X1 U775 ( .A1(n1084), .A2(G104), .ZN(n1083) );
XOR2_X1 U776 ( .A(n1085), .B(KEYINPUT61), .Z(n1082) );
NAND2_X1 U777 ( .A1(G104), .A2(n1084), .ZN(n1085) );
NOR2_X1 U778 ( .A1(n1064), .A2(n1086), .ZN(G57) );
XOR2_X1 U779 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U780 ( .A(n1089), .B(n1090), .ZN(n1088) );
XNOR2_X1 U781 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U782 ( .A1(KEYINPUT5), .A2(n1093), .ZN(n1092) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(n1087) );
XOR2_X1 U784 ( .A(KEYINPUT26), .B(G101), .Z(n1095) );
XOR2_X1 U785 ( .A(n1096), .B(n1097), .Z(n1094) );
NOR2_X1 U786 ( .A1(n1031), .A2(n1081), .ZN(n1097) );
INV_X1 U787 ( .A(G472), .ZN(n1031) );
NOR2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(G54) );
XOR2_X1 U789 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U791 ( .A1(n1023), .A2(n1081), .ZN(n1102) );
XOR2_X1 U792 ( .A(n1104), .B(KEYINPUT8), .Z(n1098) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
INV_X1 U794 ( .A(G952), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1035), .B(KEYINPUT9), .Z(n1105) );
NOR2_X1 U796 ( .A1(n1064), .A2(n1107), .ZN(G51) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1107) );
XNOR2_X1 U798 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U799 ( .A1(KEYINPUT43), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U800 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND3_X1 U801 ( .A1(n1069), .A2(n1115), .A3(KEYINPUT11), .ZN(n1110) );
INV_X1 U802 ( .A(n1081), .ZN(n1069) );
NAND2_X1 U803 ( .A1(G902), .A2(n978), .ZN(n1081) );
NAND4_X1 U804 ( .A1(n1061), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n978) );
NOR3_X1 U805 ( .A1(n1119), .A2(n1047), .A3(n1120), .ZN(n1118) );
XNOR2_X1 U806 ( .A(KEYINPUT0), .B(n1062), .ZN(n1120) );
NAND3_X1 U807 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1047) );
NAND3_X1 U808 ( .A1(n1124), .A2(n990), .A3(n1125), .ZN(n1123) );
XOR2_X1 U809 ( .A(KEYINPUT20), .B(n1044), .Z(n1119) );
INV_X1 U810 ( .A(n1126), .ZN(n1044) );
INV_X1 U811 ( .A(n1043), .ZN(n1117) );
NAND3_X1 U812 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1043) );
XOR2_X1 U813 ( .A(KEYINPUT45), .B(n1048), .Z(n1116) );
AND3_X1 U814 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1061) );
AND3_X1 U815 ( .A1(n1084), .A2(n973), .A3(n1133), .ZN(n1132) );
NAND3_X1 U816 ( .A1(n1001), .A2(n990), .A3(n1134), .ZN(n973) );
NAND3_X1 U817 ( .A1(n1134), .A2(n1001), .A3(n991), .ZN(n1084) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
NAND2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND3_X1 U820 ( .A1(n1001), .A2(n1139), .A3(n1140), .ZN(n1138) );
INV_X1 U821 ( .A(n992), .ZN(n1139) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n992) );
NAND2_X1 U823 ( .A1(n1143), .A2(n990), .ZN(n1130) );
NOR2_X1 U824 ( .A1(n1035), .A2(G952), .ZN(n1064) );
XNOR2_X1 U825 ( .A(G146), .B(n1129), .ZN(G48) );
NAND3_X1 U826 ( .A1(n1124), .A2(n991), .A3(n1125), .ZN(n1129) );
XOR2_X1 U827 ( .A(n1126), .B(n1144), .Z(G45) );
NAND2_X1 U828 ( .A1(KEYINPUT53), .A2(n1145), .ZN(n1144) );
XOR2_X1 U829 ( .A(KEYINPUT51), .B(G143), .Z(n1145) );
NAND4_X1 U830 ( .A1(n1124), .A2(n1142), .A3(n1146), .A4(n1147), .ZN(n1126) );
XOR2_X1 U831 ( .A(n1148), .B(n1127), .Z(G42) );
NAND3_X1 U832 ( .A1(n1141), .A2(n991), .A3(n1149), .ZN(n1127) );
XOR2_X1 U833 ( .A(n1128), .B(n1150), .Z(G39) );
NAND2_X1 U834 ( .A1(KEYINPUT31), .A2(G137), .ZN(n1150) );
NAND3_X1 U835 ( .A1(n1125), .A2(n1149), .A3(n1011), .ZN(n1128) );
XOR2_X1 U836 ( .A(G134), .B(n1048), .Z(G36) );
AND3_X1 U837 ( .A1(n1142), .A2(n990), .A3(n1149), .ZN(n1048) );
XNOR2_X1 U838 ( .A(n1121), .B(n1151), .ZN(G33) );
XOR2_X1 U839 ( .A(KEYINPUT58), .B(G131), .Z(n1151) );
NAND3_X1 U840 ( .A1(n1142), .A2(n991), .A3(n1149), .ZN(n1121) );
NOR3_X1 U841 ( .A1(n1152), .A2(n1153), .A3(n983), .ZN(n1149) );
NAND2_X1 U842 ( .A1(n1007), .A2(n1154), .ZN(n983) );
XOR2_X1 U843 ( .A(n1155), .B(n1156), .Z(G30) );
NAND4_X1 U844 ( .A1(KEYINPUT27), .A2(n1125), .A3(n1124), .A4(n990), .ZN(n1156) );
INV_X1 U845 ( .A(n1157), .ZN(n990) );
NOR3_X1 U846 ( .A1(n1009), .A2(n1153), .A3(n1152), .ZN(n1124) );
XNOR2_X1 U847 ( .A(G101), .B(n1158), .ZN(G3) );
NAND2_X1 U848 ( .A1(n1159), .A2(n1135), .ZN(n1158) );
XOR2_X1 U849 ( .A(n1160), .B(KEYINPUT13), .Z(n1159) );
NAND3_X1 U850 ( .A1(n1142), .A2(n1161), .A3(n1140), .ZN(n1160) );
XOR2_X1 U851 ( .A(KEYINPUT10), .B(n1001), .Z(n1161) );
XNOR2_X1 U852 ( .A(G125), .B(n1122), .ZN(G27) );
NAND4_X1 U853 ( .A1(n1141), .A2(n991), .A3(n1162), .A4(n1010), .ZN(n1122) );
NOR2_X1 U854 ( .A1(n1153), .A2(n1009), .ZN(n1162) );
AND2_X1 U855 ( .A1(n980), .A2(n1163), .ZN(n1153) );
NAND4_X1 U856 ( .A1(G953), .A2(G902), .A3(n1164), .A4(n1037), .ZN(n1163) );
INV_X1 U857 ( .A(G900), .ZN(n1037) );
NAND2_X1 U858 ( .A1(n1165), .A2(n1166), .ZN(G24) );
NAND2_X1 U859 ( .A1(G122), .A2(n1133), .ZN(n1166) );
XOR2_X1 U860 ( .A(n1167), .B(KEYINPUT60), .Z(n1165) );
OR2_X1 U861 ( .A1(n1133), .A2(G122), .ZN(n1167) );
NAND4_X1 U862 ( .A1(n1147), .A2(n1010), .A3(n1146), .A4(n1134), .ZN(n1133) );
AND3_X1 U863 ( .A1(n1135), .A2(n1168), .A3(n995), .ZN(n1134) );
NOR2_X1 U864 ( .A1(n1169), .A2(n1170), .ZN(n995) );
XOR2_X1 U865 ( .A(G119), .B(n1171), .Z(G21) );
NOR2_X1 U866 ( .A1(n1172), .A2(n1009), .ZN(n1171) );
XOR2_X1 U867 ( .A(n1137), .B(KEYINPUT15), .Z(n1172) );
NAND3_X1 U868 ( .A1(n1125), .A2(n1010), .A3(n1140), .ZN(n1137) );
AND2_X1 U869 ( .A1(n1170), .A2(n1169), .ZN(n1125) );
XOR2_X1 U870 ( .A(G116), .B(n1173), .Z(G18) );
NOR3_X1 U871 ( .A1(n1174), .A2(KEYINPUT23), .A3(n1157), .ZN(n1173) );
NAND2_X1 U872 ( .A1(n1146), .A2(n1175), .ZN(n1157) );
XOR2_X1 U873 ( .A(n1176), .B(n1062), .Z(G15) );
NAND2_X1 U874 ( .A1(n1143), .A2(n991), .ZN(n1062) );
NOR2_X1 U875 ( .A1(n1175), .A2(n1146), .ZN(n991) );
INV_X1 U876 ( .A(n1147), .ZN(n1175) );
INV_X1 U877 ( .A(n1174), .ZN(n1143) );
NAND4_X1 U878 ( .A1(n1142), .A2(n1010), .A3(n1135), .A4(n1168), .ZN(n1174) );
INV_X1 U879 ( .A(n1009), .ZN(n1135) );
NOR2_X1 U880 ( .A1(n1003), .A2(n1016), .ZN(n1010) );
INV_X1 U881 ( .A(n1002), .ZN(n1016) );
AND2_X1 U882 ( .A1(n1177), .A2(n1170), .ZN(n1142) );
XNOR2_X1 U883 ( .A(G110), .B(n1178), .ZN(G12) );
NAND4_X1 U884 ( .A1(n1179), .A2(n1140), .A3(n1141), .A4(n1001), .ZN(n1178) );
INV_X1 U885 ( .A(n1152), .ZN(n1001) );
NAND2_X1 U886 ( .A1(n1180), .A2(n1003), .ZN(n1152) );
XNOR2_X1 U887 ( .A(n1024), .B(n1181), .ZN(n1003) );
NOR2_X1 U888 ( .A1(KEYINPUT33), .A2(n1023), .ZN(n1181) );
INV_X1 U889 ( .A(G469), .ZN(n1023) );
NAND2_X1 U890 ( .A1(n1182), .A2(n1183), .ZN(n1024) );
XOR2_X1 U891 ( .A(n1184), .B(n1185), .Z(n1182) );
NOR2_X1 U892 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR3_X1 U893 ( .A1(KEYINPUT35), .A2(G110), .A3(n1148), .ZN(n1187) );
INV_X1 U894 ( .A(G140), .ZN(n1148) );
NOR2_X1 U895 ( .A1(n1103), .A2(n1188), .ZN(n1186) );
INV_X1 U896 ( .A(KEYINPUT35), .ZN(n1188) );
XOR2_X1 U897 ( .A(G110), .B(G140), .Z(n1103) );
XNOR2_X1 U898 ( .A(n1100), .B(KEYINPUT46), .ZN(n1184) );
XNOR2_X1 U899 ( .A(n1189), .B(n1190), .ZN(n1100) );
XOR2_X1 U900 ( .A(n1049), .B(n1191), .Z(n1189) );
NOR2_X1 U901 ( .A1(G953), .A2(n1036), .ZN(n1191) );
INV_X1 U902 ( .A(G227), .ZN(n1036) );
XOR2_X1 U903 ( .A(n1192), .B(n1193), .Z(n1049) );
XOR2_X1 U904 ( .A(n1155), .B(n1194), .Z(n1192) );
INV_X1 U905 ( .A(n1093), .ZN(n1194) );
INV_X1 U906 ( .A(G128), .ZN(n1155) );
XOR2_X1 U907 ( .A(n1002), .B(KEYINPUT16), .Z(n1180) );
NAND2_X1 U908 ( .A1(G221), .A2(n1195), .ZN(n1002) );
NOR2_X1 U909 ( .A1(n1170), .A2(n1177), .ZN(n1141) );
INV_X1 U910 ( .A(n1169), .ZN(n1177) );
NAND2_X1 U911 ( .A1(n1196), .A2(n1197), .ZN(n1169) );
OR2_X1 U912 ( .A1(n1071), .A2(n1025), .ZN(n1197) );
XOR2_X1 U913 ( .A(n1198), .B(KEYINPUT62), .Z(n1196) );
NAND2_X1 U914 ( .A1(n1025), .A2(n1071), .ZN(n1198) );
NAND2_X1 U915 ( .A1(G217), .A2(n1195), .ZN(n1071) );
NAND2_X1 U916 ( .A1(G234), .A2(n1183), .ZN(n1195) );
NOR2_X1 U917 ( .A1(n1068), .A2(G902), .ZN(n1025) );
XNOR2_X1 U918 ( .A(n1199), .B(n1200), .ZN(n1068) );
XOR2_X1 U919 ( .A(G119), .B(n1201), .Z(n1200) );
XOR2_X1 U920 ( .A(G137), .B(G128), .Z(n1201) );
XOR2_X1 U921 ( .A(n1202), .B(n1203), .Z(n1199) );
NOR2_X1 U922 ( .A1(KEYINPUT34), .A2(n1204), .ZN(n1203) );
XOR2_X1 U923 ( .A(n1205), .B(n1206), .Z(n1202) );
NOR2_X1 U924 ( .A1(G110), .A2(KEYINPUT12), .ZN(n1206) );
NAND3_X1 U925 ( .A1(n1207), .A2(n1035), .A3(G221), .ZN(n1205) );
XNOR2_X1 U926 ( .A(n1208), .B(G472), .ZN(n1170) );
NAND2_X1 U927 ( .A1(KEYINPUT14), .A2(n1030), .ZN(n1208) );
AND2_X1 U928 ( .A1(n1209), .A2(n1183), .ZN(n1030) );
XOR2_X1 U929 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U930 ( .A(n1093), .B(n1089), .Z(n1211) );
XNOR2_X1 U931 ( .A(n1212), .B(n1213), .ZN(n1089) );
XOR2_X1 U932 ( .A(KEYINPUT38), .B(G119), .Z(n1213) );
XOR2_X1 U933 ( .A(n1176), .B(G116), .Z(n1212) );
XOR2_X1 U934 ( .A(n1214), .B(n1215), .Z(n1093) );
XOR2_X1 U935 ( .A(KEYINPUT29), .B(G137), .Z(n1215) );
XNOR2_X1 U936 ( .A(G131), .B(G134), .ZN(n1214) );
XOR2_X1 U937 ( .A(n1216), .B(n1217), .Z(n1210) );
NOR2_X1 U938 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U939 ( .A(n1220), .B(KEYINPUT4), .Z(n1219) );
NAND2_X1 U940 ( .A1(n1221), .A2(n1096), .ZN(n1220) );
NOR2_X1 U941 ( .A1(n1096), .A2(n1221), .ZN(n1218) );
XOR2_X1 U942 ( .A(KEYINPUT19), .B(G101), .Z(n1221) );
NAND2_X1 U943 ( .A1(n1222), .A2(n1223), .ZN(n1096) );
XNOR2_X1 U944 ( .A(G210), .B(KEYINPUT41), .ZN(n1222) );
NAND2_X1 U945 ( .A1(KEYINPUT54), .A2(n1091), .ZN(n1216) );
AND2_X1 U946 ( .A1(n1011), .A2(n1168), .ZN(n1140) );
NAND2_X1 U947 ( .A1(n980), .A2(n1224), .ZN(n1168) );
NAND4_X1 U948 ( .A1(G953), .A2(G902), .A3(n1164), .A4(n1057), .ZN(n1224) );
INV_X1 U949 ( .A(G898), .ZN(n1057) );
NAND3_X1 U950 ( .A1(n1164), .A2(n1035), .A3(G952), .ZN(n980) );
NAND2_X1 U951 ( .A1(G237), .A2(G234), .ZN(n1164) );
NOR2_X1 U952 ( .A1(n1146), .A2(n1147), .ZN(n1011) );
XOR2_X1 U953 ( .A(n1225), .B(n1029), .Z(n1147) );
NOR2_X1 U954 ( .A1(n1078), .A2(G902), .ZN(n1029) );
XOR2_X1 U955 ( .A(n1226), .B(n1227), .Z(n1078) );
XOR2_X1 U956 ( .A(n1228), .B(n1204), .Z(n1227) );
XNOR2_X1 U957 ( .A(G146), .B(n1050), .ZN(n1204) );
XOR2_X1 U958 ( .A(G125), .B(G140), .Z(n1050) );
NAND3_X1 U959 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
NAND2_X1 U960 ( .A1(KEYINPUT47), .A2(G122), .ZN(n1231) );
NAND3_X1 U961 ( .A1(n1232), .A2(n1233), .A3(G113), .ZN(n1230) );
NAND2_X1 U962 ( .A1(n1234), .A2(n1176), .ZN(n1229) );
INV_X1 U963 ( .A(G113), .ZN(n1176) );
NAND2_X1 U964 ( .A1(n1235), .A2(n1233), .ZN(n1234) );
INV_X1 U965 ( .A(KEYINPUT47), .ZN(n1233) );
XOR2_X1 U966 ( .A(n1232), .B(KEYINPUT42), .Z(n1235) );
XOR2_X1 U967 ( .A(n1236), .B(n1237), .Z(n1226) );
NOR2_X1 U968 ( .A1(KEYINPUT3), .A2(n1238), .ZN(n1237) );
XOR2_X1 U969 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U970 ( .A(n1241), .B(G131), .Z(n1239) );
NAND2_X1 U971 ( .A1(G214), .A2(n1223), .ZN(n1241) );
NOR2_X1 U972 ( .A1(G953), .A2(G237), .ZN(n1223) );
XNOR2_X1 U973 ( .A(G104), .B(KEYINPUT22), .ZN(n1236) );
NAND2_X1 U974 ( .A1(KEYINPUT28), .A2(n1028), .ZN(n1225) );
INV_X1 U975 ( .A(G475), .ZN(n1028) );
XNOR2_X1 U976 ( .A(n1019), .B(n1242), .ZN(n1146) );
NOR2_X1 U977 ( .A1(G478), .A2(KEYINPUT18), .ZN(n1242) );
NOR2_X1 U978 ( .A1(n1075), .A2(G902), .ZN(n1019) );
XOR2_X1 U979 ( .A(n1243), .B(n1244), .Z(n1075) );
XOR2_X1 U980 ( .A(n1245), .B(n1246), .Z(n1244) );
NAND2_X1 U981 ( .A1(KEYINPUT30), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U982 ( .A(G107), .B(n1248), .ZN(n1247) );
NAND2_X1 U983 ( .A1(n1249), .A2(KEYINPUT1), .ZN(n1248) );
XOR2_X1 U984 ( .A(n1232), .B(n1250), .Z(n1249) );
NOR2_X1 U985 ( .A1(G116), .A2(KEYINPUT50), .ZN(n1250) );
XOR2_X1 U986 ( .A(n1251), .B(n1252), .Z(n1243) );
XOR2_X1 U987 ( .A(G134), .B(G128), .Z(n1252) );
NAND3_X1 U988 ( .A1(n1207), .A2(n1035), .A3(G217), .ZN(n1251) );
XNOR2_X1 U989 ( .A(G234), .B(KEYINPUT63), .ZN(n1207) );
XOR2_X1 U990 ( .A(n1009), .B(KEYINPUT48), .Z(n1179) );
NAND2_X1 U991 ( .A1(n1154), .A2(n1018), .ZN(n1009) );
INV_X1 U992 ( .A(n1007), .ZN(n1018) );
XOR2_X1 U993 ( .A(n1253), .B(n1115), .Z(n1007) );
AND2_X1 U994 ( .A1(G210), .A2(n1254), .ZN(n1115) );
NAND2_X1 U995 ( .A1(n1255), .A2(n1183), .ZN(n1253) );
INV_X1 U996 ( .A(G902), .ZN(n1183) );
XOR2_X1 U997 ( .A(n1256), .B(n1108), .Z(n1255) );
XOR2_X1 U998 ( .A(n1058), .B(n1257), .Z(n1108) );
NOR2_X1 U999 ( .A1(KEYINPUT17), .A2(n1059), .ZN(n1257) );
XNOR2_X1 U1000 ( .A(n1258), .B(G113), .ZN(n1059) );
NAND2_X1 U1001 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND2_X1 U1002 ( .A1(G119), .A2(n1261), .ZN(n1260) );
XOR2_X1 U1003 ( .A(KEYINPUT55), .B(n1262), .Z(n1259) );
NOR2_X1 U1004 ( .A1(G119), .A2(n1261), .ZN(n1262) );
XOR2_X1 U1005 ( .A(KEYINPUT2), .B(G116), .Z(n1261) );
XOR2_X1 U1006 ( .A(n1263), .B(n1264), .Z(n1058) );
XOR2_X1 U1007 ( .A(n1232), .B(n1265), .Z(n1264) );
XNOR2_X1 U1008 ( .A(KEYINPUT57), .B(KEYINPUT44), .ZN(n1265) );
INV_X1 U1009 ( .A(G122), .ZN(n1232) );
XNOR2_X1 U1010 ( .A(G110), .B(n1190), .ZN(n1263) );
XNOR2_X1 U1011 ( .A(n1266), .B(n1267), .ZN(n1190) );
XOR2_X1 U1012 ( .A(G104), .B(G101), .Z(n1267) );
XNOR2_X1 U1013 ( .A(G107), .B(KEYINPUT25), .ZN(n1266) );
NAND2_X1 U1014 ( .A1(n1268), .A2(KEYINPUT6), .ZN(n1256) );
XOR2_X1 U1015 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U1016 ( .A(KEYINPUT21), .B(n1113), .ZN(n1270) );
NAND2_X1 U1017 ( .A1(G224), .A2(n1035), .ZN(n1113) );
INV_X1 U1018 ( .A(G953), .ZN(n1035) );
NAND2_X1 U1019 ( .A1(KEYINPUT36), .A2(n1114), .ZN(n1269) );
XOR2_X1 U1020 ( .A(n1091), .B(G125), .Z(n1114) );
XOR2_X1 U1021 ( .A(n1193), .B(n1271), .Z(n1091) );
NOR2_X1 U1022 ( .A1(G128), .A2(KEYINPUT7), .ZN(n1271) );
XOR2_X1 U1023 ( .A(G146), .B(n1240), .Z(n1193) );
INV_X1 U1024 ( .A(n1246), .ZN(n1240) );
XNOR2_X1 U1025 ( .A(G143), .B(KEYINPUT59), .ZN(n1246) );
XNOR2_X1 U1026 ( .A(n1008), .B(KEYINPUT52), .ZN(n1154) );
AND2_X1 U1027 ( .A1(G214), .A2(n1254), .ZN(n1008) );
OR2_X1 U1028 ( .A1(G902), .A2(G237), .ZN(n1254) );
endmodule


