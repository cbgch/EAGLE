//Key = 1001000010011001100100110011110111001111100101110010000011100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U736 ( .A(G107), .B(n1023), .Z(G9) );
NOR2_X1 U737 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025) );
XOR2_X1 U739 ( .A(n1030), .B(KEYINPUT20), .Z(n1029) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U741 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND3_X1 U743 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
XOR2_X1 U744 ( .A(n1040), .B(KEYINPUT40), .Z(n1039) );
NAND3_X1 U745 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1035) );
NAND4_X1 U746 ( .A1(n1044), .A2(n1045), .A3(n1042), .A4(n1046), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
INV_X1 U748 ( .A(n1049), .ZN(n1048) );
NAND3_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
INV_X1 U750 ( .A(n1053), .ZN(n1044) );
NOR2_X1 U751 ( .A1(n1054), .A2(n1055), .ZN(n1028) );
NOR2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
AND2_X1 U753 ( .A1(n1058), .A2(n1033), .ZN(n1057) );
NOR3_X1 U754 ( .A1(n1053), .A2(n1059), .A3(n1040), .ZN(n1056) );
NOR2_X1 U755 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
AND3_X1 U757 ( .A1(n1052), .A2(n1064), .A3(n1065), .ZN(n1060) );
NAND3_X1 U758 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1026) );
NAND3_X1 U759 ( .A1(n1045), .A2(n1069), .A3(n1033), .ZN(n1068) );
NOR3_X1 U760 ( .A1(n1070), .A2(n1063), .A3(n1053), .ZN(n1033) );
NOR3_X1 U761 ( .A1(n1071), .A2(G953), .A3(G952), .ZN(n1024) );
INV_X1 U762 ( .A(n1066), .ZN(n1071) );
NAND4_X1 U763 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1066) );
NOR4_X1 U764 ( .A1(n1076), .A2(n1051), .A3(n1043), .A4(n1077), .ZN(n1075) );
XNOR2_X1 U765 ( .A(n1078), .B(KEYINPUT57), .ZN(n1077) );
NOR2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
AND2_X1 U770 ( .A1(n1083), .A2(KEYINPUT10), .ZN(n1086) );
NOR4_X1 U771 ( .A1(KEYINPUT10), .A2(n1085), .A3(n1083), .A4(n1084), .ZN(n1079) );
INV_X1 U772 ( .A(KEYINPUT31), .ZN(n1084) );
NOR2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1074) );
XOR2_X1 U774 ( .A(n1089), .B(n1090), .Z(n1072) );
NAND2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(G72) );
NAND2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U777 ( .A1(G953), .A2(n1095), .ZN(n1094) );
INV_X1 U778 ( .A(n1096), .ZN(n1093) );
NAND3_X1 U779 ( .A1(G953), .A2(n1097), .A3(n1096), .ZN(n1091) );
XOR2_X1 U780 ( .A(n1098), .B(n1099), .Z(n1096) );
NOR3_X1 U781 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NOR2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
INV_X1 U783 ( .A(n1105), .ZN(n1104) );
XNOR2_X1 U784 ( .A(KEYINPUT25), .B(n1106), .ZN(n1103) );
XOR2_X1 U785 ( .A(KEYINPUT41), .B(n1107), .Z(n1100) );
NOR2_X1 U786 ( .A1(n1105), .A2(n1108), .ZN(n1107) );
XOR2_X1 U787 ( .A(KEYINPUT25), .B(n1106), .Z(n1108) );
XOR2_X1 U788 ( .A(n1109), .B(n1110), .Z(n1105) );
XOR2_X1 U789 ( .A(n1111), .B(G131), .Z(n1109) );
NAND2_X1 U790 ( .A1(n1112), .A2(KEYINPUT38), .ZN(n1111) );
XOR2_X1 U791 ( .A(G137), .B(n1113), .Z(n1112) );
NAND2_X1 U792 ( .A1(n1067), .A2(n1114), .ZN(n1098) );
NAND4_X1 U793 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1114) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1097) );
XOR2_X1 U795 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U798 ( .A(KEYINPUT44), .B(G953), .Z(n1124) );
NAND2_X1 U799 ( .A1(G953), .A2(n1125), .ZN(n1121) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1125) );
NAND2_X1 U801 ( .A1(n1126), .A2(n1127), .ZN(n1119) );
INV_X1 U802 ( .A(n1128), .ZN(n1127) );
NOR2_X1 U803 ( .A1(n1129), .A2(n1130), .ZN(G66) );
NOR3_X1 U804 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
NOR4_X1 U805 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
NOR2_X1 U806 ( .A1(n1138), .A2(n1139), .ZN(n1132) );
NOR3_X1 U807 ( .A1(n1135), .A2(n1140), .A3(n1136), .ZN(n1138) );
INV_X1 U808 ( .A(KEYINPUT47), .ZN(n1135) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1141), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U811 ( .A1(n1144), .A2(n1137), .ZN(n1143) );
INV_X1 U812 ( .A(G478), .ZN(n1144) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1145), .ZN(G60) );
XOR2_X1 U814 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U815 ( .A1(n1148), .A2(n1137), .ZN(n1146) );
INV_X1 U816 ( .A(G475), .ZN(n1148) );
XNOR2_X1 U817 ( .A(G104), .B(n1149), .ZN(G6) );
OR2_X1 U818 ( .A1(n1062), .A2(n1150), .ZN(n1149) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1151), .ZN(G57) );
XOR2_X1 U820 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U821 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U822 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U823 ( .A1(n1158), .A2(n1137), .ZN(n1157) );
INV_X1 U824 ( .A(G472), .ZN(n1158) );
XOR2_X1 U825 ( .A(n1159), .B(n1160), .Z(n1152) );
XNOR2_X1 U826 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U827 ( .A1(KEYINPUT59), .A2(n1163), .ZN(n1162) );
NOR2_X1 U828 ( .A1(KEYINPUT21), .A2(n1164), .ZN(n1161) );
XOR2_X1 U829 ( .A(n1165), .B(KEYINPUT28), .Z(n1159) );
NOR2_X1 U830 ( .A1(n1129), .A2(n1166), .ZN(G54) );
XOR2_X1 U831 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U832 ( .A1(n1169), .A2(n1137), .ZN(n1168) );
INV_X1 U833 ( .A(G469), .ZN(n1169) );
NAND2_X1 U834 ( .A1(KEYINPUT0), .A2(n1170), .ZN(n1167) );
XOR2_X1 U835 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND2_X1 U837 ( .A1(n1164), .A2(n1175), .ZN(n1174) );
NAND2_X1 U838 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U839 ( .A1(KEYINPUT9), .A2(KEYINPUT3), .ZN(n1177) );
NAND3_X1 U840 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1173) );
INV_X1 U841 ( .A(KEYINPUT9), .ZN(n1180) );
NAND2_X1 U842 ( .A1(KEYINPUT3), .A2(n1181), .ZN(n1179) );
NAND2_X1 U843 ( .A1(n1176), .A2(n1182), .ZN(n1181) );
NAND2_X1 U844 ( .A1(n1176), .A2(n1183), .ZN(n1178) );
INV_X1 U845 ( .A(KEYINPUT3), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1129), .A2(n1184), .ZN(G51) );
XOR2_X1 U847 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND3_X1 U848 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NAND2_X1 U849 ( .A1(KEYINPUT7), .A2(n1126), .ZN(n1189) );
OR3_X1 U850 ( .A1(n1126), .A2(KEYINPUT7), .A3(n1190), .ZN(n1188) );
NAND2_X1 U851 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
INV_X1 U853 ( .A(KEYINPUT7), .ZN(n1193) );
XNOR2_X1 U854 ( .A(KEYINPUT1), .B(n1126), .ZN(n1192) );
XOR2_X1 U855 ( .A(n1194), .B(n1195), .Z(n1190) );
XOR2_X1 U856 ( .A(n1196), .B(KEYINPUT24), .Z(n1194) );
NAND3_X1 U857 ( .A1(n1197), .A2(n1198), .A3(n1083), .ZN(n1185) );
NAND2_X1 U858 ( .A1(n1137), .A2(n1199), .ZN(n1198) );
INV_X1 U859 ( .A(KEYINPUT51), .ZN(n1199) );
NAND2_X1 U860 ( .A1(G902), .A2(n1027), .ZN(n1137) );
NAND2_X1 U861 ( .A1(KEYINPUT51), .A2(n1200), .ZN(n1197) );
NAND2_X1 U862 ( .A1(n1140), .A2(G902), .ZN(n1200) );
INV_X1 U863 ( .A(n1027), .ZN(n1140) );
NAND3_X1 U864 ( .A1(n1123), .A2(n1201), .A3(n1202), .ZN(n1027) );
AND3_X1 U865 ( .A1(n1116), .A2(n1118), .A3(n1117), .ZN(n1202) );
NAND2_X1 U866 ( .A1(n1045), .A2(n1203), .ZN(n1117) );
NAND2_X1 U867 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
INV_X1 U868 ( .A(n1206), .ZN(n1205) );
XOR2_X1 U869 ( .A(KEYINPUT27), .B(n1207), .Z(n1204) );
INV_X1 U870 ( .A(n1208), .ZN(n1118) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1058), .ZN(n1116) );
XOR2_X1 U872 ( .A(KEYINPUT55), .B(n1115), .Z(n1201) );
AND3_X1 U873 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1115) );
NAND4_X1 U874 ( .A1(n1045), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1212) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U876 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U877 ( .A1(n1069), .A2(n1220), .ZN(n1219) );
XOR2_X1 U878 ( .A(n1221), .B(KEYINPUT48), .Z(n1216) );
NAND2_X1 U879 ( .A1(n1222), .A2(n1223), .ZN(n1214) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1220), .ZN(n1222) );
INV_X1 U881 ( .A(KEYINPUT19), .ZN(n1220) );
AND4_X1 U882 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1123) );
AND4_X1 U883 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
OR2_X1 U884 ( .A1(n1150), .A2(n1232), .ZN(n1231) );
XOR2_X1 U885 ( .A(KEYINPUT58), .B(n1218), .Z(n1232) );
NOR2_X1 U886 ( .A1(n1233), .A2(n1023), .ZN(n1226) );
NOR2_X1 U887 ( .A1(n1221), .A2(n1150), .ZN(n1023) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1042), .ZN(n1150) );
NOR2_X1 U889 ( .A1(n1067), .A2(G952), .ZN(n1129) );
XOR2_X1 U890 ( .A(G146), .B(n1208), .Z(G48) );
NOR3_X1 U891 ( .A1(n1235), .A2(n1236), .A3(n1062), .ZN(n1208) );
XOR2_X1 U892 ( .A(G143), .B(n1237), .Z(G45) );
NOR3_X1 U893 ( .A1(n1238), .A2(KEYINPUT60), .A3(n1236), .ZN(n1237) );
XOR2_X1 U894 ( .A(KEYINPUT37), .B(n1209), .Z(n1238) );
AND4_X1 U895 ( .A1(n1069), .A2(n1213), .A3(n1088), .A4(n1078), .ZN(n1209) );
XNOR2_X1 U896 ( .A(G140), .B(n1239), .ZN(G42) );
NAND2_X1 U897 ( .A1(n1045), .A2(n1207), .ZN(n1239) );
AND2_X1 U898 ( .A1(n1240), .A2(n1213), .ZN(n1207) );
XNOR2_X1 U899 ( .A(G137), .B(n1241), .ZN(G39) );
NAND2_X1 U900 ( .A1(n1242), .A2(n1206), .ZN(n1241) );
NOR2_X1 U901 ( .A1(n1070), .A2(n1235), .ZN(n1206) );
INV_X1 U902 ( .A(n1052), .ZN(n1070) );
XOR2_X1 U903 ( .A(n1040), .B(KEYINPUT39), .Z(n1242) );
XOR2_X1 U904 ( .A(G134), .B(n1243), .Z(G36) );
NOR2_X1 U905 ( .A1(n1221), .A2(n1244), .ZN(n1243) );
XOR2_X1 U906 ( .A(G131), .B(n1245), .Z(G33) );
NOR2_X1 U907 ( .A1(n1062), .A2(n1244), .ZN(n1245) );
NAND3_X1 U908 ( .A1(n1069), .A2(n1213), .A3(n1045), .ZN(n1244) );
INV_X1 U909 ( .A(n1040), .ZN(n1045) );
NAND2_X1 U910 ( .A1(n1041), .A2(n1246), .ZN(n1040) );
NAND3_X1 U911 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(G30) );
NAND2_X1 U912 ( .A1(KEYINPUT14), .A2(n1211), .ZN(n1249) );
INV_X1 U913 ( .A(n1250), .ZN(n1211) );
NAND3_X1 U914 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1248) );
NAND2_X1 U915 ( .A1(G128), .A2(n1253), .ZN(n1247) );
NAND2_X1 U916 ( .A1(n1254), .A2(n1251), .ZN(n1253) );
INV_X1 U917 ( .A(KEYINPUT14), .ZN(n1251) );
XOR2_X1 U918 ( .A(KEYINPUT6), .B(n1250), .Z(n1254) );
NOR3_X1 U919 ( .A1(n1221), .A2(n1236), .A3(n1235), .ZN(n1250) );
NAND3_X1 U920 ( .A1(n1255), .A2(n1037), .A3(n1213), .ZN(n1235) );
AND3_X1 U921 ( .A1(n1064), .A2(n1256), .A3(n1065), .ZN(n1213) );
INV_X1 U922 ( .A(n1058), .ZN(n1236) );
XOR2_X1 U923 ( .A(n1165), .B(n1230), .Z(G3) );
NAND3_X1 U924 ( .A1(n1069), .A2(n1234), .A3(n1052), .ZN(n1230) );
XNOR2_X1 U925 ( .A(G125), .B(n1210), .ZN(G27) );
NAND4_X1 U926 ( .A1(n1240), .A2(n1257), .A3(n1058), .A4(n1256), .ZN(n1210) );
NAND2_X1 U927 ( .A1(n1053), .A2(n1258), .ZN(n1256) );
NAND2_X1 U928 ( .A1(n1102), .A2(n1259), .ZN(n1258) );
NOR2_X1 U929 ( .A1(n1067), .A2(G900), .ZN(n1102) );
NOR3_X1 U930 ( .A1(n1260), .A2(n1261), .A3(n1062), .ZN(n1240) );
INV_X1 U931 ( .A(n1218), .ZN(n1062) );
XNOR2_X1 U932 ( .A(G122), .B(n1229), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1262), .A2(n1042), .A3(n1088), .A4(n1078), .ZN(n1229) );
INV_X1 U934 ( .A(n1055), .ZN(n1042) );
NAND2_X1 U935 ( .A1(n1038), .A2(n1260), .ZN(n1055) );
XOR2_X1 U936 ( .A(n1228), .B(n1263), .Z(G21) );
XOR2_X1 U937 ( .A(KEYINPUT33), .B(G119), .Z(n1263) );
NAND4_X1 U938 ( .A1(n1262), .A2(n1052), .A3(n1255), .A4(n1037), .ZN(n1228) );
AND3_X1 U939 ( .A1(n1058), .A2(n1264), .A3(n1257), .ZN(n1262) );
XOR2_X1 U940 ( .A(G116), .B(n1233), .Z(G18) );
AND4_X1 U941 ( .A1(n1049), .A2(n1069), .A3(n1058), .A4(n1264), .ZN(n1233) );
NOR2_X1 U942 ( .A1(n1063), .A2(n1221), .ZN(n1049) );
NAND2_X1 U943 ( .A1(n1265), .A2(n1078), .ZN(n1221) );
XOR2_X1 U944 ( .A(KEYINPUT63), .B(n1088), .Z(n1265) );
INV_X1 U945 ( .A(n1257), .ZN(n1063) );
XOR2_X1 U946 ( .A(n1266), .B(n1224), .Z(G15) );
NAND4_X1 U947 ( .A1(n1069), .A2(n1257), .A3(n1218), .A4(n1267), .ZN(n1224) );
NOR2_X1 U948 ( .A1(n1078), .A2(n1268), .ZN(n1218) );
NOR2_X1 U949 ( .A1(n1064), .A2(n1051), .ZN(n1257) );
INV_X1 U950 ( .A(n1223), .ZN(n1069) );
NAND2_X1 U951 ( .A1(n1255), .A2(n1260), .ZN(n1223) );
XOR2_X1 U952 ( .A(n1261), .B(KEYINPUT42), .Z(n1255) );
XNOR2_X1 U953 ( .A(G110), .B(n1225), .ZN(G12) );
NAND4_X1 U954 ( .A1(n1052), .A2(n1037), .A3(n1234), .A4(n1038), .ZN(n1225) );
INV_X1 U955 ( .A(n1261), .ZN(n1038) );
XOR2_X1 U956 ( .A(n1073), .B(KEYINPUT15), .Z(n1261) );
XOR2_X1 U957 ( .A(n1269), .B(G472), .Z(n1073) );
NAND2_X1 U958 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XNOR2_X1 U959 ( .A(n1272), .B(n1163), .ZN(n1270) );
NAND3_X1 U960 ( .A1(n1273), .A2(n1067), .A3(G210), .ZN(n1163) );
XOR2_X1 U961 ( .A(n1274), .B(G101), .Z(n1272) );
NAND3_X1 U962 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1274) );
NAND2_X1 U963 ( .A1(n1156), .A2(n1278), .ZN(n1277) );
INV_X1 U964 ( .A(KEYINPUT23), .ZN(n1278) );
NAND3_X1 U965 ( .A1(KEYINPUT23), .A2(n1279), .A3(n1280), .ZN(n1276) );
OR2_X1 U966 ( .A1(n1280), .A2(n1279), .ZN(n1275) );
NOR2_X1 U967 ( .A1(KEYINPUT2), .A2(n1156), .ZN(n1279) );
XOR2_X1 U968 ( .A(n1281), .B(n1282), .Z(n1156) );
XOR2_X1 U969 ( .A(G116), .B(n1283), .Z(n1282) );
NOR2_X1 U970 ( .A1(G113), .A2(KEYINPUT13), .ZN(n1283) );
NAND2_X1 U971 ( .A1(KEYINPUT43), .A2(G119), .ZN(n1281) );
XNOR2_X1 U972 ( .A(n1284), .B(n1154), .ZN(n1280) );
XOR2_X1 U973 ( .A(n1182), .B(KEYINPUT8), .Z(n1284) );
AND3_X1 U974 ( .A1(n1065), .A2(n1064), .A3(n1267), .ZN(n1234) );
AND2_X1 U975 ( .A1(n1285), .A2(n1264), .ZN(n1267) );
NAND2_X1 U976 ( .A1(n1053), .A2(n1286), .ZN(n1264) );
NAND2_X1 U977 ( .A1(n1259), .A2(n1128), .ZN(n1286) );
NOR2_X1 U978 ( .A1(n1067), .A2(G898), .ZN(n1128) );
AND2_X1 U979 ( .A1(n1287), .A2(n1288), .ZN(n1259) );
XOR2_X1 U980 ( .A(n1271), .B(KEYINPUT46), .Z(n1287) );
NAND3_X1 U981 ( .A1(n1288), .A2(n1067), .A3(G952), .ZN(n1053) );
NAND2_X1 U982 ( .A1(G237), .A2(G234), .ZN(n1288) );
XOR2_X1 U983 ( .A(KEYINPUT34), .B(n1058), .Z(n1285) );
NOR2_X1 U984 ( .A1(n1041), .A2(n1043), .ZN(n1058) );
INV_X1 U985 ( .A(n1246), .ZN(n1043) );
NAND2_X1 U986 ( .A1(G214), .A2(n1289), .ZN(n1246) );
XNOR2_X1 U987 ( .A(n1085), .B(n1083), .ZN(n1041) );
AND2_X1 U988 ( .A1(G210), .A2(n1289), .ZN(n1083) );
NAND2_X1 U989 ( .A1(n1273), .A2(n1271), .ZN(n1289) );
AND2_X1 U990 ( .A1(n1290), .A2(n1271), .ZN(n1085) );
XOR2_X1 U991 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U992 ( .A(n1126), .B(n1293), .Z(n1292) );
NOR2_X1 U993 ( .A1(KEYINPUT18), .A2(n1195), .ZN(n1293) );
XOR2_X1 U994 ( .A(G125), .B(n1154), .Z(n1195) );
XOR2_X1 U995 ( .A(n1294), .B(n1295), .Z(n1126) );
XOR2_X1 U996 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U997 ( .A(n1298), .B(n1299), .ZN(n1297) );
NAND2_X1 U998 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND2_X1 U999 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U1000 ( .A1(KEYINPUT32), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1001 ( .A1(KEYINPUT11), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1002 ( .A1(G107), .A2(n1306), .ZN(n1300) );
NAND2_X1 U1003 ( .A1(KEYINPUT11), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1004 ( .A1(KEYINPUT32), .A2(n1308), .ZN(n1307) );
XOR2_X1 U1005 ( .A(n1309), .B(n1310), .Z(n1294) );
XOR2_X1 U1006 ( .A(G113), .B(G101), .Z(n1310) );
NAND2_X1 U1007 ( .A1(KEYINPUT50), .A2(G119), .ZN(n1309) );
XOR2_X1 U1008 ( .A(n1196), .B(KEYINPUT30), .Z(n1291) );
NAND2_X1 U1009 ( .A1(G224), .A2(n1067), .ZN(n1196) );
INV_X1 U1010 ( .A(n1050), .ZN(n1064) );
XNOR2_X1 U1011 ( .A(n1087), .B(KEYINPUT52), .ZN(n1050) );
XNOR2_X1 U1012 ( .A(n1311), .B(G469), .ZN(n1087) );
NAND2_X1 U1013 ( .A1(n1312), .A2(n1271), .ZN(n1311) );
XOR2_X1 U1014 ( .A(n1172), .B(n1313), .Z(n1312) );
XOR2_X1 U1015 ( .A(n1176), .B(n1164), .Z(n1313) );
INV_X1 U1016 ( .A(n1182), .ZN(n1164) );
XOR2_X1 U1017 ( .A(n1314), .B(G131), .Z(n1182) );
NAND3_X1 U1018 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1314) );
NAND2_X1 U1019 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1020 ( .A1(KEYINPUT45), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1021 ( .A(KEYINPUT36), .B(G137), .ZN(n1318) );
NAND4_X1 U1022 ( .A1(n1320), .A2(n1321), .A3(KEYINPUT45), .A4(n1322), .ZN(n1316) );
XOR2_X1 U1023 ( .A(KEYINPUT36), .B(G137), .Z(n1321) );
OR2_X1 U1024 ( .A1(n1320), .A2(n1322), .ZN(n1315) );
INV_X1 U1025 ( .A(KEYINPUT4), .ZN(n1322) );
XOR2_X1 U1026 ( .A(n1113), .B(KEYINPUT26), .Z(n1320) );
XOR2_X1 U1027 ( .A(n1323), .B(n1324), .Z(n1176) );
XOR2_X1 U1028 ( .A(n1308), .B(n1110), .Z(n1324) );
XNOR2_X1 U1029 ( .A(n1154), .B(KEYINPUT17), .ZN(n1110) );
XNOR2_X1 U1030 ( .A(G143), .B(n1325), .ZN(n1154) );
INV_X1 U1031 ( .A(n1302), .ZN(n1308) );
XOR2_X1 U1032 ( .A(n1165), .B(n1326), .Z(n1323) );
XOR2_X1 U1033 ( .A(KEYINPUT49), .B(G107), .Z(n1326) );
INV_X1 U1034 ( .A(G101), .ZN(n1165) );
XNOR2_X1 U1035 ( .A(n1299), .B(n1327), .ZN(n1172) );
XOR2_X1 U1036 ( .A(G140), .B(n1328), .Z(n1327) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1095), .ZN(n1328) );
INV_X1 U1038 ( .A(G227), .ZN(n1095) );
XNOR2_X1 U1039 ( .A(n1051), .B(KEYINPUT35), .ZN(n1065) );
AND2_X1 U1040 ( .A1(n1329), .A2(n1330), .ZN(n1051) );
XOR2_X1 U1041 ( .A(KEYINPUT5), .B(G221), .Z(n1329) );
INV_X1 U1042 ( .A(n1260), .ZN(n1037) );
NAND3_X1 U1043 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1260) );
OR2_X1 U1044 ( .A1(n1131), .A2(KEYINPUT29), .ZN(n1333) );
INV_X1 U1045 ( .A(n1089), .ZN(n1131) );
NAND3_X1 U1046 ( .A1(KEYINPUT29), .A2(n1090), .A3(n1334), .ZN(n1332) );
OR2_X1 U1047 ( .A1(n1334), .A2(n1090), .ZN(n1331) );
INV_X1 U1048 ( .A(n1136), .ZN(n1090) );
NAND2_X1 U1049 ( .A1(G217), .A2(n1330), .ZN(n1136) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1271), .ZN(n1330) );
NOR2_X1 U1051 ( .A1(KEYINPUT53), .A2(n1089), .ZN(n1334) );
NAND2_X1 U1052 ( .A1(n1134), .A2(n1271), .ZN(n1089) );
INV_X1 U1053 ( .A(n1139), .ZN(n1134) );
XOR2_X1 U1054 ( .A(n1335), .B(n1336), .Z(n1139) );
XOR2_X1 U1055 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1056 ( .A(G119), .B(G137), .ZN(n1338) );
NAND2_X1 U1057 ( .A1(G221), .A2(n1339), .ZN(n1337) );
XNOR2_X1 U1058 ( .A(n1325), .B(n1340), .ZN(n1335) );
XOR2_X1 U1059 ( .A(n1299), .B(n1106), .Z(n1340) );
XOR2_X1 U1060 ( .A(G110), .B(KEYINPUT54), .Z(n1299) );
XNOR2_X1 U1061 ( .A(n1341), .B(G128), .ZN(n1325) );
INV_X1 U1062 ( .A(G146), .ZN(n1341) );
NOR2_X1 U1063 ( .A1(n1078), .A2(n1088), .ZN(n1052) );
INV_X1 U1064 ( .A(n1268), .ZN(n1088) );
XOR2_X1 U1065 ( .A(n1342), .B(G475), .Z(n1268) );
OR2_X1 U1066 ( .A1(n1147), .A2(G902), .ZN(n1342) );
XNOR2_X1 U1067 ( .A(n1343), .B(n1344), .ZN(n1147) );
XOR2_X1 U1068 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1069 ( .A(G131), .B(G122), .Z(n1346) );
XOR2_X1 U1070 ( .A(KEYINPUT61), .B(G146), .Z(n1345) );
XOR2_X1 U1071 ( .A(n1347), .B(n1348), .Z(n1343) );
XOR2_X1 U1072 ( .A(n1266), .B(n1349), .Z(n1348) );
NAND2_X1 U1073 ( .A1(KEYINPUT12), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1074 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND2_X1 U1075 ( .A1(KEYINPUT56), .A2(n1353), .ZN(n1352) );
INV_X1 U1076 ( .A(G143), .ZN(n1353) );
NAND3_X1 U1077 ( .A1(n1273), .A2(n1067), .A3(G214), .ZN(n1351) );
INV_X1 U1078 ( .A(G237), .ZN(n1273) );
INV_X1 U1079 ( .A(G113), .ZN(n1266) );
XOR2_X1 U1080 ( .A(n1302), .B(n1106), .Z(n1347) );
XOR2_X1 U1081 ( .A(G125), .B(G140), .Z(n1106) );
XNOR2_X1 U1082 ( .A(G104), .B(KEYINPUT62), .ZN(n1302) );
XNOR2_X1 U1083 ( .A(n1354), .B(G478), .ZN(n1078) );
NAND2_X1 U1084 ( .A1(n1142), .A2(n1271), .ZN(n1354) );
INV_X1 U1085 ( .A(G902), .ZN(n1271) );
XNOR2_X1 U1086 ( .A(n1355), .B(n1356), .ZN(n1142) );
XOR2_X1 U1087 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1088 ( .A(n1305), .B(G143), .Z(n1358) );
INV_X1 U1089 ( .A(G107), .ZN(n1305) );
NAND2_X1 U1090 ( .A1(KEYINPUT16), .A2(n1252), .ZN(n1357) );
INV_X1 U1091 ( .A(G128), .ZN(n1252) );
XOR2_X1 U1092 ( .A(n1359), .B(n1296), .Z(n1355) );
XOR2_X1 U1093 ( .A(G116), .B(G122), .Z(n1296) );
XOR2_X1 U1094 ( .A(n1360), .B(n1361), .Z(n1359) );
INV_X1 U1095 ( .A(n1113), .ZN(n1361) );
XNOR2_X1 U1096 ( .A(G134), .B(KEYINPUT22), .ZN(n1113) );
NAND2_X1 U1097 ( .A1(G217), .A2(n1339), .ZN(n1360) );
AND2_X1 U1098 ( .A1(G234), .A2(n1067), .ZN(n1339) );
INV_X1 U1099 ( .A(G953), .ZN(n1067) );
endmodule


