//Key = 0100100110111001111101010101110001100011010110101110011101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345;

XNOR2_X1 U742 ( .A(n1022), .B(n1023), .ZN(G9) );
NOR2_X1 U743 ( .A1(KEYINPUT3), .A2(n1024), .ZN(n1023) );
NOR2_X1 U744 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U746 ( .A(n1031), .B(KEYINPUT27), .Z(n1030) );
NAND4_X1 U747 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR3_X1 U748 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1029) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
AND3_X1 U754 ( .A1(n1049), .A2(n1050), .A3(G214), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
AND3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1039) );
NAND3_X1 U759 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1027) );
NAND3_X1 U760 ( .A1(n1063), .A2(n1064), .A3(n1033), .ZN(n1062) );
NOR3_X1 U761 ( .A1(n1052), .A2(n1046), .A3(n1036), .ZN(n1033) );
OR2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR3_X1 U763 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1025) );
INV_X1 U764 ( .A(n1060), .ZN(n1067) );
NAND4_X1 U765 ( .A1(n1063), .A2(n1057), .A3(n1068), .A4(n1069), .ZN(n1060) );
NOR4_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1055), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1073), .B(KEYINPUT16), .Z(n1071) );
NOR2_X1 U768 ( .A1(G475), .A2(n1074), .ZN(n1070) );
XOR2_X1 U769 ( .A(n1075), .B(G478), .Z(n1068) );
XOR2_X1 U770 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1082), .B(n1083), .Z(n1081) );
XNOR2_X1 U774 ( .A(n1084), .B(n1085), .ZN(n1083) );
XOR2_X1 U775 ( .A(n1086), .B(G125), .Z(n1082) );
NAND3_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND2_X1 U777 ( .A1(G134), .A2(n1090), .ZN(n1089) );
NAND2_X1 U778 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
INV_X1 U779 ( .A(KEYINPUT12), .ZN(n1092) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
INV_X1 U781 ( .A(G134), .ZN(n1094) );
XNOR2_X1 U782 ( .A(KEYINPUT2), .B(n1090), .ZN(n1093) );
NAND2_X1 U783 ( .A1(KEYINPUT12), .A2(n1095), .ZN(n1087) );
NAND2_X1 U784 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
OR3_X1 U785 ( .A1(n1090), .A2(G134), .A3(KEYINPUT2), .ZN(n1097) );
NAND2_X1 U786 ( .A1(KEYINPUT2), .A2(n1090), .ZN(n1096) );
XNOR2_X1 U787 ( .A(n1098), .B(KEYINPUT25), .ZN(n1090) );
INV_X1 U788 ( .A(G137), .ZN(n1098) );
NOR2_X1 U789 ( .A1(G900), .A2(n1061), .ZN(n1080) );
NAND2_X1 U790 ( .A1(n1099), .A2(n1061), .ZN(n1078) );
NAND2_X1 U791 ( .A1(G953), .A2(n1100), .ZN(n1076) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1100) );
XOR2_X1 U793 ( .A(n1101), .B(n1102), .Z(G69) );
XOR2_X1 U794 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U796 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1107) );
NAND2_X1 U798 ( .A1(KEYINPUT59), .A2(n1111), .ZN(n1109) );
NOR2_X1 U799 ( .A1(G898), .A2(n1061), .ZN(n1105) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1103) );
XOR2_X1 U801 ( .A(KEYINPUT42), .B(G953), .Z(n1113) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR3_X1 U803 ( .A1(n1061), .A2(KEYINPUT47), .A3(n1116), .ZN(n1101) );
NOR2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XNOR2_X1 U806 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1125), .ZN(G63) );
NOR3_X1 U809 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
NOR3_X1 U810 ( .A1(n1129), .A2(n1130), .A3(n1124), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1130), .ZN(n1132) );
INV_X1 U813 ( .A(n1129), .ZN(n1131) );
NOR3_X1 U814 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(G60) );
NOR3_X1 U815 ( .A1(n1137), .A2(G953), .A3(G952), .ZN(n1136) );
AND2_X1 U816 ( .A1(n1137), .A2(n1119), .ZN(n1135) );
INV_X1 U817 ( .A(KEYINPUT32), .ZN(n1137) );
XNOR2_X1 U818 ( .A(n1138), .B(n1139), .ZN(n1134) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1124), .ZN(n1139) );
INV_X1 U820 ( .A(G475), .ZN(n1140) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(G6) );
NOR2_X1 U822 ( .A1(n1119), .A2(n1143), .ZN(G57) );
XOR2_X1 U823 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U824 ( .A(n1146), .B(n1147), .ZN(n1145) );
XNOR2_X1 U825 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1144) );
XOR2_X1 U827 ( .A(KEYINPUT10), .B(n1152), .Z(n1151) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1124), .ZN(n1152) );
INV_X1 U829 ( .A(G472), .ZN(n1153) );
NAND2_X1 U830 ( .A1(KEYINPUT15), .A2(n1154), .ZN(n1150) );
NOR2_X1 U831 ( .A1(n1119), .A2(n1155), .ZN(G54) );
XOR2_X1 U832 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U834 ( .A1(KEYINPUT13), .A2(n1160), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1161), .B(n1162), .Z(n1156) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1124), .ZN(n1162) );
INV_X1 U837 ( .A(G469), .ZN(n1163) );
NAND2_X1 U838 ( .A1(KEYINPUT48), .A2(n1149), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1061), .A2(G952), .ZN(n1119) );
NOR2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(G51) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1124), .ZN(n1167) );
NAND2_X1 U843 ( .A1(G902), .A2(n1028), .ZN(n1124) );
INV_X1 U844 ( .A(n1133), .ZN(n1028) );
NOR3_X1 U845 ( .A1(n1099), .A2(n1115), .A3(n1169), .ZN(n1133) );
XNOR2_X1 U846 ( .A(n1114), .B(KEYINPUT28), .ZN(n1169) );
NAND3_X1 U847 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1114) );
NAND2_X1 U848 ( .A1(n1048), .A2(n1173), .ZN(n1172) );
NAND2_X1 U849 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND4_X1 U850 ( .A1(n1142), .A2(n1176), .A3(n1177), .A4(n1022), .ZN(n1115) );
NAND3_X1 U851 ( .A1(n1066), .A2(n1059), .A3(n1178), .ZN(n1022) );
NAND3_X1 U852 ( .A1(n1178), .A2(n1059), .A3(n1065), .ZN(n1142) );
NAND4_X1 U853 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1099) );
NOR4_X1 U854 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1181) );
NOR3_X1 U856 ( .A1(n1038), .A2(n1052), .A3(n1189), .ZN(n1188) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1180) );
NAND2_X1 U858 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND3_X1 U859 ( .A1(n1052), .A2(n1194), .A3(n1065), .ZN(n1193) );
INV_X1 U860 ( .A(KEYINPUT38), .ZN(n1194) );
INV_X1 U861 ( .A(n1057), .ZN(n1052) );
NAND3_X1 U862 ( .A1(n1048), .A2(n1195), .A3(n1196), .ZN(n1192) );
NAND2_X1 U863 ( .A1(KEYINPUT38), .A2(n1197), .ZN(n1179) );
NOR2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1166) );
XOR2_X1 U865 ( .A(KEYINPUT31), .B(n1200), .Z(n1199) );
NOR2_X1 U866 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
AND2_X1 U867 ( .A1(n1202), .A2(n1201), .ZN(n1198) );
NOR2_X1 U868 ( .A1(n1061), .A2(n1203), .ZN(n1164) );
XOR2_X1 U869 ( .A(KEYINPUT51), .B(G952), .Z(n1203) );
XOR2_X1 U870 ( .A(G146), .B(n1187), .Z(G48) );
AND3_X1 U871 ( .A1(n1065), .A2(n1048), .A3(n1204), .ZN(n1187) );
XOR2_X1 U872 ( .A(n1205), .B(n1206), .Z(G45) );
NOR2_X1 U873 ( .A1(KEYINPUT37), .A2(n1207), .ZN(n1206) );
INV_X1 U874 ( .A(G143), .ZN(n1207) );
NOR4_X1 U875 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1205) );
XOR2_X1 U876 ( .A(n1212), .B(KEYINPUT26), .Z(n1209) );
XOR2_X1 U877 ( .A(G140), .B(n1186), .Z(G42) );
AND3_X1 U878 ( .A1(n1057), .A2(n1058), .A3(n1213), .ZN(n1186) );
XOR2_X1 U879 ( .A(G137), .B(n1214), .Z(G39) );
NOR3_X1 U880 ( .A1(n1215), .A2(n1189), .A3(n1038), .ZN(n1214) );
XOR2_X1 U881 ( .A(KEYINPUT4), .B(n1057), .Z(n1215) );
XOR2_X1 U882 ( .A(G134), .B(n1185), .Z(G36) );
AND3_X1 U883 ( .A1(n1057), .A2(n1066), .A3(n1190), .ZN(n1185) );
XOR2_X1 U884 ( .A(n1197), .B(n1216), .Z(G33) );
NOR2_X1 U885 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U886 ( .A(KEYINPUT63), .B(KEYINPUT40), .Z(n1218) );
AND3_X1 U887 ( .A1(n1065), .A2(n1057), .A3(n1190), .ZN(n1197) );
INV_X1 U888 ( .A(n1210), .ZN(n1190) );
NAND3_X1 U889 ( .A1(n1058), .A2(n1219), .A3(n1054), .ZN(n1210) );
NOR2_X1 U890 ( .A1(n1220), .A2(n1221), .ZN(n1057) );
AND2_X1 U891 ( .A1(G214), .A2(n1050), .ZN(n1221) );
XOR2_X1 U892 ( .A(G128), .B(n1184), .Z(G30) );
AND3_X1 U893 ( .A1(n1066), .A2(n1048), .A3(n1204), .ZN(n1184) );
INV_X1 U894 ( .A(n1189), .ZN(n1204) );
NAND4_X1 U895 ( .A1(n1222), .A2(n1058), .A3(n1055), .A4(n1219), .ZN(n1189) );
INV_X1 U896 ( .A(n1223), .ZN(n1055) );
XOR2_X1 U897 ( .A(n1176), .B(n1224), .Z(G3) );
NAND2_X1 U898 ( .A1(KEYINPUT8), .A2(G101), .ZN(n1224) );
NAND3_X1 U899 ( .A1(n1054), .A2(n1178), .A3(n1035), .ZN(n1176) );
XOR2_X1 U900 ( .A(n1183), .B(n1225), .Z(G27) );
XOR2_X1 U901 ( .A(KEYINPUT0), .B(G125), .Z(n1225) );
AND3_X1 U902 ( .A1(n1063), .A2(n1048), .A3(n1213), .ZN(n1183) );
AND4_X1 U903 ( .A1(n1222), .A2(n1065), .A3(n1223), .A4(n1219), .ZN(n1213) );
NAND2_X1 U904 ( .A1(n1036), .A2(n1226), .ZN(n1219) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1228), .ZN(n1226) );
INV_X1 U906 ( .A(G900), .ZN(n1228) );
XOR2_X1 U907 ( .A(n1229), .B(n1230), .Z(G24) );
NAND2_X1 U908 ( .A1(n1231), .A2(n1048), .ZN(n1230) );
XOR2_X1 U909 ( .A(n1174), .B(KEYINPUT7), .Z(n1231) );
NAND4_X1 U910 ( .A1(n1232), .A2(n1059), .A3(n1196), .A4(n1195), .ZN(n1174) );
INV_X1 U911 ( .A(n1046), .ZN(n1059) );
NAND2_X1 U912 ( .A1(n1223), .A2(n1056), .ZN(n1046) );
INV_X1 U913 ( .A(n1222), .ZN(n1056) );
XNOR2_X1 U914 ( .A(G119), .B(n1170), .ZN(G21) );
NAND4_X1 U915 ( .A1(n1232), .A2(n1035), .A3(n1233), .A4(n1222), .ZN(n1170) );
NOR2_X1 U916 ( .A1(n1223), .A2(n1212), .ZN(n1233) );
XNOR2_X1 U917 ( .A(G116), .B(n1171), .ZN(G18) );
NAND4_X1 U918 ( .A1(n1232), .A2(n1054), .A3(n1066), .A4(n1048), .ZN(n1171) );
NOR2_X1 U919 ( .A1(n1195), .A2(n1211), .ZN(n1066) );
XOR2_X1 U920 ( .A(G113), .B(n1234), .Z(G15) );
NOR2_X1 U921 ( .A1(n1235), .A2(n1212), .ZN(n1234) );
XOR2_X1 U922 ( .A(n1175), .B(KEYINPUT36), .Z(n1235) );
NAND3_X1 U923 ( .A1(n1054), .A2(n1065), .A3(n1232), .ZN(n1175) );
AND2_X1 U924 ( .A1(n1063), .A2(n1236), .ZN(n1232) );
INV_X1 U925 ( .A(n1042), .ZN(n1063) );
NAND2_X1 U926 ( .A1(n1034), .A2(n1237), .ZN(n1042) );
NOR2_X1 U927 ( .A1(n1196), .A2(n1208), .ZN(n1065) );
NOR2_X1 U928 ( .A1(n1222), .A2(n1223), .ZN(n1054) );
XNOR2_X1 U929 ( .A(G110), .B(n1177), .ZN(G12) );
NAND4_X1 U930 ( .A1(n1222), .A2(n1035), .A3(n1223), .A4(n1178), .ZN(n1177) );
AND3_X1 U931 ( .A1(n1058), .A2(n1236), .A3(n1048), .ZN(n1178) );
INV_X1 U932 ( .A(n1212), .ZN(n1048) );
NAND2_X1 U933 ( .A1(n1220), .A2(n1238), .ZN(n1212) );
NAND2_X1 U934 ( .A1(G214), .A2(n1050), .ZN(n1238) );
INV_X1 U935 ( .A(n1049), .ZN(n1220) );
XNOR2_X1 U936 ( .A(n1239), .B(n1168), .ZN(n1049) );
NAND2_X1 U937 ( .A1(G210), .A2(n1050), .ZN(n1168) );
NAND2_X1 U938 ( .A1(n1240), .A2(n1241), .ZN(n1050) );
XNOR2_X1 U939 ( .A(G237), .B(KEYINPUT6), .ZN(n1240) );
NAND2_X1 U940 ( .A1(n1242), .A2(n1241), .ZN(n1239) );
XNOR2_X1 U941 ( .A(n1243), .B(n1201), .ZN(n1242) );
XNOR2_X1 U942 ( .A(n1146), .B(n1244), .ZN(n1201) );
XOR2_X1 U943 ( .A(G125), .B(n1245), .Z(n1244) );
NOR2_X1 U944 ( .A1(G953), .A2(n1117), .ZN(n1245) );
INV_X1 U945 ( .A(G224), .ZN(n1117) );
XNOR2_X1 U946 ( .A(n1202), .B(KEYINPUT43), .ZN(n1243) );
XOR2_X1 U947 ( .A(n1111), .B(n1246), .Z(n1202) );
XNOR2_X1 U948 ( .A(n1247), .B(n1110), .ZN(n1246) );
XNOR2_X1 U949 ( .A(n1248), .B(n1249), .ZN(n1110) );
NAND2_X1 U950 ( .A1(n1250), .A2(KEYINPUT46), .ZN(n1248) );
XOR2_X1 U951 ( .A(n1229), .B(KEYINPUT30), .Z(n1250) );
NAND2_X1 U952 ( .A1(KEYINPUT61), .A2(n1108), .ZN(n1247) );
XOR2_X1 U953 ( .A(n1251), .B(n1252), .Z(n1108) );
XOR2_X1 U954 ( .A(KEYINPUT23), .B(G107), .Z(n1252) );
XNOR2_X1 U955 ( .A(G101), .B(n1253), .ZN(n1251) );
XOR2_X1 U956 ( .A(n1254), .B(n1255), .Z(n1111) );
NOR2_X1 U957 ( .A1(G113), .A2(KEYINPUT60), .ZN(n1255) );
NAND2_X1 U958 ( .A1(n1036), .A2(n1256), .ZN(n1236) );
NAND4_X1 U959 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1118), .ZN(n1256) );
INV_X1 U960 ( .A(G898), .ZN(n1118) );
NAND3_X1 U961 ( .A1(n1227), .A2(n1061), .A3(n1257), .ZN(n1036) );
XNOR2_X1 U962 ( .A(G952), .B(KEYINPUT49), .ZN(n1257) );
NAND2_X1 U963 ( .A1(G237), .A2(n1258), .ZN(n1227) );
NOR2_X1 U964 ( .A1(n1034), .A2(n1032), .ZN(n1058) );
INV_X1 U965 ( .A(n1237), .ZN(n1032) );
NAND2_X1 U966 ( .A1(G221), .A2(n1259), .ZN(n1237) );
XOR2_X1 U967 ( .A(n1260), .B(G469), .Z(n1034) );
NAND2_X1 U968 ( .A1(n1261), .A2(n1241), .ZN(n1260) );
XOR2_X1 U969 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U970 ( .A(n1159), .B(n1160), .Z(n1263) );
XOR2_X1 U971 ( .A(G140), .B(n1249), .Z(n1160) );
XNOR2_X1 U972 ( .A(n1264), .B(n1265), .ZN(n1159) );
XOR2_X1 U973 ( .A(n1266), .B(n1085), .Z(n1265) );
XOR2_X1 U974 ( .A(G128), .B(n1267), .Z(n1085) );
NOR2_X1 U975 ( .A1(KEYINPUT20), .A2(n1268), .ZN(n1267) );
XOR2_X1 U976 ( .A(G146), .B(G143), .Z(n1268) );
AND2_X1 U977 ( .A1(n1061), .A2(G227), .ZN(n1266) );
XOR2_X1 U978 ( .A(n1269), .B(G101), .Z(n1264) );
NAND2_X1 U979 ( .A1(n1270), .A2(KEYINPUT33), .ZN(n1269) );
XOR2_X1 U980 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U981 ( .A1(KEYINPUT62), .A2(n1253), .ZN(n1272) );
XOR2_X1 U982 ( .A(G104), .B(KEYINPUT17), .Z(n1253) );
XOR2_X1 U983 ( .A(n1024), .B(KEYINPUT39), .Z(n1271) );
XNOR2_X1 U984 ( .A(KEYINPUT56), .B(n1149), .ZN(n1262) );
XOR2_X1 U985 ( .A(n1273), .B(G472), .Z(n1223) );
NAND2_X1 U986 ( .A1(n1274), .A2(n1241), .ZN(n1273) );
XOR2_X1 U987 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR2_X1 U988 ( .A1(KEYINPUT24), .A2(n1148), .ZN(n1276) );
XOR2_X1 U989 ( .A(n1277), .B(G101), .Z(n1148) );
NAND2_X1 U990 ( .A1(n1278), .A2(G210), .ZN(n1277) );
NAND2_X1 U991 ( .A1(n1279), .A2(n1280), .ZN(n1275) );
NAND2_X1 U992 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U993 ( .A1(KEYINPUT50), .A2(n1283), .ZN(n1282) );
OR2_X1 U994 ( .A1(n1154), .A2(KEYINPUT45), .ZN(n1283) );
INV_X1 U995 ( .A(n1284), .ZN(n1281) );
NAND2_X1 U996 ( .A1(n1154), .A2(n1285), .ZN(n1279) );
NAND2_X1 U997 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U998 ( .A1(n1284), .A2(KEYINPUT50), .ZN(n1287) );
XOR2_X1 U999 ( .A(n1149), .B(n1288), .Z(n1284) );
NOR2_X1 U1000 ( .A1(KEYINPUT58), .A2(n1146), .ZN(n1288) );
AND2_X1 U1001 ( .A1(n1289), .A2(n1290), .ZN(n1146) );
NAND2_X1 U1002 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
INV_X1 U1003 ( .A(G146), .ZN(n1292) );
XOR2_X1 U1004 ( .A(n1293), .B(KEYINPUT1), .Z(n1291) );
NAND2_X1 U1005 ( .A1(n1294), .A2(G146), .ZN(n1289) );
XOR2_X1 U1006 ( .A(KEYINPUT34), .B(n1295), .Z(n1294) );
INV_X1 U1007 ( .A(n1293), .ZN(n1295) );
XOR2_X1 U1008 ( .A(n1296), .B(G143), .Z(n1293) );
NAND2_X1 U1009 ( .A1(KEYINPUT57), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1010 ( .A(n1298), .B(G131), .Z(n1149) );
NAND2_X1 U1011 ( .A1(KEYINPUT54), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1012 ( .A(G137), .B(G134), .Z(n1299) );
INV_X1 U1013 ( .A(KEYINPUT45), .ZN(n1286) );
XOR2_X1 U1014 ( .A(n1300), .B(n1254), .Z(n1154) );
XOR2_X1 U1015 ( .A(G116), .B(G119), .Z(n1254) );
INV_X1 U1016 ( .A(n1038), .ZN(n1035) );
NAND2_X1 U1017 ( .A1(n1208), .A2(n1211), .ZN(n1038) );
INV_X1 U1018 ( .A(n1196), .ZN(n1211) );
XOR2_X1 U1019 ( .A(n1301), .B(n1126), .Z(n1196) );
INV_X1 U1020 ( .A(n1075), .ZN(n1126) );
NAND2_X1 U1021 ( .A1(n1241), .A2(n1129), .ZN(n1075) );
NAND3_X1 U1022 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1129) );
OR2_X1 U1023 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND3_X1 U1024 ( .A1(n1306), .A2(n1305), .A3(n1307), .ZN(n1303) );
INV_X1 U1025 ( .A(n1308), .ZN(n1307) );
NAND2_X1 U1026 ( .A1(n1308), .A2(n1309), .ZN(n1302) );
NAND2_X1 U1027 ( .A1(n1310), .A2(n1305), .ZN(n1309) );
INV_X1 U1028 ( .A(KEYINPUT35), .ZN(n1305) );
XNOR2_X1 U1029 ( .A(KEYINPUT55), .B(n1306), .ZN(n1310) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1311), .ZN(n1306) );
XOR2_X1 U1031 ( .A(n1312), .B(n1313), .Z(n1308) );
XOR2_X1 U1032 ( .A(n1024), .B(n1314), .Z(n1313) );
NAND2_X1 U1033 ( .A1(n1315), .A2(KEYINPUT11), .ZN(n1314) );
XOR2_X1 U1034 ( .A(n1297), .B(n1316), .Z(n1315) );
XOR2_X1 U1035 ( .A(G143), .B(G134), .Z(n1316) );
INV_X1 U1036 ( .A(G107), .ZN(n1024) );
XNOR2_X1 U1037 ( .A(G116), .B(n1317), .ZN(n1312) );
XOR2_X1 U1038 ( .A(KEYINPUT19), .B(G122), .Z(n1317) );
NAND2_X1 U1039 ( .A1(KEYINPUT53), .A2(n1130), .ZN(n1301) );
INV_X1 U1040 ( .A(G478), .ZN(n1130) );
INV_X1 U1041 ( .A(n1195), .ZN(n1208) );
NAND2_X1 U1042 ( .A1(n1318), .A2(n1073), .ZN(n1195) );
NAND2_X1 U1043 ( .A1(G475), .A2(n1074), .ZN(n1073) );
OR2_X1 U1044 ( .A1(n1074), .A2(G475), .ZN(n1318) );
NAND2_X1 U1045 ( .A1(n1138), .A2(n1241), .ZN(n1074) );
XNOR2_X1 U1046 ( .A(n1319), .B(n1320), .ZN(n1138) );
XOR2_X1 U1047 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1048 ( .A(KEYINPUT41), .B(G143), .Z(n1322) );
NOR3_X1 U1049 ( .A1(n1323), .A2(KEYINPUT52), .A3(n1324), .ZN(n1321) );
NOR2_X1 U1050 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1051 ( .A(KEYINPUT9), .B(n1327), .Z(n1326) );
NOR2_X1 U1052 ( .A1(n1328), .A2(n1327), .ZN(n1325) );
NOR2_X1 U1053 ( .A1(G104), .A2(n1329), .ZN(n1328) );
NOR2_X1 U1054 ( .A1(n1330), .A2(n1141), .ZN(n1323) );
INV_X1 U1055 ( .A(G104), .ZN(n1141) );
NOR2_X1 U1056 ( .A1(n1327), .A2(n1329), .ZN(n1330) );
INV_X1 U1057 ( .A(KEYINPUT44), .ZN(n1329) );
AND2_X1 U1058 ( .A1(n1331), .A2(n1332), .ZN(n1327) );
NAND2_X1 U1059 ( .A1(n1333), .A2(n1300), .ZN(n1332) );
INV_X1 U1060 ( .A(G113), .ZN(n1300) );
XOR2_X1 U1061 ( .A(n1229), .B(KEYINPUT21), .Z(n1333) );
XOR2_X1 U1062 ( .A(n1334), .B(KEYINPUT5), .Z(n1331) );
NAND2_X1 U1063 ( .A1(G113), .A2(n1229), .ZN(n1334) );
INV_X1 U1064 ( .A(G122), .ZN(n1229) );
XOR2_X1 U1065 ( .A(n1335), .B(n1084), .Z(n1319) );
XNOR2_X1 U1066 ( .A(n1217), .B(G140), .ZN(n1084) );
INV_X1 U1067 ( .A(G131), .ZN(n1217) );
XOR2_X1 U1068 ( .A(n1336), .B(n1337), .Z(n1335) );
NAND2_X1 U1069 ( .A1(n1278), .A2(G214), .ZN(n1336) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1278) );
XNOR2_X1 U1071 ( .A(n1072), .B(KEYINPUT29), .ZN(n1222) );
XOR2_X1 U1072 ( .A(n1338), .B(n1123), .Z(n1072) );
NAND2_X1 U1073 ( .A1(G217), .A2(n1259), .ZN(n1123) );
NAND2_X1 U1074 ( .A1(n1258), .A2(n1241), .ZN(n1259) );
XOR2_X1 U1075 ( .A(G234), .B(KEYINPUT22), .Z(n1258) );
NAND2_X1 U1076 ( .A1(n1121), .A2(n1241), .ZN(n1338) );
INV_X1 U1077 ( .A(G902), .ZN(n1241) );
XNOR2_X1 U1078 ( .A(n1339), .B(n1340), .ZN(n1121) );
XOR2_X1 U1079 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1080 ( .A(n1343), .B(G119), .Z(n1342) );
NAND2_X1 U1081 ( .A1(n1311), .A2(G221), .ZN(n1343) );
AND2_X1 U1082 ( .A1(G234), .A2(n1061), .ZN(n1311) );
INV_X1 U1083 ( .A(G953), .ZN(n1061) );
XOR2_X1 U1084 ( .A(n1297), .B(G137), .Z(n1341) );
INV_X1 U1085 ( .A(G128), .ZN(n1297) );
XNOR2_X1 U1086 ( .A(n1337), .B(n1344), .ZN(n1339) );
XOR2_X1 U1087 ( .A(n1345), .B(n1249), .Z(n1344) );
XOR2_X1 U1088 ( .A(G110), .B(KEYINPUT18), .Z(n1249) );
NOR2_X1 U1089 ( .A1(G140), .A2(KEYINPUT14), .ZN(n1345) );
XOR2_X1 U1090 ( .A(G125), .B(G146), .Z(n1337) );
endmodule


