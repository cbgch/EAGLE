//Key = 1110010110101100000000101001101000001000001110011100011010110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284;

XOR2_X1 U710 ( .A(G107), .B(n977), .Z(G9) );
NOR2_X1 U711 ( .A1(n978), .A2(n979), .ZN(n977) );
NOR2_X1 U712 ( .A1(n980), .A2(n981), .ZN(G75) );
NOR3_X1 U713 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n981) );
NAND3_X1 U714 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n982) );
NAND2_X1 U715 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND2_X1 U716 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND3_X1 U717 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND2_X1 U718 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND3_X1 U719 ( .A1(n997), .A2(n998), .A3(KEYINPUT11), .ZN(n995) );
NAND3_X1 U720 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n992) );
NAND2_X1 U721 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
OR2_X1 U722 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U723 ( .A1(n997), .A2(n1006), .ZN(n999) );
NAND2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
OR2_X1 U725 ( .A1(n1009), .A2(KEYINPUT11), .ZN(n1008) );
NAND2_X1 U726 ( .A1(n1010), .A2(n1011), .ZN(n1007) );
NAND3_X1 U727 ( .A1(n997), .A2(n1012), .A3(n1002), .ZN(n990) );
NAND2_X1 U728 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U729 ( .A1(n1001), .A2(n1015), .ZN(n1014) );
OR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U731 ( .A1(n994), .A2(n1018), .ZN(n1013) );
NAND2_X1 U732 ( .A1(n979), .A2(n1019), .ZN(n1018) );
NAND2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
INV_X1 U734 ( .A(n1022), .ZN(n988) );
NOR3_X1 U735 ( .A1(n1023), .A2(G953), .A3(n1024), .ZN(n980) );
INV_X1 U736 ( .A(n985), .ZN(n1024) );
NAND4_X1 U737 ( .A1(n1010), .A2(n1025), .A3(n997), .A4(n1026), .ZN(n985) );
NOR4_X1 U738 ( .A1(n1021), .A2(n1011), .A3(n1027), .A4(n1028), .ZN(n1026) );
XOR2_X1 U739 ( .A(n1029), .B(n1030), .Z(n1027) );
NOR2_X1 U740 ( .A1(n1031), .A2(KEYINPUT3), .ZN(n1030) );
INV_X1 U741 ( .A(n1032), .ZN(n1031) );
XOR2_X1 U742 ( .A(KEYINPUT14), .B(G952), .Z(n1023) );
XOR2_X1 U743 ( .A(n1033), .B(n1034), .Z(G72) );
NOR2_X1 U744 ( .A1(n1035), .A2(n986), .ZN(n1034) );
NOR2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U746 ( .A(n1038), .B(n1039), .Z(n1033) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XOR2_X1 U748 ( .A(n1042), .B(n1043), .Z(n1041) );
XOR2_X1 U749 ( .A(n1044), .B(n1045), .Z(n1043) );
NAND2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U752 ( .A(KEYINPUT5), .B(n1050), .Z(n1046) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1050) );
XOR2_X1 U754 ( .A(n1051), .B(G134), .Z(n1048) );
NAND2_X1 U755 ( .A1(KEYINPUT49), .A2(G137), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n986), .A2(n1052), .ZN(n1040) );
XOR2_X1 U757 ( .A(KEYINPUT33), .B(G900), .Z(n1052) );
NAND2_X1 U758 ( .A1(KEYINPUT0), .A2(n1053), .ZN(n1038) );
NAND2_X1 U759 ( .A1(n1054), .A2(n986), .ZN(n1053) );
NAND3_X1 U760 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
XOR2_X1 U761 ( .A(n1058), .B(KEYINPUT23), .Z(n1057) );
XOR2_X1 U762 ( .A(n1059), .B(n1060), .Z(G69) );
XOR2_X1 U763 ( .A(n1061), .B(n1062), .Z(n1060) );
NOR4_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
INV_X1 U766 ( .A(KEYINPUT63), .ZN(n1067) );
NOR2_X1 U767 ( .A1(KEYINPUT63), .A2(n1069), .ZN(n1063) );
NOR2_X1 U768 ( .A1(KEYINPUT60), .A2(n1070), .ZN(n1061) );
NOR2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U770 ( .A(KEYINPUT58), .B(G953), .Z(n1072) );
AND2_X1 U771 ( .A1(G224), .A2(G898), .ZN(n1071) );
NAND3_X1 U772 ( .A1(n1073), .A2(n986), .A3(KEYINPUT56), .ZN(n1059) );
NAND2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U774 ( .A(n1076), .ZN(n1075) );
XOR2_X1 U775 ( .A(n1077), .B(KEYINPUT35), .Z(n1074) );
NOR2_X1 U776 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XOR2_X1 U777 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U778 ( .A1(n1032), .A2(n1082), .ZN(n1081) );
NAND2_X1 U779 ( .A1(KEYINPUT13), .A2(n1083), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1078), .A2(n1084), .ZN(G63) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND3_X1 U782 ( .A1(n1087), .A2(n1088), .A3(G478), .ZN(n1085) );
OR2_X1 U783 ( .A1(n1089), .A2(KEYINPUT41), .ZN(n1088) );
NAND2_X1 U784 ( .A1(KEYINPUT41), .A2(n1090), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1091), .A2(n984), .ZN(n1090) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(G60) );
XOR2_X1 U787 ( .A(KEYINPUT4), .B(n1078), .Z(n1093) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1092) );
AND2_X1 U789 ( .A1(G475), .A2(n1089), .ZN(n1095) );
NAND2_X1 U790 ( .A1(KEYINPUT42), .A2(n1096), .ZN(n1094) );
XNOR2_X1 U791 ( .A(G104), .B(n1077), .ZN(G6) );
NOR2_X1 U792 ( .A1(n1078), .A2(n1097), .ZN(G57) );
XOR2_X1 U793 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U794 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U795 ( .A1(n1089), .A2(G472), .ZN(n1100) );
XOR2_X1 U796 ( .A(n1102), .B(KEYINPUT27), .Z(n1098) );
NAND2_X1 U797 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U798 ( .A1(n1078), .A2(n1105), .ZN(G54) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U801 ( .A1(n1089), .A2(G469), .ZN(n1108) );
XNOR2_X1 U802 ( .A(n1110), .B(n1111), .ZN(n1106) );
NOR2_X1 U803 ( .A1(KEYINPUT34), .A2(n1112), .ZN(n1111) );
NAND2_X1 U804 ( .A1(n1113), .A2(KEYINPUT28), .ZN(n1110) );
XOR2_X1 U805 ( .A(n1114), .B(KEYINPUT7), .Z(n1113) );
NOR2_X1 U806 ( .A1(n1078), .A2(n1115), .ZN(G51) );
XOR2_X1 U807 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U808 ( .A(n1118), .B(KEYINPUT53), .ZN(n1117) );
NAND3_X1 U809 ( .A1(n1089), .A2(n1119), .A3(KEYINPUT24), .ZN(n1118) );
XOR2_X1 U810 ( .A(KEYINPUT16), .B(G210), .Z(n1119) );
INV_X1 U811 ( .A(n1082), .ZN(n1089) );
NAND2_X1 U812 ( .A1(G902), .A2(n984), .ZN(n1082) );
NAND4_X1 U813 ( .A1(n1058), .A2(n1077), .A3(n1055), .A4(n1120), .ZN(n984) );
NOR2_X1 U814 ( .A1(n1076), .A2(n1121), .ZN(n1120) );
XNOR2_X1 U815 ( .A(KEYINPUT21), .B(n1056), .ZN(n1121) );
NAND4_X1 U816 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1076) );
AND2_X1 U817 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
NAND2_X1 U818 ( .A1(n1128), .A2(n1129), .ZN(n1122) );
NAND2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND4_X1 U820 ( .A1(n997), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1131) );
NAND3_X1 U821 ( .A1(n1135), .A2(n1136), .A3(n1009), .ZN(n1134) );
INV_X1 U822 ( .A(n998), .ZN(n1009) );
NAND2_X1 U823 ( .A1(n1017), .A2(n1137), .ZN(n1136) );
INV_X1 U824 ( .A(KEYINPUT10), .ZN(n1137) );
OR2_X1 U825 ( .A1(n1138), .A2(KEYINPUT44), .ZN(n1135) );
NAND3_X1 U826 ( .A1(n1139), .A2(n1140), .A3(n998), .ZN(n1133) );
NAND2_X1 U827 ( .A1(KEYINPUT10), .A2(n1017), .ZN(n1140) );
NAND2_X1 U828 ( .A1(KEYINPUT44), .A2(n1016), .ZN(n1139) );
XNOR2_X1 U829 ( .A(KEYINPUT54), .B(n978), .ZN(n1130) );
NAND4_X1 U830 ( .A1(n998), .A2(n1005), .A3(n994), .A4(n1132), .ZN(n978) );
AND4_X1 U831 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1055) );
NOR3_X1 U832 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
OR2_X1 U833 ( .A1(n1148), .A2(n979), .ZN(n1143) );
NAND3_X1 U834 ( .A1(n1004), .A2(n994), .A3(n1149), .ZN(n1077) );
AND2_X1 U835 ( .A1(n1150), .A2(G953), .ZN(n1078) );
XOR2_X1 U836 ( .A(n983), .B(KEYINPUT15), .Z(n1150) );
INV_X1 U837 ( .A(G952), .ZN(n983) );
XOR2_X1 U838 ( .A(G146), .B(n1145), .Z(G48) );
AND3_X1 U839 ( .A1(n1004), .A2(n1128), .A3(n1151), .ZN(n1145) );
XOR2_X1 U840 ( .A(n1152), .B(n1141), .Z(G45) );
NAND3_X1 U841 ( .A1(n1017), .A2(n1153), .A3(n1154), .ZN(n1141) );
NOR3_X1 U842 ( .A1(n979), .A2(n1155), .A3(n1156), .ZN(n1154) );
XNOR2_X1 U843 ( .A(G140), .B(n1056), .ZN(G42) );
NAND2_X1 U844 ( .A1(n1157), .A2(n1016), .ZN(n1056) );
XOR2_X1 U845 ( .A(G137), .B(n1147), .Z(G39) );
AND3_X1 U846 ( .A1(n1001), .A2(n997), .A3(n1151), .ZN(n1147) );
XOR2_X1 U847 ( .A(n1158), .B(n1058), .Z(G36) );
NAND4_X1 U848 ( .A1(n1017), .A2(n1153), .A3(n1001), .A4(n1005), .ZN(n1058) );
XOR2_X1 U849 ( .A(n1049), .B(n1142), .Z(G33) );
NAND2_X1 U850 ( .A1(n1157), .A2(n1017), .ZN(n1142) );
AND3_X1 U851 ( .A1(n1001), .A2(n1004), .A3(n1153), .ZN(n1157) );
INV_X1 U852 ( .A(n996), .ZN(n1001) );
NAND2_X1 U853 ( .A1(n1020), .A2(n1159), .ZN(n996) );
INV_X1 U854 ( .A(n1028), .ZN(n1020) );
XOR2_X1 U855 ( .A(G128), .B(n1146), .Z(G30) );
AND3_X1 U856 ( .A1(n1128), .A2(n1005), .A3(n1151), .ZN(n1146) );
AND3_X1 U857 ( .A1(n1160), .A2(n1161), .A3(n1153), .ZN(n1151) );
AND2_X1 U858 ( .A1(n998), .A2(n1162), .ZN(n1153) );
XOR2_X1 U859 ( .A(n1163), .B(n1164), .Z(G3) );
NAND3_X1 U860 ( .A1(n1017), .A2(n1149), .A3(n1165), .ZN(n1164) );
XNOR2_X1 U861 ( .A(n997), .B(KEYINPUT36), .ZN(n1165) );
XOR2_X1 U862 ( .A(G125), .B(n1166), .Z(G27) );
NOR2_X1 U863 ( .A1(n1167), .A2(n979), .ZN(n1166) );
XOR2_X1 U864 ( .A(n1148), .B(KEYINPUT19), .Z(n1167) );
NAND4_X1 U865 ( .A1(n1016), .A2(n1002), .A3(n1004), .A4(n1162), .ZN(n1148) );
NAND2_X1 U866 ( .A1(n1168), .A2(n1022), .ZN(n1162) );
NAND4_X1 U867 ( .A1(n1169), .A2(G953), .A3(G902), .A4(n1170), .ZN(n1168) );
XOR2_X1 U868 ( .A(n1037), .B(KEYINPUT33), .Z(n1169) );
INV_X1 U869 ( .A(G900), .ZN(n1037) );
XNOR2_X1 U870 ( .A(G122), .B(n1123), .ZN(G24) );
NAND4_X1 U871 ( .A1(n1171), .A2(n994), .A3(n1172), .A4(n1173), .ZN(n1123) );
NOR2_X1 U872 ( .A1(n1174), .A2(n1175), .ZN(n994) );
XNOR2_X1 U873 ( .A(n1125), .B(n1176), .ZN(G21) );
NOR2_X1 U874 ( .A1(KEYINPUT39), .A2(n1177), .ZN(n1176) );
NAND4_X1 U875 ( .A1(n1171), .A2(n997), .A3(n1160), .A4(n1161), .ZN(n1125) );
NAND2_X1 U876 ( .A1(KEYINPUT38), .A2(n1138), .ZN(n1161) );
NAND2_X1 U877 ( .A1(n1178), .A2(n1179), .ZN(n1160) );
INV_X1 U878 ( .A(KEYINPUT38), .ZN(n1179) );
NAND2_X1 U879 ( .A1(n1175), .A2(n1174), .ZN(n1178) );
INV_X1 U880 ( .A(n1025), .ZN(n1174) );
XOR2_X1 U881 ( .A(n1180), .B(n1127), .Z(G18) );
NAND3_X1 U882 ( .A1(n1017), .A2(n1005), .A3(n1171), .ZN(n1127) );
NOR2_X1 U883 ( .A1(n1173), .A2(n1156), .ZN(n1005) );
XOR2_X1 U884 ( .A(n1181), .B(n1126), .Z(G15) );
NAND3_X1 U885 ( .A1(n1017), .A2(n1004), .A3(n1171), .ZN(n1126) );
AND3_X1 U886 ( .A1(n1128), .A2(n1132), .A3(n1002), .ZN(n1171) );
NOR2_X1 U887 ( .A1(n1182), .A2(n1183), .ZN(n1002) );
NOR2_X1 U888 ( .A1(n1172), .A2(n1155), .ZN(n1004) );
NOR2_X1 U889 ( .A1(n1175), .A2(n1025), .ZN(n1017) );
XNOR2_X1 U890 ( .A(G110), .B(n1184), .ZN(G12) );
NAND3_X1 U891 ( .A1(n1149), .A2(n997), .A3(n1016), .ZN(n1184) );
INV_X1 U892 ( .A(n1138), .ZN(n1016) );
NAND2_X1 U893 ( .A1(n1025), .A2(n1175), .ZN(n1138) );
XOR2_X1 U894 ( .A(n1185), .B(n1032), .Z(n1175) );
NAND2_X1 U895 ( .A1(G217), .A2(n1186), .ZN(n1032) );
XOR2_X1 U896 ( .A(n1029), .B(KEYINPUT31), .Z(n1185) );
NAND2_X1 U897 ( .A1(n1083), .A2(n1091), .ZN(n1029) );
XNOR2_X1 U898 ( .A(n1187), .B(n1188), .ZN(n1083) );
XOR2_X1 U899 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U900 ( .A(n1177), .B(G137), .Z(n1190) );
INV_X1 U901 ( .A(G119), .ZN(n1177) );
NAND2_X1 U902 ( .A1(KEYINPUT30), .A2(n1191), .ZN(n1189) );
XOR2_X1 U903 ( .A(n1042), .B(n1192), .Z(n1191) );
XOR2_X1 U904 ( .A(KEYINPUT26), .B(G146), .Z(n1192) );
XNOR2_X1 U905 ( .A(n1193), .B(n1194), .ZN(n1187) );
XOR2_X1 U906 ( .A(n1195), .B(n1196), .Z(n1194) );
AND3_X1 U907 ( .A1(G221), .A2(n986), .A3(G234), .ZN(n1196) );
NOR2_X1 U908 ( .A1(G128), .A2(KEYINPUT18), .ZN(n1195) );
XOR2_X1 U909 ( .A(n1197), .B(G472), .Z(n1025) );
NAND2_X1 U910 ( .A1(n1198), .A2(n1091), .ZN(n1197) );
XOR2_X1 U911 ( .A(n1101), .B(n1199), .Z(n1198) );
XOR2_X1 U912 ( .A(KEYINPUT20), .B(n1200), .Z(n1199) );
NOR2_X1 U913 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U914 ( .A(KEYINPUT61), .B(n1103), .ZN(n1202) );
NAND2_X1 U915 ( .A1(n1163), .A2(n1203), .ZN(n1103) );
NAND2_X1 U916 ( .A1(n1204), .A2(G210), .ZN(n1203) );
INV_X1 U917 ( .A(G101), .ZN(n1163) );
INV_X1 U918 ( .A(n1104), .ZN(n1201) );
NAND3_X1 U919 ( .A1(G101), .A2(G210), .A3(n1204), .ZN(n1104) );
XOR2_X1 U920 ( .A(n1205), .B(n1206), .Z(n1101) );
XOR2_X1 U921 ( .A(G113), .B(n1207), .Z(n1206) );
NOR2_X1 U922 ( .A1(KEYINPUT50), .A2(n1208), .ZN(n1207) );
XOR2_X1 U923 ( .A(n1112), .B(n1209), .Z(n1205) );
NOR2_X1 U924 ( .A1(n1172), .A2(n1173), .ZN(n997) );
INV_X1 U925 ( .A(n1155), .ZN(n1173) );
XNOR2_X1 U926 ( .A(G475), .B(n1210), .ZN(n1155) );
NOR2_X1 U927 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U928 ( .A(KEYINPUT32), .B(G902), .Z(n1212) );
INV_X1 U929 ( .A(n1096), .ZN(n1211) );
NAND2_X1 U930 ( .A1(n1213), .A2(n1214), .ZN(n1096) );
NAND2_X1 U931 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U932 ( .A(KEYINPUT43), .B(n1217), .Z(n1213) );
NOR2_X1 U933 ( .A1(n1216), .A2(n1215), .ZN(n1217) );
XOR2_X1 U934 ( .A(n1218), .B(n1219), .Z(n1215) );
XNOR2_X1 U935 ( .A(n1220), .B(n1221), .ZN(n1219) );
XOR2_X1 U936 ( .A(n1049), .B(n1222), .Z(n1221) );
NAND2_X1 U937 ( .A1(n1204), .A2(G214), .ZN(n1222) );
NOR2_X1 U938 ( .A1(G953), .A2(G237), .ZN(n1204) );
NAND2_X1 U939 ( .A1(KEYINPUT2), .A2(G143), .ZN(n1220) );
XOR2_X1 U940 ( .A(n1223), .B(n1042), .Z(n1218) );
XOR2_X1 U941 ( .A(G125), .B(G140), .Z(n1042) );
NAND2_X1 U942 ( .A1(KEYINPUT1), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U943 ( .A(G104), .B(n1225), .ZN(n1216) );
XOR2_X1 U944 ( .A(G122), .B(G113), .Z(n1225) );
INV_X1 U945 ( .A(n1156), .ZN(n1172) );
XOR2_X1 U946 ( .A(n1226), .B(G478), .Z(n1156) );
NAND2_X1 U947 ( .A1(n1086), .A2(n1091), .ZN(n1226) );
XNOR2_X1 U948 ( .A(n1227), .B(n1228), .ZN(n1086) );
XNOR2_X1 U949 ( .A(n1229), .B(n1230), .ZN(n1228) );
AND4_X1 U950 ( .A1(n1231), .A2(n986), .A3(G234), .A4(G217), .ZN(n1230) );
INV_X1 U951 ( .A(KEYINPUT37), .ZN(n1231) );
NAND2_X1 U952 ( .A1(KEYINPUT47), .A2(G107), .ZN(n1229) );
NAND2_X1 U953 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
NAND2_X1 U954 ( .A1(n1234), .A2(n1180), .ZN(n1233) );
XOR2_X1 U955 ( .A(KEYINPUT6), .B(n1235), .Z(n1234) );
NAND2_X1 U956 ( .A1(n1236), .A2(G116), .ZN(n1232) );
XOR2_X1 U957 ( .A(KEYINPUT8), .B(n1235), .Z(n1236) );
XNOR2_X1 U958 ( .A(n1237), .B(G122), .ZN(n1235) );
NAND3_X1 U959 ( .A1(n1238), .A2(n1239), .A3(KEYINPUT59), .ZN(n1237) );
NAND2_X1 U960 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND2_X1 U961 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U962 ( .A(G134), .B(n1244), .Z(n1240) );
NOR2_X1 U963 ( .A1(G143), .A2(KEYINPUT52), .ZN(n1244) );
NAND3_X1 U964 ( .A1(n1242), .A2(n1243), .A3(n1245), .ZN(n1238) );
XOR2_X1 U965 ( .A(n1158), .B(n1246), .Z(n1245) );
OR2_X1 U966 ( .A1(n1152), .A2(KEYINPUT52), .ZN(n1246) );
INV_X1 U967 ( .A(G143), .ZN(n1152) );
INV_X1 U968 ( .A(G134), .ZN(n1158) );
INV_X1 U969 ( .A(KEYINPUT55), .ZN(n1243) );
AND3_X1 U970 ( .A1(n998), .A2(n1132), .A3(n1128), .ZN(n1149) );
INV_X1 U971 ( .A(n979), .ZN(n1128) );
NAND2_X1 U972 ( .A1(n1247), .A2(n1159), .ZN(n979) );
XOR2_X1 U973 ( .A(n1021), .B(KEYINPUT12), .Z(n1159) );
AND2_X1 U974 ( .A1(n1248), .A2(G214), .ZN(n1021) );
XOR2_X1 U975 ( .A(n1249), .B(KEYINPUT40), .Z(n1248) );
OR2_X1 U976 ( .A1(G902), .A2(G237), .ZN(n1249) );
XOR2_X1 U977 ( .A(n1028), .B(KEYINPUT57), .Z(n1247) );
NAND3_X1 U978 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1028) );
OR2_X1 U979 ( .A1(n1253), .A2(n1116), .ZN(n1252) );
NAND3_X1 U980 ( .A1(n1116), .A2(n1253), .A3(n1091), .ZN(n1251) );
NAND2_X1 U981 ( .A1(G237), .A2(G210), .ZN(n1253) );
XNOR2_X1 U982 ( .A(n1254), .B(n1255), .ZN(n1116) );
XOR2_X1 U983 ( .A(G125), .B(n1256), .Z(n1255) );
AND2_X1 U984 ( .A1(n986), .A2(G224), .ZN(n1256) );
XOR2_X1 U985 ( .A(n1257), .B(n1209), .Z(n1254) );
XNOR2_X1 U986 ( .A(n1258), .B(n1259), .ZN(n1209) );
XOR2_X1 U987 ( .A(G143), .B(G128), .Z(n1259) );
XOR2_X1 U988 ( .A(n1224), .B(KEYINPUT62), .Z(n1258) );
INV_X1 U989 ( .A(G146), .ZN(n1224) );
NAND2_X1 U990 ( .A1(n1260), .A2(n1068), .ZN(n1257) );
NAND2_X1 U991 ( .A1(n1261), .A2(n1069), .ZN(n1068) );
INV_X1 U992 ( .A(n1065), .ZN(n1260) );
NOR2_X1 U993 ( .A1(n1069), .A2(n1261), .ZN(n1065) );
XOR2_X1 U994 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U995 ( .A(n1264), .B(n1208), .ZN(n1263) );
XOR2_X1 U996 ( .A(G119), .B(n1180), .Z(n1208) );
INV_X1 U997 ( .A(G116), .ZN(n1180) );
NOR2_X1 U998 ( .A1(KEYINPUT25), .A2(n1181), .ZN(n1264) );
INV_X1 U999 ( .A(G113), .ZN(n1181) );
XNOR2_X1 U1000 ( .A(G122), .B(n1193), .ZN(n1069) );
NAND2_X1 U1001 ( .A1(G902), .A2(G210), .ZN(n1250) );
NAND2_X1 U1002 ( .A1(n1022), .A2(n1265), .ZN(n1132) );
NAND3_X1 U1003 ( .A1(G902), .A2(n1170), .A3(n1066), .ZN(n1265) );
NOR2_X1 U1004 ( .A1(n986), .A2(G898), .ZN(n1066) );
NAND3_X1 U1005 ( .A1(n1170), .A2(n986), .A3(G952), .ZN(n1022) );
INV_X1 U1006 ( .A(G953), .ZN(n986) );
NAND2_X1 U1007 ( .A1(G234), .A2(G237), .ZN(n1170) );
NOR2_X1 U1008 ( .A1(n1183), .A2(n1010), .ZN(n998) );
INV_X1 U1009 ( .A(n1182), .ZN(n1010) );
XNOR2_X1 U1010 ( .A(n1266), .B(G469), .ZN(n1182) );
NAND2_X1 U1011 ( .A1(n1267), .A2(n1091), .ZN(n1266) );
XOR2_X1 U1012 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U1013 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
AND3_X1 U1014 ( .A1(KEYINPUT9), .A2(n1044), .A3(n1262), .ZN(n1271) );
NOR2_X1 U1015 ( .A1(KEYINPUT9), .A2(n1109), .ZN(n1270) );
XNOR2_X1 U1016 ( .A(n1044), .B(n1262), .ZN(n1109) );
XNOR2_X1 U1017 ( .A(G101), .B(n1272), .ZN(n1262) );
XOR2_X1 U1018 ( .A(G107), .B(G104), .Z(n1272) );
NAND2_X1 U1019 ( .A1(n1273), .A2(n1274), .ZN(n1044) );
NAND2_X1 U1020 ( .A1(n1275), .A2(n1242), .ZN(n1274) );
XOR2_X1 U1021 ( .A(KEYINPUT22), .B(n1276), .Z(n1273) );
NOR2_X1 U1022 ( .A1(n1242), .A2(n1275), .ZN(n1276) );
XOR2_X1 U1023 ( .A(G143), .B(n1277), .Z(n1275) );
NOR2_X1 U1024 ( .A1(G146), .A2(KEYINPUT46), .ZN(n1277) );
INV_X1 U1025 ( .A(G128), .ZN(n1242) );
XNOR2_X1 U1026 ( .A(n1278), .B(n1279), .ZN(n1268) );
NOR2_X1 U1027 ( .A1(KEYINPUT45), .A2(n1112), .ZN(n1279) );
XOR2_X1 U1028 ( .A(n1049), .B(n1280), .Z(n1112) );
XOR2_X1 U1029 ( .A(G137), .B(G134), .Z(n1280) );
INV_X1 U1030 ( .A(G131), .ZN(n1049) );
NOR2_X1 U1031 ( .A1(KEYINPUT17), .A2(n1281), .ZN(n1278) );
XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n1282), .Z(n1281) );
INV_X1 U1033 ( .A(n1114), .ZN(n1282) );
XNOR2_X1 U1034 ( .A(n1193), .B(n1283), .ZN(n1114) );
XOR2_X1 U1035 ( .A(G140), .B(n1284), .Z(n1283) );
NOR2_X1 U1036 ( .A1(G953), .A2(n1036), .ZN(n1284) );
INV_X1 U1037 ( .A(G227), .ZN(n1036) );
XOR2_X1 U1038 ( .A(G110), .B(KEYINPUT48), .Z(n1193) );
XOR2_X1 U1039 ( .A(n1011), .B(KEYINPUT29), .Z(n1183) );
AND2_X1 U1040 ( .A1(G221), .A2(n1186), .ZN(n1011) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1091), .ZN(n1186) );
INV_X1 U1042 ( .A(G902), .ZN(n1091) );
endmodule


