//Key = 1001100110111000011110000101000011000010100111100101010011011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277;

XOR2_X1 U726 ( .A(n984), .B(n985), .Z(G9) );
NAND2_X1 U727 ( .A1(KEYINPUT43), .A2(n986), .ZN(n985) );
XOR2_X1 U728 ( .A(KEYINPUT14), .B(G107), .Z(n986) );
NOR2_X1 U729 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U730 ( .A1(G953), .A2(n989), .A3(n990), .A4(n991), .ZN(n988) );
NOR2_X1 U731 ( .A1(n992), .A2(n993), .ZN(n990) );
NOR2_X1 U732 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR3_X1 U733 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NOR2_X1 U734 ( .A1(n999), .A2(n1000), .ZN(n997) );
AND2_X1 U735 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NOR2_X1 U736 ( .A1(n1003), .A2(n1004), .ZN(n999) );
NOR2_X1 U737 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U738 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U739 ( .A1(n1009), .A2(n1010), .ZN(n1005) );
NOR2_X1 U740 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR4_X1 U741 ( .A1(n1013), .A2(n1010), .A3(n1008), .A4(n1004), .ZN(n994) );
INV_X1 U742 ( .A(n1002), .ZN(n1008) );
NOR3_X1 U743 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U744 ( .A1(n1017), .A2(n998), .ZN(n1016) );
NOR2_X1 U745 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR3_X1 U746 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1015) );
XOR2_X1 U747 ( .A(KEYINPUT17), .B(n1023), .Z(n1020) );
NOR2_X1 U748 ( .A1(n1024), .A2(n996), .ZN(n1014) );
NOR3_X1 U749 ( .A1(n989), .A2(G953), .A3(G952), .ZN(n987) );
AND4_X1 U750 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n989) );
NOR4_X1 U751 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1004), .ZN(n1028) );
INV_X1 U752 ( .A(n1032), .ZN(n1004) );
XOR2_X1 U753 ( .A(n1033), .B(KEYINPUT32), .Z(n1029) );
NOR3_X1 U754 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1027) );
INV_X1 U755 ( .A(n1007), .ZN(n1036) );
NOR2_X1 U756 ( .A1(n1037), .A2(n1038), .ZN(n1034) );
XOR2_X1 U757 ( .A(KEYINPUT20), .B(n1039), .Z(n1026) );
XOR2_X1 U758 ( .A(KEYINPUT59), .B(n1040), .Z(n1025) );
AND2_X1 U759 ( .A1(n1038), .A2(n1037), .ZN(n1040) );
XOR2_X1 U760 ( .A(n1041), .B(n1042), .Z(G72) );
XOR2_X1 U761 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U762 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XOR2_X1 U763 ( .A(n1047), .B(n1048), .Z(n1046) );
NAND2_X1 U764 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U765 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U766 ( .A(KEYINPUT51), .B(n1053), .Z(n1049) );
NOR2_X1 U767 ( .A1(n1051), .A2(n1052), .ZN(n1053) );
XOR2_X1 U768 ( .A(n1054), .B(n1055), .Z(n1051) );
NOR2_X1 U769 ( .A1(KEYINPUT24), .A2(n1056), .ZN(n1055) );
NAND2_X1 U770 ( .A1(n1057), .A2(n1058), .ZN(n1043) );
NAND2_X1 U771 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U772 ( .A1(G953), .A2(n1061), .A3(KEYINPUT19), .ZN(n1041) );
NAND2_X1 U773 ( .A1(G900), .A2(G227), .ZN(n1061) );
NAND2_X1 U774 ( .A1(n1062), .A2(n1063), .ZN(G69) );
NAND2_X1 U775 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U776 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NAND2_X1 U777 ( .A1(KEYINPUT62), .A2(n1068), .ZN(n1067) );
OR3_X1 U778 ( .A1(n1069), .A2(KEYINPUT62), .A3(n1065), .ZN(n1062) );
NAND2_X1 U779 ( .A1(G953), .A2(n1070), .ZN(n1065) );
NAND2_X1 U780 ( .A1(G224), .A2(G898), .ZN(n1070) );
XOR2_X1 U781 ( .A(n1068), .B(n1066), .Z(n1069) );
AND2_X1 U782 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
NAND3_X1 U783 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NAND2_X1 U784 ( .A1(n1076), .A2(G953), .ZN(n1074) );
XOR2_X1 U785 ( .A(KEYINPUT56), .B(n1077), .Z(n1071) );
NOR3_X1 U786 ( .A1(n1073), .A2(G953), .A3(n1075), .ZN(n1077) );
XNOR2_X1 U787 ( .A(n1078), .B(n1079), .ZN(n1073) );
NAND2_X1 U788 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND2_X1 U789 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U790 ( .A(n1084), .B(KEYINPUT5), .Z(n1082) );
INV_X1 U791 ( .A(n1085), .ZN(n1080) );
INV_X1 U792 ( .A(KEYINPUT52), .ZN(n1068) );
NOR2_X1 U793 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XNOR2_X1 U794 ( .A(n1088), .B(n1089), .ZN(n1087) );
NOR2_X1 U795 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U796 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XOR2_X1 U797 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U798 ( .A1(n1095), .A2(n1091), .ZN(n1093) );
INV_X1 U799 ( .A(G478), .ZN(n1095) );
NOR2_X1 U800 ( .A1(n1086), .A2(n1096), .ZN(G60) );
XNOR2_X1 U801 ( .A(n1097), .B(n1098), .ZN(n1096) );
NOR2_X1 U802 ( .A1(n1099), .A2(n1091), .ZN(n1098) );
INV_X1 U803 ( .A(G475), .ZN(n1099) );
NAND2_X1 U804 ( .A1(n1100), .A2(n1101), .ZN(G6) );
NAND2_X1 U805 ( .A1(G104), .A2(n1102), .ZN(n1101) );
XOR2_X1 U806 ( .A(KEYINPUT27), .B(n1103), .Z(n1100) );
NOR2_X1 U807 ( .A1(G104), .A2(n1102), .ZN(n1103) );
NOR2_X1 U808 ( .A1(n1086), .A2(n1104), .ZN(G57) );
XOR2_X1 U809 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U810 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U811 ( .A1(KEYINPUT38), .A2(n1109), .ZN(n1107) );
XOR2_X1 U812 ( .A(n1110), .B(n1111), .Z(n1105) );
NOR2_X1 U813 ( .A1(n1112), .A2(n1091), .ZN(n1111) );
INV_X1 U814 ( .A(G472), .ZN(n1112) );
NAND2_X1 U815 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XOR2_X1 U816 ( .A(n1115), .B(KEYINPUT58), .Z(n1113) );
NOR2_X1 U817 ( .A1(n1086), .A2(n1116), .ZN(G54) );
XOR2_X1 U818 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U819 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND3_X1 U820 ( .A1(G902), .A2(G469), .A3(n1121), .ZN(n1119) );
XOR2_X1 U821 ( .A(n991), .B(KEYINPUT16), .Z(n1121) );
XOR2_X1 U822 ( .A(n1122), .B(KEYINPUT39), .Z(n1117) );
NAND2_X1 U823 ( .A1(n1123), .A2(KEYINPUT49), .ZN(n1122) );
XOR2_X1 U824 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U825 ( .A(G140), .B(G110), .Z(n1125) );
NAND2_X1 U826 ( .A1(n1126), .A2(KEYINPUT44), .ZN(n1124) );
XOR2_X1 U827 ( .A(n1127), .B(KEYINPUT33), .Z(n1126) );
NOR2_X1 U828 ( .A1(n1086), .A2(n1128), .ZN(G51) );
XOR2_X1 U829 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U830 ( .A1(n1038), .A2(n1091), .ZN(n1130) );
NAND2_X1 U831 ( .A1(G902), .A2(n991), .ZN(n1091) );
NAND3_X1 U832 ( .A1(n1075), .A2(n1059), .A3(n1131), .ZN(n991) );
XOR2_X1 U833 ( .A(n1060), .B(KEYINPUT37), .Z(n1131) );
AND4_X1 U834 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1059) );
NOR4_X1 U835 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
NOR3_X1 U836 ( .A1(n1140), .A2(n1141), .A3(n996), .ZN(n1139) );
XOR2_X1 U837 ( .A(n998), .B(KEYINPUT21), .Z(n1141) );
INV_X1 U838 ( .A(n1142), .ZN(n998) );
INV_X1 U839 ( .A(n1143), .ZN(n1138) );
NAND2_X1 U840 ( .A1(n1144), .A2(n1018), .ZN(n1134) );
AND4_X1 U841 ( .A1(n1102), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1075) );
AND4_X1 U842 ( .A1(n984), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1147) );
NAND3_X1 U843 ( .A1(n1002), .A2(n1019), .A3(n1151), .ZN(n984) );
NAND2_X1 U844 ( .A1(n1152), .A2(n1153), .ZN(n1146) );
NAND2_X1 U845 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND3_X1 U846 ( .A1(n1151), .A2(n1002), .A3(n1018), .ZN(n1102) );
NOR2_X1 U847 ( .A1(n1156), .A2(n1157), .ZN(n1129) );
XOR2_X1 U848 ( .A(KEYINPUT41), .B(n1158), .Z(n1157) );
NOR2_X1 U849 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND2_X1 U850 ( .A1(n1160), .A2(n1159), .ZN(n1156) );
XNOR2_X1 U851 ( .A(n1161), .B(n1162), .ZN(n1160) );
NAND2_X1 U852 ( .A1(KEYINPUT12), .A2(n1163), .ZN(n1161) );
XOR2_X1 U853 ( .A(n1164), .B(n1052), .Z(n1163) );
NOR2_X1 U854 ( .A1(G125), .A2(KEYINPUT31), .ZN(n1164) );
NOR2_X1 U855 ( .A1(n1057), .A2(G952), .ZN(n1086) );
XOR2_X1 U856 ( .A(n1165), .B(n1060), .Z(G48) );
NAND3_X1 U857 ( .A1(n1018), .A2(n1152), .A3(n1166), .ZN(n1060) );
XOR2_X1 U858 ( .A(n1167), .B(n1143), .Z(G45) );
NAND4_X1 U859 ( .A1(n1012), .A2(n1168), .A3(n1001), .A4(n1169), .ZN(n1143) );
XOR2_X1 U860 ( .A(G140), .B(n1137), .Z(G42) );
AND3_X1 U861 ( .A1(n1018), .A2(n1011), .A3(n1170), .ZN(n1137) );
XOR2_X1 U862 ( .A(n1171), .B(G137), .Z(G39) );
NAND2_X1 U863 ( .A1(KEYINPUT18), .A2(n1172), .ZN(n1171) );
NAND3_X1 U864 ( .A1(n1023), .A2(n1142), .A3(n1166), .ZN(n1172) );
XOR2_X1 U865 ( .A(n1173), .B(G134), .Z(G36) );
NAND2_X1 U866 ( .A1(KEYINPUT60), .A2(n1132), .ZN(n1173) );
NAND2_X1 U867 ( .A1(n1144), .A2(n1019), .ZN(n1132) );
XOR2_X1 U868 ( .A(n1174), .B(n1175), .Z(G33) );
NAND2_X1 U869 ( .A1(n1144), .A2(n1176), .ZN(n1175) );
XOR2_X1 U870 ( .A(KEYINPUT26), .B(n1018), .Z(n1176) );
AND2_X1 U871 ( .A1(n1170), .A2(n1012), .ZN(n1144) );
AND3_X1 U872 ( .A1(n1142), .A2(n1169), .A3(n1001), .ZN(n1170) );
XOR2_X1 U873 ( .A(G128), .B(n1136), .Z(G30) );
AND3_X1 U874 ( .A1(n1019), .A2(n1152), .A3(n1166), .ZN(n1136) );
INV_X1 U875 ( .A(n1140), .ZN(n1166) );
NAND4_X1 U876 ( .A1(n1001), .A2(n1030), .A3(n1177), .A4(n1169), .ZN(n1140) );
XOR2_X1 U877 ( .A(n1178), .B(n1145), .Z(G3) );
NAND3_X1 U878 ( .A1(n1151), .A2(n1023), .A3(n1012), .ZN(n1145) );
XNOR2_X1 U879 ( .A(G125), .B(n1133), .ZN(G27) );
NAND4_X1 U880 ( .A1(n1152), .A2(n1169), .A3(n1179), .A4(n1180), .ZN(n1133) );
AND3_X1 U881 ( .A1(n1018), .A2(n1011), .A3(n1032), .ZN(n1180) );
NAND2_X1 U882 ( .A1(n993), .A2(n1181), .ZN(n1169) );
NAND3_X1 U883 ( .A1(G902), .A2(n1182), .A3(n1045), .ZN(n1181) );
NOR2_X1 U884 ( .A1(n1057), .A2(G900), .ZN(n1045) );
XNOR2_X1 U885 ( .A(G122), .B(n1150), .ZN(G24) );
NAND3_X1 U886 ( .A1(n1183), .A2(n1002), .A3(n1168), .ZN(n1150) );
AND3_X1 U887 ( .A1(n1031), .A2(n1152), .A3(n1184), .ZN(n1168) );
NOR2_X1 U888 ( .A1(n1177), .A2(n1185), .ZN(n1002) );
XOR2_X1 U889 ( .A(KEYINPUT11), .B(n1186), .Z(n1185) );
XNOR2_X1 U890 ( .A(G119), .B(n1149), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1177), .A2(n1152), .A3(n1030), .A4(n1187), .ZN(n1149) );
NOR2_X1 U892 ( .A1(n996), .A2(n1188), .ZN(n1187) );
INV_X1 U893 ( .A(n1023), .ZN(n996) );
XOR2_X1 U894 ( .A(G116), .B(n1189), .Z(G18) );
NOR3_X1 U895 ( .A1(n1190), .A2(KEYINPUT35), .A3(n1024), .ZN(n1189) );
XNOR2_X1 U896 ( .A(KEYINPUT57), .B(n1154), .ZN(n1190) );
NAND3_X1 U897 ( .A1(n1183), .A2(n1019), .A3(n1012), .ZN(n1154) );
NAND2_X1 U898 ( .A1(n1191), .A2(n1192), .ZN(n1019) );
OR3_X1 U899 ( .A1(n1033), .A2(n1031), .A3(KEYINPUT28), .ZN(n1192) );
NAND2_X1 U900 ( .A1(KEYINPUT28), .A2(n1023), .ZN(n1191) );
XOR2_X1 U901 ( .A(G113), .B(n1193), .Z(G15) );
NOR2_X1 U902 ( .A1(n1024), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U903 ( .A(KEYINPUT4), .B(n1155), .ZN(n1194) );
NAND3_X1 U904 ( .A1(n1012), .A2(n1183), .A3(n1018), .ZN(n1155) );
AND2_X1 U905 ( .A1(n1033), .A2(n1031), .ZN(n1018) );
INV_X1 U906 ( .A(n1188), .ZN(n1183) );
NAND3_X1 U907 ( .A1(n1179), .A2(n1195), .A3(n1032), .ZN(n1188) );
AND2_X1 U908 ( .A1(n1196), .A2(n1177), .ZN(n1012) );
XOR2_X1 U909 ( .A(KEYINPUT11), .B(n1030), .Z(n1196) );
INV_X1 U910 ( .A(n1186), .ZN(n1030) );
INV_X1 U911 ( .A(n1152), .ZN(n1024) );
XOR2_X1 U912 ( .A(G110), .B(n1197), .Z(G12) );
NOR2_X1 U913 ( .A1(KEYINPUT23), .A2(n1148), .ZN(n1197) );
NAND3_X1 U914 ( .A1(n1151), .A2(n1023), .A3(n1011), .ZN(n1148) );
NOR2_X1 U915 ( .A1(n1177), .A2(n1186), .ZN(n1011) );
XNOR2_X1 U916 ( .A(n1198), .B(n1090), .ZN(n1186) );
NAND2_X1 U917 ( .A1(G217), .A2(n1199), .ZN(n1090) );
NAND2_X1 U918 ( .A1(n1088), .A2(n1200), .ZN(n1198) );
XNOR2_X1 U919 ( .A(n1201), .B(n1202), .ZN(n1088) );
XOR2_X1 U920 ( .A(n1048), .B(n1203), .Z(n1202) );
XOR2_X1 U921 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U922 ( .A1(KEYINPUT48), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U923 ( .A(G119), .B(n1207), .ZN(n1206) );
NAND2_X1 U924 ( .A1(n1208), .A2(G221), .ZN(n1204) );
XOR2_X1 U925 ( .A(n1209), .B(n1210), .Z(n1201) );
XOR2_X1 U926 ( .A(KEYINPUT0), .B(G146), .Z(n1210) );
XOR2_X1 U927 ( .A(G137), .B(n1211), .Z(n1209) );
XOR2_X1 U928 ( .A(n1039), .B(KEYINPUT63), .Z(n1177) );
XNOR2_X1 U929 ( .A(n1212), .B(G472), .ZN(n1039) );
NAND2_X1 U930 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U931 ( .A(n1109), .B(n1215), .Z(n1214) );
XOR2_X1 U932 ( .A(n1216), .B(n1108), .Z(n1215) );
XOR2_X1 U933 ( .A(n1217), .B(n1218), .Z(n1108) );
INV_X1 U934 ( .A(n1219), .ZN(n1218) );
NAND2_X1 U935 ( .A1(KEYINPUT45), .A2(n1220), .ZN(n1217) );
NAND2_X1 U936 ( .A1(n1115), .A2(n1114), .ZN(n1216) );
NAND4_X1 U937 ( .A1(n1221), .A2(G210), .A3(G101), .A4(n1222), .ZN(n1114) );
NAND2_X1 U938 ( .A1(n1178), .A2(n1223), .ZN(n1115) );
NAND3_X1 U939 ( .A1(n1221), .A2(n1222), .A3(G210), .ZN(n1223) );
XOR2_X1 U940 ( .A(KEYINPUT10), .B(G902), .Z(n1213) );
NOR2_X1 U941 ( .A1(n1031), .A2(n1184), .ZN(n1023) );
INV_X1 U942 ( .A(n1033), .ZN(n1184) );
XOR2_X1 U943 ( .A(n1224), .B(G478), .Z(n1033) );
OR2_X1 U944 ( .A1(n1094), .A2(G902), .ZN(n1224) );
XNOR2_X1 U945 ( .A(n1225), .B(n1226), .ZN(n1094) );
XOR2_X1 U946 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND2_X1 U947 ( .A1(n1208), .A2(G217), .ZN(n1228) );
AND2_X1 U948 ( .A1(n1221), .A2(G234), .ZN(n1208) );
NAND2_X1 U949 ( .A1(KEYINPUT7), .A2(n1229), .ZN(n1227) );
XOR2_X1 U950 ( .A(G122), .B(G116), .Z(n1229) );
XOR2_X1 U951 ( .A(n1230), .B(n1231), .Z(n1225) );
NOR2_X1 U952 ( .A1(KEYINPUT61), .A2(n1232), .ZN(n1231) );
XOR2_X1 U953 ( .A(G143), .B(n1233), .Z(n1232) );
NOR2_X1 U954 ( .A1(KEYINPUT1), .A2(n1207), .ZN(n1233) );
XNOR2_X1 U955 ( .A(G107), .B(G134), .ZN(n1230) );
XNOR2_X1 U956 ( .A(n1234), .B(G475), .ZN(n1031) );
NAND2_X1 U957 ( .A1(n1097), .A2(n1200), .ZN(n1234) );
XNOR2_X1 U958 ( .A(n1235), .B(n1236), .ZN(n1097) );
XOR2_X1 U959 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U960 ( .A(n1219), .B(n1239), .Z(n1238) );
AND3_X1 U961 ( .A1(G214), .A2(n1222), .A3(n1221), .ZN(n1239) );
NAND2_X1 U962 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
NAND2_X1 U963 ( .A1(n1242), .A2(n1165), .ZN(n1241) );
INV_X1 U964 ( .A(G146), .ZN(n1165) );
XOR2_X1 U965 ( .A(n1243), .B(KEYINPUT42), .Z(n1242) );
NAND2_X1 U966 ( .A1(n1244), .A2(G146), .ZN(n1240) );
XOR2_X1 U967 ( .A(KEYINPUT15), .B(n1245), .Z(n1244) );
INV_X1 U968 ( .A(n1243), .ZN(n1245) );
XOR2_X1 U969 ( .A(n1048), .B(KEYINPUT8), .Z(n1243) );
XNOR2_X1 U970 ( .A(G125), .B(G140), .ZN(n1048) );
XOR2_X1 U971 ( .A(n1246), .B(n1247), .Z(n1235) );
XNOR2_X1 U972 ( .A(n1248), .B(n1249), .ZN(n1247) );
NOR2_X1 U973 ( .A1(KEYINPUT6), .A2(n1174), .ZN(n1249) );
NAND2_X1 U974 ( .A1(KEYINPUT46), .A2(G104), .ZN(n1248) );
XOR2_X1 U975 ( .A(G122), .B(n1167), .Z(n1246) );
AND3_X1 U976 ( .A1(n1152), .A2(n1195), .A3(n1001), .ZN(n1151) );
NOR2_X1 U977 ( .A1(n1010), .A2(n1032), .ZN(n1001) );
XOR2_X1 U978 ( .A(n1250), .B(G469), .Z(n1032) );
NAND2_X1 U979 ( .A1(n1251), .A2(n1200), .ZN(n1250) );
XOR2_X1 U980 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U981 ( .A(n1254), .B(n1127), .ZN(n1253) );
NAND2_X1 U982 ( .A1(G227), .A2(n1221), .ZN(n1127) );
NOR2_X1 U983 ( .A1(KEYINPUT54), .A2(n1255), .ZN(n1254) );
XOR2_X1 U984 ( .A(n1256), .B(G140), .Z(n1255) );
NAND2_X1 U985 ( .A1(KEYINPUT3), .A2(n1211), .ZN(n1256) );
INV_X1 U986 ( .A(n1120), .ZN(n1252) );
XOR2_X1 U987 ( .A(n1257), .B(n1109), .Z(n1120) );
XNOR2_X1 U988 ( .A(n1258), .B(n1259), .ZN(n1109) );
XNOR2_X1 U989 ( .A(n1052), .B(n1056), .ZN(n1259) );
XNOR2_X1 U990 ( .A(G134), .B(G137), .ZN(n1056) );
XOR2_X1 U991 ( .A(n1054), .B(KEYINPUT13), .Z(n1258) );
XOR2_X1 U992 ( .A(n1174), .B(KEYINPUT53), .Z(n1054) );
INV_X1 U993 ( .A(G131), .ZN(n1174) );
XOR2_X1 U994 ( .A(n1178), .B(n1260), .Z(n1257) );
NOR2_X1 U995 ( .A1(KEYINPUT2), .A2(n1261), .ZN(n1260) );
INV_X1 U996 ( .A(G101), .ZN(n1178) );
INV_X1 U997 ( .A(n1179), .ZN(n1010) );
XOR2_X1 U998 ( .A(n1007), .B(KEYINPUT50), .Z(n1179) );
NAND2_X1 U999 ( .A1(G221), .A2(n1199), .ZN(n1007) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1200), .ZN(n1199) );
NAND2_X1 U1001 ( .A1(n993), .A2(n1262), .ZN(n1195) );
NAND4_X1 U1002 ( .A1(n1076), .A2(G902), .A3(G953), .A4(n1182), .ZN(n1262) );
XNOR2_X1 U1003 ( .A(G898), .B(KEYINPUT9), .ZN(n1076) );
NAND3_X1 U1004 ( .A1(n1182), .A2(n1057), .A3(G952), .ZN(n993) );
INV_X1 U1005 ( .A(G953), .ZN(n1057) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1182) );
NAND2_X1 U1007 ( .A1(n1263), .A2(n1264), .ZN(n1152) );
NAND3_X1 U1008 ( .A1(n1022), .A2(n1021), .A3(n1265), .ZN(n1264) );
INV_X1 U1009 ( .A(KEYINPUT36), .ZN(n1265) );
NAND2_X1 U1010 ( .A1(KEYINPUT36), .A2(n1142), .ZN(n1263) );
NOR2_X1 U1011 ( .A1(n1022), .A2(n1035), .ZN(n1142) );
INV_X1 U1012 ( .A(n1021), .ZN(n1035) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1266), .ZN(n1021) );
XNOR2_X1 U1014 ( .A(n1037), .B(n1038), .ZN(n1022) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1266), .ZN(n1038) );
NAND2_X1 U1016 ( .A1(n1222), .A2(n1200), .ZN(n1266) );
INV_X1 U1017 ( .A(G237), .ZN(n1222) );
AND2_X1 U1018 ( .A1(n1267), .A2(n1200), .ZN(n1037) );
INV_X1 U1019 ( .A(G902), .ZN(n1200) );
XOR2_X1 U1020 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U1021 ( .A(n1270), .B(n1052), .Z(n1269) );
XOR2_X1 U1022 ( .A(n1271), .B(n1207), .Z(n1052) );
XNOR2_X1 U1023 ( .A(G128), .B(KEYINPUT47), .ZN(n1207) );
XOR2_X1 U1024 ( .A(n1167), .B(G146), .Z(n1271) );
INV_X1 U1025 ( .A(G143), .ZN(n1167) );
NAND2_X1 U1026 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
OR2_X1 U1027 ( .A1(KEYINPUT55), .A2(n1159), .ZN(n1273) );
NAND2_X1 U1028 ( .A1(KEYINPUT34), .A2(n1159), .ZN(n1272) );
XNOR2_X1 U1029 ( .A(n1079), .B(n1274), .ZN(n1159) );
NOR4_X1 U1030 ( .A1(n1275), .A2(n1276), .A3(KEYINPUT22), .A4(n1085), .ZN(n1274) );
NOR2_X1 U1031 ( .A1(n1083), .A2(n1084), .ZN(n1085) );
NOR2_X1 U1032 ( .A1(KEYINPUT40), .A2(n1084), .ZN(n1276) );
AND3_X1 U1033 ( .A1(n1084), .A2(n1083), .A3(KEYINPUT40), .ZN(n1275) );
XOR2_X1 U1034 ( .A(G101), .B(n1261), .Z(n1083) );
XNOR2_X1 U1035 ( .A(G107), .B(G104), .ZN(n1261) );
XOR2_X1 U1036 ( .A(n1220), .B(n1219), .Z(n1084) );
XNOR2_X1 U1037 ( .A(G113), .B(KEYINPUT25), .ZN(n1219) );
XOR2_X1 U1038 ( .A(G116), .B(n1277), .Z(n1220) );
XOR2_X1 U1039 ( .A(KEYINPUT30), .B(G119), .Z(n1277) );
XNOR2_X1 U1040 ( .A(n1211), .B(G122), .ZN(n1079) );
INV_X1 U1041 ( .A(G110), .ZN(n1211) );
XNOR2_X1 U1042 ( .A(G125), .B(n1162), .ZN(n1268) );
AND2_X1 U1043 ( .A1(G224), .A2(n1221), .ZN(n1162) );
XNOR2_X1 U1044 ( .A(G953), .B(KEYINPUT29), .ZN(n1221) );
endmodule


