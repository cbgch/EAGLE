//Key = 0100001001111100001001111010110101100101111110001101001010110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XNOR2_X1 U734 ( .A(G107), .B(n1005), .ZN(G9) );
NOR2_X1 U735 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR3_X1 U736 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
XOR2_X1 U737 ( .A(KEYINPUT44), .B(n1011), .Z(n1010) );
NAND3_X1 U738 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1008) );
NAND2_X1 U739 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND3_X1 U741 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND2_X1 U742 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NAND2_X1 U743 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
OR2_X1 U744 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1022) );
NAND2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
OR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U748 ( .A1(n1028), .A2(n1034), .A3(n1024), .ZN(n1017) );
NAND2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U750 ( .A1(n1021), .A2(n1037), .ZN(n1036) );
NAND2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U752 ( .A1(n1019), .A2(n1040), .ZN(n1035) );
NAND2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
INV_X1 U755 ( .A(n1045), .ZN(n1015) );
AND3_X1 U756 ( .A1(n1012), .A2(n1013), .A3(n1046), .ZN(n1006) );
NAND4_X1 U757 ( .A1(n1047), .A2(n1032), .A3(n1048), .A4(n1049), .ZN(n1012) );
NOR4_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
XNOR2_X1 U759 ( .A(n1054), .B(n1055), .ZN(n1051) );
NOR2_X1 U760 ( .A1(KEYINPUT55), .A2(n1056), .ZN(n1055) );
NAND3_X1 U761 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1050) );
XOR2_X1 U762 ( .A(n1060), .B(KEYINPUT60), .Z(n1059) );
OR2_X1 U763 ( .A1(n1061), .A2(G472), .ZN(n1060) );
OR2_X1 U764 ( .A1(G478), .A2(KEYINPUT31), .ZN(n1058) );
NAND3_X1 U765 ( .A1(G478), .A2(n1062), .A3(KEYINPUT31), .ZN(n1057) );
NOR3_X1 U766 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1048) );
INV_X1 U767 ( .A(n1066), .ZN(n1063) );
NAND2_X1 U768 ( .A1(G472), .A2(n1061), .ZN(n1047) );
XNOR2_X1 U769 ( .A(n1067), .B(KEYINPUT63), .ZN(n1061) );
XOR2_X1 U770 ( .A(n1068), .B(n1069), .Z(G72) );
NOR2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
AND2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U773 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1070) );
NOR2_X1 U774 ( .A1(G900), .A2(n1013), .ZN(n1074) );
AND2_X1 U775 ( .A1(n1075), .A2(n1013), .ZN(n1073) );
NAND3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
INV_X1 U777 ( .A(n1079), .ZN(n1076) );
XNOR2_X1 U778 ( .A(n1080), .B(n1081), .ZN(n1072) );
NOR2_X1 U779 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U780 ( .A1(KEYINPUT46), .A2(n1084), .ZN(n1083) );
NOR2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
INV_X1 U782 ( .A(KEYINPUT46), .ZN(n1085) );
XNOR2_X1 U783 ( .A(n1087), .B(n1088), .ZN(n1080) );
NOR2_X1 U784 ( .A1(KEYINPUT53), .A2(n1089), .ZN(n1068) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1013), .ZN(n1089) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1091), .A2(n1092), .ZN(G69) );
NAND2_X1 U788 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U789 ( .A1(G953), .A2(n1095), .ZN(n1094) );
NAND3_X1 U790 ( .A1(G953), .A2(n1096), .A3(n1097), .ZN(n1091) );
XNOR2_X1 U791 ( .A(n1093), .B(KEYINPUT45), .ZN(n1097) );
XNOR2_X1 U792 ( .A(n1098), .B(n1099), .ZN(n1093) );
NOR3_X1 U793 ( .A1(n1100), .A2(KEYINPUT38), .A3(G953), .ZN(n1099) );
XNOR2_X1 U794 ( .A(n1101), .B(KEYINPUT58), .ZN(n1100) );
NAND2_X1 U795 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
NAND2_X1 U796 ( .A1(G953), .A2(n1104), .ZN(n1103) );
XOR2_X1 U797 ( .A(n1105), .B(n1106), .Z(n1102) );
NOR2_X1 U798 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U799 ( .A(KEYINPUT56), .B(KEYINPUT35), .ZN(n1107) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1096) );
NOR2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U802 ( .A(n1111), .B(KEYINPUT39), .Z(n1110) );
NAND2_X1 U803 ( .A1(n1112), .A2(n1046), .ZN(n1111) );
INV_X1 U804 ( .A(G952), .ZN(n1046) );
XNOR2_X1 U805 ( .A(KEYINPUT32), .B(n1013), .ZN(n1112) );
XNOR2_X1 U806 ( .A(n1113), .B(n1114), .ZN(n1109) );
NOR2_X1 U807 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1118), .ZN(G63) );
XOR2_X1 U809 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U810 ( .A1(KEYINPUT48), .A2(n1121), .ZN(n1120) );
NAND2_X1 U811 ( .A1(n1122), .A2(G478), .ZN(n1119) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1123), .ZN(G60) );
XOR2_X1 U813 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U814 ( .A1(n1126), .A2(n1116), .ZN(n1125) );
NAND2_X1 U815 ( .A1(KEYINPUT28), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U816 ( .A(G104), .B(n1128), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1117), .A2(n1129), .ZN(G57) );
XOR2_X1 U818 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U819 ( .A(G101), .B(n1132), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1130) );
AND2_X1 U821 ( .A1(G472), .A2(n1122), .ZN(n1134) );
INV_X1 U822 ( .A(n1116), .ZN(n1122) );
NAND2_X1 U823 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NAND2_X1 U824 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U825 ( .A(KEYINPUT12), .B(n1139), .Z(n1135) );
NOR2_X1 U826 ( .A1(n1137), .A2(n1138), .ZN(n1139) );
NOR2_X1 U827 ( .A1(n1117), .A2(n1140), .ZN(G54) );
XOR2_X1 U828 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U829 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U830 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U831 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U832 ( .A1(n1149), .A2(KEYINPUT50), .ZN(n1147) );
INV_X1 U833 ( .A(n1150), .ZN(n1149) );
NOR2_X1 U834 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
NOR3_X1 U835 ( .A1(n1153), .A2(n1151), .A3(n1152), .ZN(n1143) );
INV_X1 U836 ( .A(KEYINPUT43), .ZN(n1152) );
XOR2_X1 U837 ( .A(n1154), .B(KEYINPUT51), .Z(n1151) );
XOR2_X1 U838 ( .A(n1155), .B(n1148), .Z(n1153) );
XNOR2_X1 U839 ( .A(n1156), .B(KEYINPUT24), .ZN(n1148) );
NOR2_X1 U840 ( .A1(KEYINPUT50), .A2(n1150), .ZN(n1155) );
NOR2_X1 U841 ( .A1(n1056), .A2(n1116), .ZN(n1141) );
NOR2_X1 U842 ( .A1(n1117), .A2(n1157), .ZN(G51) );
XOR2_X1 U843 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U844 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U845 ( .A1(n1162), .A2(n1116), .ZN(n1160) );
NAND2_X1 U846 ( .A1(G902), .A2(n1163), .ZN(n1116) );
NAND2_X1 U847 ( .A1(n1101), .A2(n1011), .ZN(n1163) );
AND2_X1 U848 ( .A1(n1078), .A2(n1164), .ZN(n1011) );
XOR2_X1 U849 ( .A(KEYINPUT30), .B(n1165), .Z(n1164) );
NOR2_X1 U850 ( .A1(n1166), .A2(n1079), .ZN(n1165) );
NAND3_X1 U851 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1079) );
NAND4_X1 U852 ( .A1(n1170), .A2(n1026), .A3(n1171), .A4(n1024), .ZN(n1169) );
NOR2_X1 U853 ( .A1(n1041), .A2(n1039), .ZN(n1171) );
INV_X1 U854 ( .A(n1172), .ZN(n1039) );
INV_X1 U855 ( .A(n1173), .ZN(n1041) );
XOR2_X1 U856 ( .A(n1174), .B(KEYINPUT17), .Z(n1170) );
XOR2_X1 U857 ( .A(n1077), .B(KEYINPUT9), .Z(n1166) );
AND4_X1 U858 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1078) );
INV_X1 U859 ( .A(n1009), .ZN(n1101) );
NAND2_X1 U860 ( .A1(n1179), .A2(n1180), .ZN(n1009) );
NOR4_X1 U861 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
AND4_X1 U862 ( .A1(n1005), .A2(n1185), .A3(n1186), .A4(n1128), .ZN(n1179) );
NAND3_X1 U863 ( .A1(n1187), .A2(n1019), .A3(n1026), .ZN(n1128) );
NAND3_X1 U864 ( .A1(n1187), .A2(n1019), .A3(n1027), .ZN(n1005) );
XNOR2_X1 U865 ( .A(KEYINPUT13), .B(n1188), .ZN(n1158) );
NOR2_X1 U866 ( .A1(n1013), .A2(G952), .ZN(n1117) );
XNOR2_X1 U867 ( .A(G146), .B(n1175), .ZN(G48) );
NAND3_X1 U868 ( .A1(n1026), .A2(n1173), .A3(n1189), .ZN(n1175) );
XNOR2_X1 U869 ( .A(G143), .B(n1176), .ZN(G45) );
NAND4_X1 U870 ( .A1(n1190), .A2(n1173), .A3(n1191), .A4(n1192), .ZN(n1176) );
XNOR2_X1 U871 ( .A(G140), .B(n1177), .ZN(G42) );
NAND3_X1 U872 ( .A1(n1021), .A2(n1193), .A3(n1194), .ZN(n1177) );
XNOR2_X1 U873 ( .A(G137), .B(n1178), .ZN(G39) );
NAND3_X1 U874 ( .A1(n1028), .A2(n1021), .A3(n1189), .ZN(n1178) );
XNOR2_X1 U875 ( .A(G134), .B(n1167), .ZN(G36) );
NAND3_X1 U876 ( .A1(n1021), .A2(n1027), .A3(n1190), .ZN(n1167) );
XNOR2_X1 U877 ( .A(G131), .B(n1168), .ZN(G33) );
NAND3_X1 U878 ( .A1(n1026), .A2(n1021), .A3(n1190), .ZN(n1168) );
AND3_X1 U879 ( .A1(n1193), .A2(n1174), .A3(n1195), .ZN(n1190) );
INV_X1 U880 ( .A(n1052), .ZN(n1021) );
NAND2_X1 U881 ( .A1(n1044), .A2(n1196), .ZN(n1052) );
XOR2_X1 U882 ( .A(G128), .B(n1197), .Z(G30) );
NOR2_X1 U883 ( .A1(KEYINPUT47), .A2(n1077), .ZN(n1197) );
NAND3_X1 U884 ( .A1(n1027), .A2(n1173), .A3(n1189), .ZN(n1077) );
AND4_X1 U885 ( .A1(n1193), .A2(n1053), .A3(n1174), .A4(n1198), .ZN(n1189) );
XNOR2_X1 U886 ( .A(n1184), .B(n1199), .ZN(G3) );
NOR2_X1 U887 ( .A1(G101), .A2(KEYINPUT4), .ZN(n1199) );
AND3_X1 U888 ( .A1(n1187), .A2(n1195), .A3(n1028), .ZN(n1184) );
XNOR2_X1 U889 ( .A(G125), .B(n1200), .ZN(G27) );
NAND4_X1 U890 ( .A1(KEYINPUT6), .A2(n1194), .A3(n1024), .A4(n1173), .ZN(n1200) );
AND3_X1 U891 ( .A1(n1172), .A2(n1174), .A3(n1026), .ZN(n1194) );
NAND2_X1 U892 ( .A1(n1045), .A2(n1201), .ZN(n1174) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1203), .ZN(n1201) );
INV_X1 U894 ( .A(G900), .ZN(n1203) );
NAND3_X1 U895 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(G24) );
NAND2_X1 U896 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U897 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
INV_X1 U898 ( .A(KEYINPUT1), .ZN(n1210) );
NAND2_X1 U899 ( .A1(n1211), .A2(G122), .ZN(n1209) );
XNOR2_X1 U900 ( .A(n1207), .B(KEYINPUT0), .ZN(n1211) );
NAND2_X1 U901 ( .A1(KEYINPUT1), .A2(n1212), .ZN(n1204) );
NAND2_X1 U902 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR3_X1 U903 ( .A1(n1208), .A2(n1207), .A3(KEYINPUT0), .ZN(n1214) );
NAND2_X1 U904 ( .A1(KEYINPUT0), .A2(n1207), .ZN(n1213) );
INV_X1 U905 ( .A(n1186), .ZN(n1207) );
NAND3_X1 U906 ( .A1(n1024), .A2(n1215), .A3(n1216), .ZN(n1186) );
AND3_X1 U907 ( .A1(n1019), .A2(n1192), .A3(n1191), .ZN(n1216) );
NAND2_X1 U908 ( .A1(n1217), .A2(n1218), .ZN(n1019) );
OR2_X1 U909 ( .A1(n1038), .A2(KEYINPUT29), .ZN(n1218) );
INV_X1 U910 ( .A(n1195), .ZN(n1038) );
NAND3_X1 U911 ( .A1(n1219), .A2(n1220), .A3(KEYINPUT29), .ZN(n1217) );
XOR2_X1 U912 ( .A(G119), .B(n1221), .Z(G21) );
NOR2_X1 U913 ( .A1(KEYINPUT27), .A2(n1185), .ZN(n1221) );
NAND4_X1 U914 ( .A1(n1024), .A2(n1028), .A3(n1222), .A4(n1215), .ZN(n1185) );
NOR2_X1 U915 ( .A1(n1219), .A2(n1220), .ZN(n1222) );
XOR2_X1 U916 ( .A(G116), .B(n1183), .Z(G18) );
AND2_X1 U917 ( .A1(n1223), .A2(n1027), .ZN(n1183) );
NOR2_X1 U918 ( .A1(n1191), .A2(n1224), .ZN(n1027) );
XNOR2_X1 U919 ( .A(G113), .B(n1225), .ZN(G15) );
NOR2_X1 U920 ( .A1(n1182), .A2(KEYINPUT20), .ZN(n1225) );
AND2_X1 U921 ( .A1(n1026), .A2(n1223), .ZN(n1182) );
AND3_X1 U922 ( .A1(n1195), .A2(n1215), .A3(n1024), .ZN(n1223) );
NOR2_X1 U923 ( .A1(n1033), .A2(n1226), .ZN(n1024) );
INV_X1 U924 ( .A(n1032), .ZN(n1226) );
NOR2_X1 U925 ( .A1(n1053), .A2(n1219), .ZN(n1195) );
INV_X1 U926 ( .A(n1198), .ZN(n1219) );
AND2_X1 U927 ( .A1(n1224), .A2(n1191), .ZN(n1026) );
XOR2_X1 U928 ( .A(n1181), .B(n1227), .Z(G12) );
NOR2_X1 U929 ( .A1(KEYINPUT61), .A2(n1228), .ZN(n1227) );
INV_X1 U930 ( .A(G110), .ZN(n1228) );
AND3_X1 U931 ( .A1(n1172), .A2(n1187), .A3(n1028), .ZN(n1181) );
NOR2_X1 U932 ( .A1(n1192), .A2(n1191), .ZN(n1028) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1066), .ZN(n1191) );
NAND3_X1 U934 ( .A1(n1126), .A2(n1230), .A3(n1127), .ZN(n1066) );
INV_X1 U935 ( .A(G475), .ZN(n1126) );
XOR2_X1 U936 ( .A(KEYINPUT26), .B(n1064), .Z(n1229) );
AND2_X1 U937 ( .A1(G475), .A2(n1231), .ZN(n1064) );
NAND2_X1 U938 ( .A1(n1127), .A2(n1230), .ZN(n1231) );
XOR2_X1 U939 ( .A(n1232), .B(n1233), .Z(n1127) );
NOR3_X1 U940 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NOR2_X1 U941 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
AND3_X1 U942 ( .A1(n1238), .A2(n1239), .A3(n1237), .ZN(n1235) );
AND2_X1 U943 ( .A1(n1240), .A2(KEYINPUT54), .ZN(n1237) );
XNOR2_X1 U944 ( .A(n1241), .B(n1242), .ZN(n1238) );
XNOR2_X1 U945 ( .A(n1243), .B(G131), .ZN(n1242) );
INV_X1 U946 ( .A(G143), .ZN(n1243) );
NAND2_X1 U947 ( .A1(G214), .A2(n1244), .ZN(n1241) );
NOR2_X1 U948 ( .A1(n1240), .A2(n1239), .ZN(n1234) );
INV_X1 U949 ( .A(KEYINPUT16), .ZN(n1239) );
XOR2_X1 U950 ( .A(n1245), .B(G146), .Z(n1240) );
NAND2_X1 U951 ( .A1(KEYINPUT21), .A2(n1084), .ZN(n1245) );
XNOR2_X1 U952 ( .A(n1246), .B(G140), .ZN(n1084) );
NAND2_X1 U953 ( .A1(n1247), .A2(KEYINPUT18), .ZN(n1232) );
XOR2_X1 U954 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U955 ( .A(G104), .B(G122), .ZN(n1248) );
INV_X1 U956 ( .A(n1224), .ZN(n1192) );
NOR2_X1 U957 ( .A1(n1065), .A2(n1250), .ZN(n1224) );
AND2_X1 U958 ( .A1(G478), .A2(n1062), .ZN(n1250) );
NOR2_X1 U959 ( .A1(n1062), .A2(G478), .ZN(n1065) );
OR2_X1 U960 ( .A1(n1121), .A2(G902), .ZN(n1062) );
XOR2_X1 U961 ( .A(n1251), .B(n1252), .Z(n1121) );
AND2_X1 U962 ( .A1(n1253), .A2(G217), .ZN(n1252) );
NAND2_X1 U963 ( .A1(KEYINPUT40), .A2(n1254), .ZN(n1251) );
XOR2_X1 U964 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U965 ( .A(G107), .B(n1257), .Z(n1256) );
XOR2_X1 U966 ( .A(G116), .B(n1258), .Z(n1255) );
XNOR2_X1 U967 ( .A(G134), .B(n1208), .ZN(n1258) );
AND2_X1 U968 ( .A1(n1193), .A2(n1215), .ZN(n1187) );
AND2_X1 U969 ( .A1(n1173), .A2(n1259), .ZN(n1215) );
NAND2_X1 U970 ( .A1(n1045), .A2(n1260), .ZN(n1259) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1104), .ZN(n1260) );
INV_X1 U972 ( .A(G898), .ZN(n1104) );
NAND3_X1 U973 ( .A1(n1202), .A2(n1013), .A3(G952), .ZN(n1045) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1202) );
NOR2_X1 U975 ( .A1(n1044), .A2(n1043), .ZN(n1173) );
INV_X1 U976 ( .A(n1196), .ZN(n1043) );
NAND2_X1 U977 ( .A1(G214), .A2(n1261), .ZN(n1196) );
XNOR2_X1 U978 ( .A(n1262), .B(n1162), .ZN(n1044) );
NAND2_X1 U979 ( .A1(G210), .A2(n1261), .ZN(n1162) );
NAND2_X1 U980 ( .A1(n1263), .A2(n1230), .ZN(n1261) );
INV_X1 U981 ( .A(G237), .ZN(n1263) );
NAND2_X1 U982 ( .A1(n1264), .A2(n1230), .ZN(n1262) );
XOR2_X1 U983 ( .A(n1265), .B(n1161), .Z(n1264) );
XNOR2_X1 U984 ( .A(n1266), .B(n1267), .ZN(n1161) );
XNOR2_X1 U985 ( .A(n1246), .B(n1268), .ZN(n1267) );
NOR2_X1 U986 ( .A1(G953), .A2(n1095), .ZN(n1268) );
INV_X1 U987 ( .A(G224), .ZN(n1095) );
XNOR2_X1 U988 ( .A(KEYINPUT37), .B(n1269), .ZN(n1265) );
NOR2_X1 U989 ( .A1(KEYINPUT19), .A2(n1188), .ZN(n1269) );
NAND3_X1 U990 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1188) );
NAND2_X1 U991 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U992 ( .A1(KEYINPUT10), .A2(n1275), .ZN(n1274) );
XOR2_X1 U993 ( .A(n1105), .B(KEYINPUT3), .Z(n1273) );
NAND4_X1 U994 ( .A1(n1275), .A2(n1276), .A3(KEYINPUT10), .A4(n1277), .ZN(n1271) );
XNOR2_X1 U995 ( .A(KEYINPUT3), .B(n1105), .ZN(n1276) );
XOR2_X1 U996 ( .A(n1278), .B(n1279), .Z(n1105) );
XOR2_X1 U997 ( .A(n1137), .B(n1280), .Z(n1279) );
XOR2_X1 U998 ( .A(n1281), .B(G107), .Z(n1278) );
NAND2_X1 U999 ( .A1(KEYINPUT62), .A2(n1282), .ZN(n1281) );
INV_X1 U1000 ( .A(G104), .ZN(n1282) );
OR2_X1 U1001 ( .A1(n1275), .A2(n1277), .ZN(n1270) );
INV_X1 U1002 ( .A(KEYINPUT14), .ZN(n1277) );
XNOR2_X1 U1003 ( .A(n1108), .B(KEYINPUT25), .ZN(n1275) );
XNOR2_X1 U1004 ( .A(G110), .B(n1208), .ZN(n1108) );
INV_X1 U1005 ( .A(G122), .ZN(n1208) );
INV_X1 U1006 ( .A(n1030), .ZN(n1193) );
NAND2_X1 U1007 ( .A1(n1033), .A2(n1032), .ZN(n1030) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1283), .ZN(n1032) );
XOR2_X1 U1009 ( .A(n1054), .B(n1056), .Z(n1033) );
INV_X1 U1010 ( .A(G469), .ZN(n1056) );
NAND2_X1 U1011 ( .A1(n1284), .A2(n1230), .ZN(n1054) );
XNOR2_X1 U1012 ( .A(n1285), .B(n1156), .ZN(n1284) );
XOR2_X1 U1013 ( .A(n1286), .B(n1287), .Z(n1156) );
XNOR2_X1 U1014 ( .A(n1288), .B(n1289), .ZN(n1287) );
NOR2_X1 U1015 ( .A1(KEYINPUT15), .A2(n1280), .ZN(n1288) );
XNOR2_X1 U1016 ( .A(G101), .B(KEYINPUT11), .ZN(n1280) );
XNOR2_X1 U1017 ( .A(G104), .B(n1290), .ZN(n1286) );
XOR2_X1 U1018 ( .A(KEYINPUT36), .B(G107), .Z(n1290) );
NAND2_X1 U1019 ( .A1(n1291), .A2(KEYINPUT41), .ZN(n1285) );
XNOR2_X1 U1020 ( .A(n1154), .B(n1150), .ZN(n1291) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1013), .ZN(n1150) );
XNOR2_X1 U1022 ( .A(G110), .B(n1292), .ZN(n1154) );
XOR2_X1 U1023 ( .A(KEYINPUT23), .B(G140), .Z(n1292) );
NOR2_X1 U1024 ( .A1(n1198), .A2(n1220), .ZN(n1172) );
INV_X1 U1025 ( .A(n1053), .ZN(n1220) );
XOR2_X1 U1026 ( .A(n1293), .B(n1115), .Z(n1053) );
NAND2_X1 U1027 ( .A1(G217), .A2(n1283), .ZN(n1115) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1230), .ZN(n1283) );
NAND2_X1 U1029 ( .A1(n1113), .A2(n1230), .ZN(n1293) );
XNOR2_X1 U1030 ( .A(n1294), .B(n1295), .ZN(n1113) );
XOR2_X1 U1031 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND2_X1 U1032 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
OR2_X1 U1033 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U1034 ( .A(n1302), .B(KEYINPUT57), .Z(n1298) );
NAND2_X1 U1035 ( .A1(n1301), .A2(n1300), .ZN(n1302) );
XOR2_X1 U1036 ( .A(G110), .B(n1303), .Z(n1300) );
XOR2_X1 U1037 ( .A(G128), .B(G119), .Z(n1303) );
XNOR2_X1 U1038 ( .A(n1304), .B(G146), .ZN(n1301) );
NAND2_X1 U1039 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1040 ( .A1(G140), .A2(n1246), .ZN(n1306) );
XOR2_X1 U1041 ( .A(n1086), .B(KEYINPUT7), .Z(n1305) );
OR2_X1 U1042 ( .A1(n1246), .A2(G140), .ZN(n1086) );
INV_X1 U1043 ( .A(G125), .ZN(n1246) );
NAND2_X1 U1044 ( .A1(n1307), .A2(KEYINPUT34), .ZN(n1296) );
XNOR2_X1 U1045 ( .A(G137), .B(KEYINPUT8), .ZN(n1307) );
NAND2_X1 U1046 ( .A1(G221), .A2(n1253), .ZN(n1294) );
AND2_X1 U1047 ( .A1(G234), .A2(n1013), .ZN(n1253) );
INV_X1 U1048 ( .A(G953), .ZN(n1013) );
NAND3_X1 U1049 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1198) );
NAND2_X1 U1050 ( .A1(G472), .A2(n1311), .ZN(n1310) );
OR3_X1 U1051 ( .A1(n1311), .A2(G472), .A3(KEYINPUT5), .ZN(n1309) );
AND2_X1 U1052 ( .A1(KEYINPUT42), .A2(n1067), .ZN(n1311) );
NAND2_X1 U1053 ( .A1(KEYINPUT5), .A2(n1312), .ZN(n1308) );
OR2_X1 U1054 ( .A1(n1067), .A2(G472), .ZN(n1312) );
NAND2_X1 U1055 ( .A1(n1313), .A2(n1230), .ZN(n1067) );
INV_X1 U1056 ( .A(G902), .ZN(n1230) );
XNOR2_X1 U1057 ( .A(n1314), .B(n1137), .ZN(n1313) );
XOR2_X1 U1058 ( .A(n1315), .B(n1249), .Z(n1137) );
XOR2_X1 U1059 ( .A(G113), .B(KEYINPUT33), .Z(n1249) );
XNOR2_X1 U1060 ( .A(G116), .B(G119), .ZN(n1315) );
XOR2_X1 U1061 ( .A(n1316), .B(n1317), .Z(n1314) );
NOR3_X1 U1062 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1317) );
NOR2_X1 U1063 ( .A1(G101), .A2(n1321), .ZN(n1320) );
AND3_X1 U1064 ( .A1(G101), .A2(n1321), .A3(KEYINPUT22), .ZN(n1319) );
AND2_X1 U1065 ( .A1(KEYINPUT59), .A2(n1132), .ZN(n1321) );
NOR2_X1 U1066 ( .A1(KEYINPUT22), .A2(n1132), .ZN(n1318) );
NAND2_X1 U1067 ( .A1(G210), .A2(n1244), .ZN(n1132) );
NOR2_X1 U1068 ( .A1(G953), .A2(G237), .ZN(n1244) );
NAND2_X1 U1069 ( .A1(n1289), .A2(n1322), .ZN(n1316) );
XOR2_X1 U1070 ( .A(KEYINPUT52), .B(KEYINPUT49), .Z(n1322) );
INV_X1 U1071 ( .A(n1138), .ZN(n1289) );
XNOR2_X1 U1072 ( .A(n1087), .B(n1323), .ZN(n1138) );
NOR2_X1 U1073 ( .A1(KEYINPUT2), .A2(n1088), .ZN(n1323) );
INV_X1 U1074 ( .A(G131), .ZN(n1088) );
XOR2_X1 U1075 ( .A(n1266), .B(n1324), .Z(n1087) );
XOR2_X1 U1076 ( .A(G137), .B(G134), .Z(n1324) );
XNOR2_X1 U1077 ( .A(G146), .B(n1257), .ZN(n1266) );
XOR2_X1 U1078 ( .A(G128), .B(G143), .Z(n1257) );
endmodule


