//Key = 1111010110110000000101100100001000101011011111010101000110111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350;

XNOR2_X1 U731 ( .A(G107), .B(n1020), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U733 ( .A1(G953), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1022) );
NOR2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
INV_X1 U735 ( .A(n1028), .ZN(n1027) );
NOR2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1026) );
NOR3_X1 U737 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1034) );
NOR2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U743 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR4_X1 U744 ( .A1(n1046), .A2(n1047), .A3(n1037), .A4(n1041), .ZN(n1029) );
NOR3_X1 U745 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
NOR2_X1 U747 ( .A1(n1053), .A2(n1050), .ZN(n1046) );
AND2_X1 U748 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR3_X1 U751 ( .A1(n1023), .A2(G953), .A3(G952), .ZN(n1021) );
AND4_X1 U752 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1023) );
NOR4_X1 U753 ( .A1(n1064), .A2(n1058), .A3(n1065), .A4(n1066), .ZN(n1063) );
XNOR2_X1 U754 ( .A(n1067), .B(n1068), .ZN(n1066) );
NAND2_X1 U755 ( .A1(KEYINPUT55), .A2(n1069), .ZN(n1067) );
AND2_X1 U756 ( .A1(n1070), .A2(G472), .ZN(n1065) );
NOR2_X1 U757 ( .A1(n1071), .A2(n1072), .ZN(n1062) );
INV_X1 U758 ( .A(n1051), .ZN(n1072) );
XOR2_X1 U759 ( .A(n1073), .B(n1074), .Z(n1071) );
XNOR2_X1 U760 ( .A(n1075), .B(n1076), .ZN(n1060) );
XNOR2_X1 U761 ( .A(KEYINPUT15), .B(n1077), .ZN(n1076) );
XOR2_X1 U762 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U763 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U764 ( .A1(G227), .A2(n1082), .ZN(n1080) );
NOR3_X1 U765 ( .A1(KEYINPUT14), .A2(n1083), .A3(n1084), .ZN(n1078) );
NOR2_X1 U766 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
AND3_X1 U767 ( .A1(n1086), .A2(n1087), .A3(n1085), .ZN(n1083) );
XNOR2_X1 U768 ( .A(n1088), .B(n1089), .ZN(n1085) );
XOR2_X1 U769 ( .A(G140), .B(G125), .Z(n1089) );
NAND2_X1 U770 ( .A1(n1090), .A2(KEYINPUT10), .ZN(n1088) );
XOR2_X1 U771 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U772 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U773 ( .A(KEYINPUT24), .B(n1095), .Z(n1094) );
NOR2_X1 U774 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
AND2_X1 U775 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND3_X1 U776 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U777 ( .A1(KEYINPUT54), .A2(G134), .ZN(n1100) );
NAND3_X1 U778 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1099) );
INV_X1 U779 ( .A(KEYINPUT54), .ZN(n1102) );
OR2_X1 U780 ( .A1(n1103), .A2(n1101), .ZN(n1098) );
NOR2_X1 U781 ( .A1(n1104), .A2(G134), .ZN(n1101) );
INV_X1 U782 ( .A(KEYINPUT45), .ZN(n1104) );
INV_X1 U783 ( .A(n1081), .ZN(n1087) );
NAND2_X1 U784 ( .A1(n1082), .A2(n1105), .ZN(n1086) );
NAND3_X1 U785 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
XOR2_X1 U786 ( .A(n1109), .B(KEYINPUT57), .Z(n1108) );
XOR2_X1 U787 ( .A(KEYINPUT62), .B(n1110), .Z(n1107) );
NAND2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(G69) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1082), .ZN(n1112) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U791 ( .A1(KEYINPUT36), .A2(n1116), .ZN(n1115) );
NAND2_X1 U792 ( .A1(n1117), .A2(G953), .ZN(n1111) );
XOR2_X1 U793 ( .A(n1114), .B(n1118), .Z(n1117) );
AND2_X1 U794 ( .A1(G224), .A2(G898), .ZN(n1118) );
NAND2_X1 U795 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U797 ( .A(n1082), .B(KEYINPUT47), .Z(n1121) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NOR2_X1 U801 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XOR2_X1 U802 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND3_X1 U803 ( .A1(n1132), .A2(n1025), .A3(G478), .ZN(n1130) );
XOR2_X1 U804 ( .A(KEYINPUT20), .B(n1133), .Z(n1132) );
NOR2_X1 U805 ( .A1(n1123), .A2(n1134), .ZN(G60) );
XOR2_X1 U806 ( .A(n1135), .B(n1136), .Z(n1134) );
AND2_X1 U807 ( .A1(G475), .A2(n1137), .ZN(n1136) );
XOR2_X1 U808 ( .A(G104), .B(n1138), .Z(G6) );
AND2_X1 U809 ( .A1(n1139), .A2(n1039), .ZN(n1138) );
NOR2_X1 U810 ( .A1(n1123), .A2(n1140), .ZN(G57) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U812 ( .A(n1143), .B(n1144), .ZN(n1142) );
NAND2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
OR2_X1 U814 ( .A1(KEYINPUT5), .A2(n1147), .ZN(n1146) );
NAND2_X1 U815 ( .A1(KEYINPUT43), .A2(n1147), .ZN(n1145) );
NAND2_X1 U816 ( .A1(n1137), .A2(G472), .ZN(n1147) );
XOR2_X1 U817 ( .A(n1148), .B(n1149), .Z(n1141) );
NOR2_X1 U818 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U819 ( .A(n1152), .B(KEYINPUT63), .Z(n1151) );
NAND2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NAND2_X1 U822 ( .A1(KEYINPUT60), .A2(n1155), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1123), .A2(n1156), .ZN(G54) );
XOR2_X1 U824 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U825 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U826 ( .A1(G469), .A2(n1137), .ZN(n1159) );
INV_X1 U827 ( .A(n1128), .ZN(n1137) );
XOR2_X1 U828 ( .A(KEYINPUT40), .B(G140), .Z(n1157) );
NOR2_X1 U829 ( .A1(n1123), .A2(n1161), .ZN(G51) );
XOR2_X1 U830 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U831 ( .A(n1119), .B(n1164), .ZN(n1163) );
NAND2_X1 U832 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
INV_X1 U834 ( .A(KEYINPUT46), .ZN(n1168) );
XOR2_X1 U835 ( .A(n1169), .B(G125), .Z(n1167) );
NAND3_X1 U836 ( .A1(G125), .A2(n1169), .A3(KEYINPUT46), .ZN(n1165) );
XNOR2_X1 U837 ( .A(n1170), .B(G122), .ZN(n1119) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1162) );
XNOR2_X1 U839 ( .A(KEYINPUT28), .B(n1173), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1077), .A2(n1128), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1133), .A2(n1025), .ZN(n1128) );
NAND4_X1 U842 ( .A1(n1110), .A2(n1174), .A3(n1106), .A4(n1109), .ZN(n1025) );
AND3_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1106) );
OR2_X1 U844 ( .A1(n1178), .A2(n1031), .ZN(n1177) );
INV_X1 U845 ( .A(n1053), .ZN(n1031) );
INV_X1 U846 ( .A(n1116), .ZN(n1174) );
NAND4_X1 U847 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1116) );
AND4_X1 U848 ( .A1(n1020), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1182) );
NAND2_X1 U849 ( .A1(n1038), .A2(n1139), .ZN(n1020) );
NOR3_X1 U850 ( .A1(n1186), .A2(n1187), .A3(n1033), .ZN(n1139) );
NOR2_X1 U851 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
NOR2_X1 U852 ( .A1(n1056), .A2(n1190), .ZN(n1189) );
NOR4_X1 U853 ( .A1(n1186), .A2(n1191), .A3(n1041), .A4(n1192), .ZN(n1188) );
XOR2_X1 U854 ( .A(KEYINPUT48), .B(n1187), .Z(n1192) );
NAND4_X1 U855 ( .A1(n1193), .A2(n1194), .A3(n1039), .A4(n1195), .ZN(n1179) );
NOR2_X1 U856 ( .A1(n1187), .A2(n1033), .ZN(n1195) );
NAND2_X1 U857 ( .A1(KEYINPUT8), .A2(n1186), .ZN(n1194) );
NAND2_X1 U858 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
INV_X1 U859 ( .A(KEYINPUT8), .ZN(n1197) );
NAND2_X1 U860 ( .A1(n1043), .A2(n1056), .ZN(n1196) );
AND4_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1110) );
XOR2_X1 U862 ( .A(G902), .B(KEYINPUT52), .Z(n1133) );
NOR2_X1 U863 ( .A1(n1082), .A2(G952), .ZN(n1123) );
XOR2_X1 U864 ( .A(n1202), .B(G146), .Z(G48) );
NAND2_X1 U865 ( .A1(KEYINPUT34), .A2(n1175), .ZN(n1202) );
NAND3_X1 U866 ( .A1(n1203), .A2(n1052), .A3(n1204), .ZN(n1175) );
XOR2_X1 U867 ( .A(n1205), .B(G143), .Z(G45) );
NAND2_X1 U868 ( .A1(KEYINPUT21), .A2(n1176), .ZN(n1205) );
NAND3_X1 U869 ( .A1(n1049), .A2(n1203), .A3(n1206), .ZN(n1176) );
AND3_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1210), .B(n1211), .Z(G42) );
NAND2_X1 U872 ( .A1(KEYINPUT11), .A2(G140), .ZN(n1211) );
NAND2_X1 U873 ( .A1(n1212), .A2(n1053), .ZN(n1210) );
XOR2_X1 U874 ( .A(n1178), .B(KEYINPUT42), .Z(n1212) );
NAND3_X1 U875 ( .A1(n1043), .A2(n1213), .A3(n1204), .ZN(n1178) );
XOR2_X1 U876 ( .A(n1103), .B(n1109), .Z(G39) );
NAND3_X1 U877 ( .A1(n1214), .A2(n1052), .A3(n1215), .ZN(n1109) );
XNOR2_X1 U878 ( .A(G134), .B(n1198), .ZN(G36) );
NAND3_X1 U879 ( .A1(n1214), .A2(n1038), .A3(n1049), .ZN(n1198) );
XOR2_X1 U880 ( .A(n1096), .B(n1199), .Z(G33) );
NAND3_X1 U881 ( .A1(n1214), .A2(n1039), .A3(n1049), .ZN(n1199) );
AND3_X1 U882 ( .A1(n1043), .A2(n1209), .A3(n1053), .ZN(n1214) );
NOR2_X1 U883 ( .A1(n1216), .A2(n1058), .ZN(n1053) );
XNOR2_X1 U884 ( .A(n1200), .B(n1217), .ZN(G30) );
NOR2_X1 U885 ( .A1(KEYINPUT16), .A2(n1218), .ZN(n1217) );
NAND3_X1 U886 ( .A1(n1038), .A2(n1203), .A3(n1219), .ZN(n1200) );
NOR3_X1 U887 ( .A1(n1051), .A2(n1213), .A3(n1220), .ZN(n1219) );
XNOR2_X1 U888 ( .A(G101), .B(n1221), .ZN(G3) );
NAND4_X1 U889 ( .A1(n1222), .A2(n1049), .A3(n1203), .A4(n1223), .ZN(n1221) );
INV_X1 U890 ( .A(n1186), .ZN(n1203) );
NAND2_X1 U891 ( .A1(n1224), .A2(n1043), .ZN(n1186) );
XOR2_X1 U892 ( .A(n1225), .B(n1201), .Z(G27) );
NAND4_X1 U893 ( .A1(n1204), .A2(n1061), .A3(n1224), .A4(n1213), .ZN(n1201) );
NOR3_X1 U894 ( .A1(n1051), .A2(n1220), .A3(n1226), .ZN(n1204) );
INV_X1 U895 ( .A(n1209), .ZN(n1220) );
NAND2_X1 U896 ( .A1(n1227), .A2(n1228), .ZN(n1209) );
NAND3_X1 U897 ( .A1(G902), .A2(n1028), .A3(n1081), .ZN(n1228) );
NOR2_X1 U898 ( .A1(G900), .A2(n1082), .ZN(n1081) );
XOR2_X1 U899 ( .A(n1229), .B(n1180), .Z(G24) );
NAND4_X1 U900 ( .A1(n1230), .A2(n1054), .A3(n1207), .A4(n1208), .ZN(n1180) );
INV_X1 U901 ( .A(n1033), .ZN(n1054) );
NAND2_X1 U902 ( .A1(n1213), .A2(n1051), .ZN(n1033) );
XNOR2_X1 U903 ( .A(G119), .B(n1185), .ZN(G21) );
NAND3_X1 U904 ( .A1(n1215), .A2(n1052), .A3(n1230), .ZN(n1185) );
XOR2_X1 U905 ( .A(n1231), .B(n1184), .Z(G18) );
NAND3_X1 U906 ( .A1(n1049), .A2(n1038), .A3(n1230), .ZN(n1184) );
NOR2_X1 U907 ( .A1(n1208), .A2(n1232), .ZN(n1038) );
XOR2_X1 U908 ( .A(n1183), .B(n1233), .Z(G15) );
NOR2_X1 U909 ( .A1(G113), .A2(KEYINPUT13), .ZN(n1233) );
NAND3_X1 U910 ( .A1(n1049), .A2(n1039), .A3(n1230), .ZN(n1183) );
NOR3_X1 U911 ( .A1(n1056), .A2(n1187), .A3(n1037), .ZN(n1230) );
INV_X1 U912 ( .A(n1061), .ZN(n1037) );
NOR2_X1 U913 ( .A1(n1044), .A2(n1234), .ZN(n1061) );
INV_X1 U914 ( .A(n1045), .ZN(n1234) );
INV_X1 U915 ( .A(n1223), .ZN(n1187) );
INV_X1 U916 ( .A(n1224), .ZN(n1056) );
INV_X1 U917 ( .A(n1226), .ZN(n1039) );
NAND2_X1 U918 ( .A1(n1235), .A2(n1208), .ZN(n1226) );
XOR2_X1 U919 ( .A(KEYINPUT23), .B(n1232), .Z(n1235) );
INV_X1 U920 ( .A(n1207), .ZN(n1232) );
INV_X1 U921 ( .A(n1191), .ZN(n1049) );
NAND2_X1 U922 ( .A1(n1051), .A2(n1052), .ZN(n1191) );
INV_X1 U923 ( .A(n1213), .ZN(n1052) );
XNOR2_X1 U924 ( .A(G110), .B(n1236), .ZN(G12) );
NAND2_X1 U925 ( .A1(n1237), .A2(n1224), .ZN(n1236) );
NOR2_X1 U926 ( .A1(n1059), .A2(n1058), .ZN(n1224) );
AND2_X1 U927 ( .A1(G214), .A2(n1238), .ZN(n1058) );
INV_X1 U928 ( .A(n1216), .ZN(n1059) );
NAND3_X1 U929 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1216) );
OR2_X1 U930 ( .A1(n1077), .A2(n1242), .ZN(n1241) );
NAND3_X1 U931 ( .A1(n1242), .A2(n1077), .A3(KEYINPUT7), .ZN(n1240) );
NAND2_X1 U932 ( .A1(KEYINPUT58), .A2(n1243), .ZN(n1242) );
NAND2_X1 U933 ( .A1(n1244), .A2(n1245), .ZN(n1239) );
INV_X1 U934 ( .A(KEYINPUT7), .ZN(n1245) );
NAND2_X1 U935 ( .A1(n1075), .A2(n1077), .ZN(n1244) );
NAND2_X1 U936 ( .A1(G210), .A2(n1238), .ZN(n1077) );
NAND2_X1 U937 ( .A1(n1246), .A2(n1247), .ZN(n1238) );
INV_X1 U938 ( .A(G237), .ZN(n1247) );
XOR2_X1 U939 ( .A(n1248), .B(KEYINPUT27), .Z(n1246) );
INV_X1 U940 ( .A(n1243), .ZN(n1075) );
NAND2_X1 U941 ( .A1(n1249), .A2(n1248), .ZN(n1243) );
XOR2_X1 U942 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U943 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U944 ( .A(KEYINPUT28), .B(n1254), .Z(n1253) );
NOR2_X1 U945 ( .A1(KEYINPUT18), .A2(n1173), .ZN(n1254) );
NAND2_X1 U946 ( .A1(G224), .A2(n1082), .ZN(n1173) );
XOR2_X1 U947 ( .A(n1170), .B(n1255), .Z(n1250) );
INV_X1 U948 ( .A(n1169), .ZN(n1255) );
XOR2_X1 U949 ( .A(n1256), .B(n1257), .Z(n1170) );
XOR2_X1 U950 ( .A(n1258), .B(n1259), .Z(n1256) );
INV_X1 U951 ( .A(n1260), .ZN(n1259) );
NAND2_X1 U952 ( .A1(KEYINPUT56), .A2(n1231), .ZN(n1258) );
XOR2_X1 U953 ( .A(n1190), .B(KEYINPUT49), .Z(n1237) );
NAND4_X1 U954 ( .A1(n1215), .A2(n1043), .A3(n1213), .A4(n1223), .ZN(n1190) );
NAND2_X1 U955 ( .A1(n1227), .A2(n1261), .ZN(n1223) );
NAND4_X1 U956 ( .A1(G953), .A2(G902), .A3(n1028), .A4(n1122), .ZN(n1261) );
INV_X1 U957 ( .A(G898), .ZN(n1122) );
NAND3_X1 U958 ( .A1(G952), .A2(n1028), .A3(n1262), .ZN(n1227) );
XOR2_X1 U959 ( .A(n1082), .B(KEYINPUT35), .Z(n1262) );
NAND2_X1 U960 ( .A1(G234), .A2(G237), .ZN(n1028) );
NOR2_X1 U961 ( .A1(n1263), .A2(n1064), .ZN(n1213) );
NOR2_X1 U962 ( .A1(n1070), .A2(G472), .ZN(n1064) );
AND2_X1 U963 ( .A1(n1264), .A2(n1070), .ZN(n1263) );
NAND2_X1 U964 ( .A1(n1265), .A2(n1248), .ZN(n1070) );
XOR2_X1 U965 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U966 ( .A(n1155), .B(n1154), .Z(n1267) );
XOR2_X1 U967 ( .A(n1268), .B(n1169), .Z(n1155) );
XOR2_X1 U968 ( .A(n1269), .B(n1270), .Z(n1169) );
XOR2_X1 U969 ( .A(n1271), .B(n1272), .Z(n1266) );
NOR2_X1 U970 ( .A1(KEYINPUT17), .A2(n1144), .ZN(n1272) );
XNOR2_X1 U971 ( .A(G116), .B(n1257), .ZN(n1144) );
XOR2_X1 U972 ( .A(G113), .B(G119), .Z(n1257) );
NAND2_X1 U973 ( .A1(n1273), .A2(KEYINPUT51), .ZN(n1271) );
XNOR2_X1 U974 ( .A(n1153), .B(KEYINPUT44), .ZN(n1273) );
AND2_X1 U975 ( .A1(G210), .A2(n1274), .ZN(n1153) );
XOR2_X1 U976 ( .A(KEYINPUT61), .B(G472), .Z(n1264) );
AND2_X1 U977 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U978 ( .A1(G221), .A2(n1275), .ZN(n1045) );
XNOR2_X1 U979 ( .A(n1276), .B(G469), .ZN(n1044) );
NAND2_X1 U980 ( .A1(n1277), .A2(n1248), .ZN(n1276) );
XOR2_X1 U981 ( .A(n1278), .B(n1160), .Z(n1277) );
XNOR2_X1 U982 ( .A(n1279), .B(n1280), .ZN(n1160) );
XOR2_X1 U983 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U984 ( .A(KEYINPUT53), .B(KEYINPUT41), .ZN(n1282) );
NAND2_X1 U985 ( .A1(G227), .A2(n1082), .ZN(n1281) );
XOR2_X1 U986 ( .A(n1260), .B(n1283), .Z(n1279) );
XOR2_X1 U987 ( .A(n1284), .B(n1268), .Z(n1283) );
XNOR2_X1 U988 ( .A(n1096), .B(n1285), .ZN(n1268) );
XOR2_X1 U989 ( .A(G137), .B(G134), .Z(n1285) );
INV_X1 U990 ( .A(G131), .ZN(n1096) );
INV_X1 U991 ( .A(n1091), .ZN(n1284) );
XOR2_X1 U992 ( .A(n1286), .B(n1287), .Z(n1091) );
NOR2_X1 U993 ( .A1(KEYINPUT37), .A2(n1288), .ZN(n1287) );
INV_X1 U994 ( .A(G143), .ZN(n1288) );
XOR2_X1 U995 ( .A(n1218), .B(G146), .Z(n1286) );
INV_X1 U996 ( .A(G128), .ZN(n1218) );
XOR2_X1 U997 ( .A(n1289), .B(n1290), .Z(n1260) );
XOR2_X1 U998 ( .A(G110), .B(G107), .Z(n1290) );
XNOR2_X1 U999 ( .A(G104), .B(n1154), .ZN(n1289) );
XOR2_X1 U1000 ( .A(G101), .B(KEYINPUT31), .Z(n1154) );
NOR2_X1 U1001 ( .A1(G140), .A2(KEYINPUT29), .ZN(n1278) );
NOR2_X1 U1002 ( .A1(n1041), .A2(n1051), .ZN(n1215) );
XNOR2_X1 U1003 ( .A(n1291), .B(n1127), .ZN(n1051) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1275), .ZN(n1127) );
NAND2_X1 U1005 ( .A1(G234), .A2(n1248), .ZN(n1275) );
OR2_X1 U1006 ( .A1(n1126), .A2(G902), .ZN(n1291) );
XNOR2_X1 U1007 ( .A(n1292), .B(n1293), .ZN(n1126) );
XOR2_X1 U1008 ( .A(G119), .B(n1294), .Z(n1293) );
XOR2_X1 U1009 ( .A(KEYINPUT9), .B(G128), .Z(n1294) );
XOR2_X1 U1010 ( .A(n1295), .B(n1296), .Z(n1292) );
XOR2_X1 U1011 ( .A(G110), .B(n1297), .Z(n1296) );
NOR2_X1 U1012 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR2_X1 U1013 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
INV_X1 U1014 ( .A(n1302), .ZN(n1301) );
NOR2_X1 U1015 ( .A1(KEYINPUT4), .A2(n1303), .ZN(n1300) );
NOR2_X1 U1016 ( .A1(G146), .A2(KEYINPUT6), .ZN(n1303) );
NOR2_X1 U1017 ( .A1(n1304), .A2(n1269), .ZN(n1298) );
INV_X1 U1018 ( .A(G146), .ZN(n1269) );
NOR2_X1 U1019 ( .A1(n1305), .A2(KEYINPUT6), .ZN(n1304) );
NOR2_X1 U1020 ( .A1(KEYINPUT4), .A2(n1302), .ZN(n1305) );
NAND3_X1 U1021 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1302) );
OR2_X1 U1022 ( .A1(n1225), .A2(KEYINPUT25), .ZN(n1308) );
NAND3_X1 U1023 ( .A1(KEYINPUT25), .A2(n1225), .A3(G140), .ZN(n1307) );
NAND2_X1 U1024 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
INV_X1 U1025 ( .A(G140), .ZN(n1310) );
NAND2_X1 U1026 ( .A1(n1311), .A2(KEYINPUT25), .ZN(n1309) );
XOR2_X1 U1027 ( .A(n1225), .B(KEYINPUT26), .Z(n1311) );
INV_X1 U1028 ( .A(G125), .ZN(n1225) );
NAND2_X1 U1029 ( .A1(n1312), .A2(n1313), .ZN(n1295) );
NAND2_X1 U1030 ( .A1(n1103), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1315), .ZN(n1314) );
INV_X1 U1032 ( .A(G137), .ZN(n1103) );
XOR2_X1 U1033 ( .A(KEYINPUT0), .B(n1316), .Z(n1312) );
NOR3_X1 U1034 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1316) );
INV_X1 U1035 ( .A(G221), .ZN(n1319) );
XOR2_X1 U1036 ( .A(KEYINPUT30), .B(G137), .Z(n1317) );
INV_X1 U1037 ( .A(n1222), .ZN(n1041) );
NOR2_X1 U1038 ( .A1(n1208), .A2(n1207), .ZN(n1222) );
XNOR2_X1 U1039 ( .A(n1074), .B(n1320), .ZN(n1207) );
XNOR2_X1 U1040 ( .A(n1321), .B(KEYINPUT59), .ZN(n1320) );
NAND2_X1 U1041 ( .A1(KEYINPUT19), .A2(n1073), .ZN(n1321) );
NAND2_X1 U1042 ( .A1(n1131), .A2(n1248), .ZN(n1073) );
XOR2_X1 U1043 ( .A(n1322), .B(n1323), .Z(n1131) );
AND2_X1 U1044 ( .A1(n1315), .A2(G217), .ZN(n1323) );
INV_X1 U1045 ( .A(n1318), .ZN(n1315) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1082), .ZN(n1318) );
NAND2_X1 U1047 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
OR2_X1 U1048 ( .A1(n1326), .A2(KEYINPUT38), .ZN(n1325) );
XOR2_X1 U1049 ( .A(n1327), .B(n1328), .Z(n1324) );
XOR2_X1 U1050 ( .A(n1329), .B(G107), .Z(n1328) );
NAND2_X1 U1051 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1052 ( .A1(G116), .A2(n1229), .ZN(n1331) );
INV_X1 U1053 ( .A(G122), .ZN(n1229) );
XOR2_X1 U1054 ( .A(n1332), .B(KEYINPUT12), .Z(n1330) );
NAND2_X1 U1055 ( .A1(G122), .A2(n1231), .ZN(n1332) );
INV_X1 U1056 ( .A(G116), .ZN(n1231) );
NAND2_X1 U1057 ( .A1(KEYINPUT38), .A2(n1326), .ZN(n1327) );
XOR2_X1 U1058 ( .A(G134), .B(n1270), .Z(n1326) );
XOR2_X1 U1059 ( .A(G128), .B(G143), .Z(n1270) );
XOR2_X1 U1060 ( .A(G478), .B(KEYINPUT39), .Z(n1074) );
NAND2_X1 U1061 ( .A1(n1333), .A2(n1334), .ZN(n1208) );
NAND2_X1 U1062 ( .A1(n1335), .A2(n1068), .ZN(n1334) );
XOR2_X1 U1063 ( .A(KEYINPUT2), .B(n1336), .Z(n1333) );
NOR2_X1 U1064 ( .A1(n1335), .A2(n1068), .ZN(n1336) );
NAND2_X1 U1065 ( .A1(n1337), .A2(n1248), .ZN(n1068) );
INV_X1 U1066 ( .A(G902), .ZN(n1248) );
XOR2_X1 U1067 ( .A(KEYINPUT32), .B(n1338), .Z(n1337) );
INV_X1 U1068 ( .A(n1135), .ZN(n1338) );
XOR2_X1 U1069 ( .A(n1339), .B(n1340), .Z(n1135) );
XOR2_X1 U1070 ( .A(n1252), .B(n1341), .Z(n1340) );
XNOR2_X1 U1071 ( .A(n1342), .B(n1343), .ZN(n1341) );
NOR2_X1 U1072 ( .A1(G104), .A2(KEYINPUT33), .ZN(n1343) );
NAND2_X1 U1073 ( .A1(KEYINPUT3), .A2(n1344), .ZN(n1342) );
INV_X1 U1074 ( .A(G113), .ZN(n1344) );
XOR2_X1 U1075 ( .A(G122), .B(G125), .Z(n1252) );
XOR2_X1 U1076 ( .A(n1345), .B(n1346), .Z(n1339) );
XOR2_X1 U1077 ( .A(G146), .B(G140), .Z(n1346) );
XOR2_X1 U1078 ( .A(n1347), .B(G131), .Z(n1345) );
NAND2_X1 U1079 ( .A1(KEYINPUT22), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1080 ( .A(G143), .B(n1349), .Z(n1348) );
AND2_X1 U1081 ( .A1(n1274), .A2(G214), .ZN(n1349) );
AND2_X1 U1082 ( .A1(n1350), .A2(n1082), .ZN(n1274) );
INV_X1 U1083 ( .A(G953), .ZN(n1082) );
XOR2_X1 U1084 ( .A(KEYINPUT1), .B(G237), .Z(n1350) );
INV_X1 U1085 ( .A(n1069), .ZN(n1335) );
XNOR2_X1 U1086 ( .A(G475), .B(KEYINPUT50), .ZN(n1069) );
endmodule


