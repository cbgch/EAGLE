//Key = 0110001110010100011000100011000111000001010100101001100011010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
n1444, n1445, n1446, n1447;

XNOR2_X1 U796 ( .A(n1114), .B(n1115), .ZN(G9) );
NAND2_X1 U797 ( .A1(KEYINPUT1), .A2(G107), .ZN(n1115) );
NAND4_X1 U798 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(G75) );
NAND2_X1 U799 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U800 ( .A1(KEYINPUT51), .A2(n1122), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND4_X1 U803 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
NAND2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NAND2_X1 U805 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
OR2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U807 ( .A1(n1137), .A2(n1138), .ZN(n1131) );
NAND2_X1 U808 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U809 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U810 ( .A(n1143), .B(KEYINPUT25), .ZN(n1141) );
INV_X1 U811 ( .A(n1144), .ZN(n1139) );
NAND3_X1 U812 ( .A1(n1133), .A2(n1145), .A3(n1137), .ZN(n1125) );
NAND2_X1 U813 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND3_X1 U814 ( .A1(n1148), .A2(n1149), .A3(n1127), .ZN(n1147) );
OR2_X1 U815 ( .A1(n1130), .A2(n1128), .ZN(n1149) );
OR3_X1 U816 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1148) );
NAND2_X1 U817 ( .A1(n1153), .A2(n1128), .ZN(n1146) );
NOR2_X1 U818 ( .A1(n1154), .A2(n1155), .ZN(n1118) );
NOR4_X1 U819 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
XOR2_X1 U820 ( .A(n1160), .B(KEYINPUT13), .Z(n1159) );
NAND2_X1 U821 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U822 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
INV_X1 U823 ( .A(n1163), .ZN(n1161) );
NAND3_X1 U824 ( .A1(n1130), .A2(n1164), .A3(n1165), .ZN(n1157) );
NAND4_X1 U825 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1156) );
NOR3_X1 U826 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
NOR3_X1 U827 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
INV_X1 U828 ( .A(KEYINPUT17), .ZN(n1173) );
NOR2_X1 U829 ( .A1(KEYINPUT17), .A2(G475), .ZN(n1171) );
XOR2_X1 U830 ( .A(n1176), .B(n1177), .Z(n1170) );
XNOR2_X1 U831 ( .A(n1178), .B(n1179), .ZN(n1168) );
XNOR2_X1 U832 ( .A(KEYINPUT43), .B(n1127), .ZN(n1167) );
NAND2_X1 U833 ( .A1(G952), .A2(n1180), .ZN(n1117) );
NAND2_X1 U834 ( .A1(KEYINPUT51), .A2(G953), .ZN(n1116) );
XOR2_X1 U835 ( .A(n1181), .B(n1182), .Z(G72) );
XOR2_X1 U836 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U837 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
AND2_X1 U838 ( .A1(G227), .A2(G900), .ZN(n1185) );
NAND2_X1 U839 ( .A1(n1187), .A2(n1188), .ZN(n1183) );
NAND2_X1 U840 ( .A1(G953), .A2(n1189), .ZN(n1188) );
XNOR2_X1 U841 ( .A(n1190), .B(n1191), .ZN(n1187) );
NAND3_X1 U842 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1190) );
NAND2_X1 U843 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
OR3_X1 U844 ( .A1(n1196), .A2(n1195), .A3(n1197), .ZN(n1193) );
INV_X1 U845 ( .A(KEYINPUT52), .ZN(n1197) );
NAND2_X1 U846 ( .A1(KEYINPUT18), .A2(n1198), .ZN(n1196) );
OR2_X1 U847 ( .A1(n1198), .A2(KEYINPUT52), .ZN(n1192) );
XOR2_X1 U848 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U849 ( .A(KEYINPUT7), .B(G131), .Z(n1200) );
XNOR2_X1 U850 ( .A(n1201), .B(n1202), .ZN(n1199) );
NOR2_X1 U851 ( .A1(KEYINPUT30), .A2(n1203), .ZN(n1202) );
NAND2_X1 U852 ( .A1(n1186), .A2(n1204), .ZN(n1181) );
NAND2_X1 U853 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U854 ( .A1(n1207), .A2(n1208), .ZN(G69) );
NAND2_X1 U855 ( .A1(n1209), .A2(n1186), .ZN(n1208) );
XOR2_X1 U856 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND2_X1 U857 ( .A1(n1212), .A2(G953), .ZN(n1207) );
NAND2_X1 U858 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U859 ( .A1(n1210), .A2(n1215), .ZN(n1214) );
INV_X1 U860 ( .A(G224), .ZN(n1215) );
NAND2_X1 U861 ( .A1(G224), .A2(n1216), .ZN(n1213) );
NAND2_X1 U862 ( .A1(G898), .A2(n1210), .ZN(n1216) );
NAND2_X1 U863 ( .A1(n1217), .A2(n1218), .ZN(n1210) );
NAND2_X1 U864 ( .A1(G953), .A2(n1219), .ZN(n1218) );
XOR2_X1 U865 ( .A(n1220), .B(n1221), .Z(n1217) );
XOR2_X1 U866 ( .A(n1222), .B(KEYINPUT50), .Z(n1220) );
NOR3_X1 U867 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(G66) );
AND3_X1 U868 ( .A1(KEYINPUT29), .A2(n1186), .A3(n1226), .ZN(n1225) );
NOR2_X1 U869 ( .A1(KEYINPUT29), .A2(n1227), .ZN(n1224) );
INV_X1 U870 ( .A(n1154), .ZN(n1227) );
XNOR2_X1 U871 ( .A(n1228), .B(n1229), .ZN(n1223) );
NOR2_X1 U872 ( .A1(n1177), .A2(n1230), .ZN(n1229) );
NOR2_X1 U873 ( .A1(n1231), .A2(n1232), .ZN(G63) );
XNOR2_X1 U874 ( .A(n1154), .B(KEYINPUT31), .ZN(n1232) );
XOR2_X1 U875 ( .A(n1233), .B(n1234), .Z(n1231) );
NOR3_X1 U876 ( .A1(n1179), .A2(n1235), .A3(n1236), .ZN(n1234) );
NOR2_X1 U877 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U878 ( .A1(n1239), .A2(n1180), .ZN(n1237) );
AND2_X1 U879 ( .A1(n1238), .A2(n1230), .ZN(n1235) );
INV_X1 U880 ( .A(KEYINPUT21), .ZN(n1238) );
INV_X1 U881 ( .A(G478), .ZN(n1179) );
NAND2_X1 U882 ( .A1(KEYINPUT8), .A2(n1240), .ZN(n1233) );
NOR2_X1 U883 ( .A1(n1154), .A2(n1241), .ZN(G60) );
XOR2_X1 U884 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U885 ( .A1(n1175), .A2(n1230), .ZN(n1242) );
XNOR2_X1 U886 ( .A(n1244), .B(n1245), .ZN(G6) );
NOR2_X1 U887 ( .A1(KEYINPUT0), .A2(n1246), .ZN(n1245) );
NOR2_X1 U888 ( .A1(n1154), .A2(n1247), .ZN(G57) );
XOR2_X1 U889 ( .A(n1248), .B(n1249), .Z(n1247) );
NOR2_X1 U890 ( .A1(KEYINPUT14), .A2(n1250), .ZN(n1248) );
XOR2_X1 U891 ( .A(n1251), .B(n1252), .Z(n1250) );
NOR2_X1 U892 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR2_X1 U893 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U894 ( .A(KEYINPUT24), .B(n1257), .Z(n1256) );
AND2_X1 U895 ( .A1(n1255), .A2(n1257), .ZN(n1253) );
XOR2_X1 U896 ( .A(n1258), .B(KEYINPUT62), .Z(n1257) );
AND2_X1 U897 ( .A1(n1259), .A2(n1260), .ZN(n1255) );
OR2_X1 U898 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U899 ( .A(KEYINPUT46), .B(n1263), .Z(n1259) );
NOR2_X1 U900 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U901 ( .A(n1262), .B(KEYINPUT2), .Z(n1265) );
NOR2_X1 U902 ( .A1(n1162), .A2(n1230), .ZN(n1251) );
INV_X1 U903 ( .A(G472), .ZN(n1162) );
NOR2_X1 U904 ( .A1(n1154), .A2(n1266), .ZN(G54) );
XOR2_X1 U905 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U906 ( .A(n1195), .B(n1269), .Z(n1268) );
XNOR2_X1 U907 ( .A(n1270), .B(n1262), .ZN(n1267) );
XOR2_X1 U908 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U909 ( .A1(n1273), .A2(n1230), .ZN(n1272) );
NAND2_X1 U910 ( .A1(KEYINPUT6), .A2(n1274), .ZN(n1271) );
NOR2_X1 U911 ( .A1(n1154), .A2(n1275), .ZN(G51) );
NOR2_X1 U912 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U913 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U914 ( .A1(KEYINPUT61), .A2(n1280), .ZN(n1279) );
NOR2_X1 U915 ( .A1(n1281), .A2(n1230), .ZN(n1278) );
NAND2_X1 U916 ( .A1(G902), .A2(n1180), .ZN(n1230) );
NAND3_X1 U917 ( .A1(n1211), .A2(n1205), .A3(n1282), .ZN(n1180) );
XOR2_X1 U918 ( .A(n1206), .B(KEYINPUT45), .Z(n1282) );
AND4_X1 U919 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1205) );
NOR4_X1 U920 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1286) );
NAND2_X1 U921 ( .A1(n1291), .A2(n1292), .ZN(n1285) );
XOR2_X1 U922 ( .A(KEYINPUT44), .B(n1135), .Z(n1292) );
AND4_X1 U923 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1211) );
NOR4_X1 U924 ( .A1(n1114), .A2(n1297), .A3(n1298), .A4(n1299), .ZN(n1296) );
AND3_X1 U925 ( .A1(n1136), .A2(n1128), .A3(n1300), .ZN(n1114) );
AND2_X1 U926 ( .A1(n1301), .A2(n1246), .ZN(n1295) );
NAND3_X1 U927 ( .A1(n1300), .A2(n1128), .A3(n1135), .ZN(n1246) );
AND2_X1 U928 ( .A1(n1280), .A2(KEYINPUT61), .ZN(n1276) );
XOR2_X1 U929 ( .A(n1264), .B(n1302), .Z(n1280) );
XOR2_X1 U930 ( .A(G125), .B(n1303), .Z(n1302) );
NOR2_X1 U931 ( .A1(n1186), .A2(G952), .ZN(n1154) );
INV_X1 U932 ( .A(G953), .ZN(n1186) );
XNOR2_X1 U933 ( .A(G146), .B(n1283), .ZN(G48) );
NAND3_X1 U934 ( .A1(n1135), .A2(n1304), .A3(n1305), .ZN(n1283) );
XNOR2_X1 U935 ( .A(G143), .B(n1206), .ZN(G45) );
NAND4_X1 U936 ( .A1(n1305), .A2(n1151), .A3(n1306), .A4(n1307), .ZN(n1206) );
XNOR2_X1 U937 ( .A(G140), .B(n1284), .ZN(G42) );
NAND3_X1 U938 ( .A1(n1135), .A2(n1150), .A3(n1308), .ZN(n1284) );
XOR2_X1 U939 ( .A(G137), .B(n1290), .Z(G39) );
AND3_X1 U940 ( .A1(n1304), .A2(n1137), .A3(n1308), .ZN(n1290) );
XOR2_X1 U941 ( .A(n1289), .B(n1309), .Z(G36) );
NOR2_X1 U942 ( .A1(KEYINPUT40), .A2(n1310), .ZN(n1309) );
INV_X1 U943 ( .A(G134), .ZN(n1310) );
AND3_X1 U944 ( .A1(n1136), .A2(n1151), .A3(n1308), .ZN(n1289) );
XOR2_X1 U945 ( .A(G131), .B(n1288), .Z(G33) );
AND3_X1 U946 ( .A1(n1135), .A2(n1151), .A3(n1308), .ZN(n1288) );
AND4_X1 U947 ( .A1(n1127), .A2(n1144), .A3(n1311), .A4(n1130), .ZN(n1308) );
XOR2_X1 U948 ( .A(G128), .B(n1287), .Z(G30) );
AND3_X1 U949 ( .A1(n1304), .A2(n1136), .A3(n1305), .ZN(n1287) );
AND3_X1 U950 ( .A1(n1144), .A2(n1311), .A3(n1153), .ZN(n1305) );
XNOR2_X1 U951 ( .A(G101), .B(n1301), .ZN(G3) );
NAND3_X1 U952 ( .A1(n1300), .A2(n1151), .A3(n1137), .ZN(n1301) );
NAND2_X1 U953 ( .A1(n1312), .A2(n1313), .ZN(G27) );
NAND4_X1 U954 ( .A1(n1291), .A2(n1135), .A3(n1314), .A4(n1315), .ZN(n1313) );
NAND2_X1 U955 ( .A1(G125), .A2(n1316), .ZN(n1315) );
OR2_X1 U956 ( .A1(n1317), .A2(G125), .ZN(n1314) );
NAND3_X1 U957 ( .A1(n1318), .A2(n1316), .A3(G125), .ZN(n1312) );
INV_X1 U958 ( .A(KEYINPUT54), .ZN(n1316) );
NAND3_X1 U959 ( .A1(n1135), .A2(n1317), .A3(n1291), .ZN(n1318) );
AND4_X1 U960 ( .A1(n1153), .A2(n1150), .A3(n1133), .A4(n1311), .ZN(n1291) );
NAND2_X1 U961 ( .A1(n1319), .A2(n1320), .ZN(n1311) );
NAND2_X1 U962 ( .A1(n1321), .A2(n1189), .ZN(n1319) );
INV_X1 U963 ( .A(G900), .ZN(n1189) );
INV_X1 U964 ( .A(KEYINPUT37), .ZN(n1317) );
XNOR2_X1 U965 ( .A(G122), .B(n1293), .ZN(G24) );
NAND4_X1 U966 ( .A1(n1306), .A2(n1322), .A3(n1128), .A4(n1307), .ZN(n1293) );
NAND2_X1 U967 ( .A1(n1323), .A2(n1324), .ZN(n1128) );
OR3_X1 U968 ( .A1(n1325), .A2(n1326), .A3(KEYINPUT58), .ZN(n1324) );
NAND2_X1 U969 ( .A1(KEYINPUT58), .A2(n1151), .ZN(n1323) );
XNOR2_X1 U970 ( .A(G119), .B(n1294), .ZN(G21) );
NAND3_X1 U971 ( .A1(n1304), .A2(n1137), .A3(n1322), .ZN(n1294) );
XOR2_X1 U972 ( .A(n1327), .B(G116), .Z(G18) );
NAND2_X1 U973 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U974 ( .A1(n1299), .A2(n1330), .ZN(n1329) );
INV_X1 U975 ( .A(KEYINPUT20), .ZN(n1330) );
AND3_X1 U976 ( .A1(n1136), .A2(n1151), .A3(n1322), .ZN(n1299) );
NAND3_X1 U977 ( .A1(n1153), .A2(n1331), .A3(KEYINPUT20), .ZN(n1328) );
NAND4_X1 U978 ( .A1(n1136), .A2(n1151), .A3(n1133), .A4(n1332), .ZN(n1331) );
NOR2_X1 U979 ( .A1(n1307), .A2(n1333), .ZN(n1136) );
XOR2_X1 U980 ( .A(G113), .B(n1298), .Z(G15) );
AND3_X1 U981 ( .A1(n1322), .A2(n1151), .A3(n1135), .ZN(n1298) );
AND2_X1 U982 ( .A1(n1333), .A2(n1307), .ZN(n1135) );
NOR2_X1 U983 ( .A1(n1325), .A2(n1334), .ZN(n1151) );
AND3_X1 U984 ( .A1(n1133), .A2(n1332), .A3(n1153), .ZN(n1322) );
NAND2_X1 U985 ( .A1(n1335), .A2(n1336), .ZN(n1133) );
OR3_X1 U986 ( .A1(n1143), .A2(n1142), .A3(KEYINPUT25), .ZN(n1336) );
NAND2_X1 U987 ( .A1(KEYINPUT25), .A2(n1144), .ZN(n1335) );
NAND3_X1 U988 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(G12) );
NAND2_X1 U989 ( .A1(n1297), .A2(n1340), .ZN(n1339) );
NAND2_X1 U990 ( .A1(n1341), .A2(n1342), .ZN(n1338) );
INV_X1 U991 ( .A(KEYINPUT32), .ZN(n1342) );
NAND2_X1 U992 ( .A1(n1343), .A2(G110), .ZN(n1341) );
XNOR2_X1 U993 ( .A(n1297), .B(KEYINPUT34), .ZN(n1343) );
NAND2_X1 U994 ( .A1(KEYINPUT32), .A2(n1344), .ZN(n1337) );
NAND2_X1 U995 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
OR3_X1 U996 ( .A1(n1340), .A2(n1297), .A3(KEYINPUT34), .ZN(n1346) );
NAND2_X1 U997 ( .A1(KEYINPUT34), .A2(n1297), .ZN(n1345) );
AND3_X1 U998 ( .A1(n1300), .A2(n1150), .A3(n1137), .ZN(n1297) );
NOR2_X1 U999 ( .A1(n1307), .A2(n1306), .ZN(n1137) );
INV_X1 U1000 ( .A(n1333), .ZN(n1306) );
XNOR2_X1 U1001 ( .A(n1178), .B(n1347), .ZN(n1333) );
NOR2_X1 U1002 ( .A1(G478), .A2(KEYINPUT15), .ZN(n1347) );
NAND2_X1 U1003 ( .A1(n1240), .A2(n1239), .ZN(n1178) );
XOR2_X1 U1004 ( .A(n1348), .B(n1349), .Z(n1240) );
XNOR2_X1 U1005 ( .A(n1201), .B(n1350), .ZN(n1349) );
XOR2_X1 U1006 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1007 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
INV_X1 U1008 ( .A(G217), .ZN(n1354) );
NAND2_X1 U1009 ( .A1(KEYINPUT11), .A2(n1355), .ZN(n1351) );
XOR2_X1 U1010 ( .A(n1356), .B(n1357), .Z(n1348) );
XOR2_X1 U1011 ( .A(G128), .B(G122), .Z(n1357) );
XNOR2_X1 U1012 ( .A(G107), .B(G116), .ZN(n1356) );
NAND2_X1 U1013 ( .A1(n1358), .A2(n1164), .ZN(n1307) );
NAND2_X1 U1014 ( .A1(n1174), .A2(n1175), .ZN(n1164) );
OR2_X1 U1015 ( .A1(n1175), .A2(n1174), .ZN(n1358) );
NOR2_X1 U1016 ( .A1(n1243), .A2(G902), .ZN(n1174) );
XNOR2_X1 U1017 ( .A(n1359), .B(n1360), .ZN(n1243) );
XOR2_X1 U1018 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1019 ( .A(n1244), .B(n1363), .ZN(n1362) );
NOR2_X1 U1020 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
INV_X1 U1021 ( .A(G214), .ZN(n1364) );
INV_X1 U1022 ( .A(G104), .ZN(n1244) );
XOR2_X1 U1023 ( .A(G122), .B(G113), .Z(n1361) );
XOR2_X1 U1024 ( .A(n1366), .B(n1367), .Z(n1359) );
XOR2_X1 U1025 ( .A(n1368), .B(n1191), .Z(n1367) );
NOR2_X1 U1026 ( .A1(G131), .A2(KEYINPUT42), .ZN(n1368) );
INV_X1 U1027 ( .A(G475), .ZN(n1175) );
NAND2_X1 U1028 ( .A1(n1369), .A2(n1370), .ZN(n1150) );
NAND3_X1 U1029 ( .A1(n1334), .A2(n1325), .A3(n1371), .ZN(n1370) );
INV_X1 U1030 ( .A(KEYINPUT58), .ZN(n1371) );
NAND2_X1 U1031 ( .A1(KEYINPUT58), .A2(n1304), .ZN(n1369) );
AND2_X1 U1032 ( .A1(n1326), .A2(n1325), .ZN(n1304) );
NAND2_X1 U1033 ( .A1(n1372), .A2(n1373), .ZN(n1325) );
NAND2_X1 U1034 ( .A1(n1374), .A2(KEYINPUT55), .ZN(n1373) );
XOR2_X1 U1035 ( .A(n1176), .B(n1375), .Z(n1372) );
NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n1374), .ZN(n1375) );
XOR2_X1 U1037 ( .A(n1177), .B(KEYINPUT28), .Z(n1374) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1376), .ZN(n1177) );
NAND2_X1 U1039 ( .A1(n1228), .A2(n1239), .ZN(n1176) );
XNOR2_X1 U1040 ( .A(n1377), .B(n1378), .ZN(n1228) );
XOR2_X1 U1041 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1042 ( .A(G128), .B(G119), .Z(n1380) );
XOR2_X1 U1043 ( .A(KEYINPUT19), .B(G146), .Z(n1379) );
XOR2_X1 U1044 ( .A(n1381), .B(n1382), .Z(n1377) );
XNOR2_X1 U1045 ( .A(n1340), .B(n1383), .ZN(n1382) );
NOR2_X1 U1046 ( .A1(n1384), .A2(n1353), .ZN(n1383) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1385), .ZN(n1353) );
INV_X1 U1048 ( .A(G221), .ZN(n1384) );
XNOR2_X1 U1049 ( .A(n1191), .B(n1203), .ZN(n1381) );
XOR2_X1 U1050 ( .A(G140), .B(G125), .Z(n1191) );
INV_X1 U1051 ( .A(n1334), .ZN(n1326) );
XNOR2_X1 U1052 ( .A(n1386), .B(n1387), .ZN(n1334) );
XNOR2_X1 U1053 ( .A(G472), .B(n1163), .ZN(n1387) );
NAND2_X1 U1054 ( .A1(n1388), .A2(n1239), .ZN(n1163) );
XNOR2_X1 U1055 ( .A(n1389), .B(n1249), .ZN(n1388) );
XOR2_X1 U1056 ( .A(G101), .B(n1390), .Z(n1249) );
NOR2_X1 U1057 ( .A1(n1391), .A2(n1365), .ZN(n1390) );
NAND2_X1 U1058 ( .A1(n1385), .A2(n1392), .ZN(n1365) );
INV_X1 U1059 ( .A(G210), .ZN(n1391) );
NAND2_X1 U1060 ( .A1(n1393), .A2(n1394), .ZN(n1389) );
NAND2_X1 U1061 ( .A1(n1258), .A2(n1395), .ZN(n1394) );
XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n1396), .Z(n1393) );
NOR2_X1 U1063 ( .A1(n1258), .A2(n1395), .ZN(n1396) );
XNOR2_X1 U1064 ( .A(n1397), .B(n1261), .ZN(n1395) );
XOR2_X1 U1065 ( .A(n1262), .B(KEYINPUT23), .Z(n1397) );
XNOR2_X1 U1066 ( .A(n1398), .B(n1399), .ZN(n1258) );
NOR2_X1 U1067 ( .A1(G119), .A2(KEYINPUT5), .ZN(n1399) );
XNOR2_X1 U1068 ( .A(KEYINPUT39), .B(KEYINPUT3), .ZN(n1386) );
AND3_X1 U1069 ( .A1(n1144), .A2(n1332), .A3(n1153), .ZN(n1300) );
NOR2_X1 U1070 ( .A1(n1127), .A2(n1152), .ZN(n1153) );
INV_X1 U1071 ( .A(n1130), .ZN(n1152) );
NAND2_X1 U1072 ( .A1(G214), .A2(n1400), .ZN(n1130) );
XNOR2_X1 U1073 ( .A(n1401), .B(n1281), .ZN(n1127) );
NAND2_X1 U1074 ( .A1(G210), .A2(n1400), .ZN(n1281) );
NAND2_X1 U1075 ( .A1(n1392), .A2(n1239), .ZN(n1400) );
INV_X1 U1076 ( .A(G237), .ZN(n1392) );
NAND2_X1 U1077 ( .A1(n1402), .A2(n1239), .ZN(n1401) );
XOR2_X1 U1078 ( .A(n1403), .B(n1303), .Z(n1402) );
XOR2_X1 U1079 ( .A(n1221), .B(n1404), .Z(n1303) );
XOR2_X1 U1080 ( .A(n1405), .B(n1406), .Z(n1404) );
AND2_X1 U1081 ( .A1(n1385), .A2(G224), .ZN(n1406) );
NOR3_X1 U1082 ( .A1(KEYINPUT60), .A2(n1407), .A3(n1408), .ZN(n1405) );
NOR2_X1 U1083 ( .A1(n1409), .A2(n1222), .ZN(n1408) );
NAND2_X1 U1084 ( .A1(n1410), .A2(n1411), .ZN(n1222) );
NAND2_X1 U1085 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
XNOR2_X1 U1086 ( .A(n1414), .B(n1415), .ZN(n1412) );
INV_X1 U1087 ( .A(G101), .ZN(n1414) );
INV_X1 U1088 ( .A(KEYINPUT48), .ZN(n1409) );
NOR2_X1 U1089 ( .A1(KEYINPUT48), .A2(n1410), .ZN(n1407) );
NAND2_X1 U1090 ( .A1(n1416), .A2(n1417), .ZN(n1410) );
INV_X1 U1091 ( .A(n1413), .ZN(n1417) );
XNOR2_X1 U1092 ( .A(n1398), .B(G119), .ZN(n1413) );
XNOR2_X1 U1093 ( .A(G113), .B(n1418), .ZN(n1398) );
XOR2_X1 U1094 ( .A(KEYINPUT4), .B(G116), .Z(n1418) );
XNOR2_X1 U1095 ( .A(G101), .B(n1415), .ZN(n1416) );
XNOR2_X1 U1096 ( .A(G122), .B(n1340), .ZN(n1221) );
INV_X1 U1097 ( .A(G110), .ZN(n1340) );
XOR2_X1 U1098 ( .A(n1419), .B(KEYINPUT38), .Z(n1403) );
NAND3_X1 U1099 ( .A1(n1420), .A2(n1421), .A3(n1422), .ZN(n1419) );
NAND2_X1 U1100 ( .A1(G125), .A2(n1423), .ZN(n1422) );
OR3_X1 U1101 ( .A1(n1423), .A2(G125), .A3(KEYINPUT16), .ZN(n1421) );
OR2_X1 U1102 ( .A1(KEYINPUT9), .A2(n1264), .ZN(n1423) );
NAND2_X1 U1103 ( .A1(KEYINPUT16), .A2(n1264), .ZN(n1420) );
INV_X1 U1104 ( .A(n1261), .ZN(n1264) );
NAND2_X1 U1105 ( .A1(n1424), .A2(n1425), .ZN(n1261) );
NAND2_X1 U1106 ( .A1(n1426), .A2(n1355), .ZN(n1425) );
INV_X1 U1107 ( .A(G143), .ZN(n1355) );
NAND2_X1 U1108 ( .A1(n1427), .A2(G143), .ZN(n1424) );
XNOR2_X1 U1109 ( .A(KEYINPUT12), .B(n1426), .ZN(n1427) );
XOR2_X1 U1110 ( .A(n1428), .B(G146), .Z(n1426) );
NAND2_X1 U1111 ( .A1(KEYINPUT22), .A2(G128), .ZN(n1428) );
NAND2_X1 U1112 ( .A1(n1429), .A2(n1320), .ZN(n1332) );
NAND2_X1 U1113 ( .A1(n1120), .A2(n1124), .ZN(n1320) );
NOR2_X1 U1114 ( .A1(n1226), .A2(G953), .ZN(n1120) );
INV_X1 U1115 ( .A(G952), .ZN(n1226) );
NAND2_X1 U1116 ( .A1(n1321), .A2(n1219), .ZN(n1429) );
INV_X1 U1117 ( .A(G898), .ZN(n1219) );
AND3_X1 U1118 ( .A1(G953), .A2(n1124), .A3(G902), .ZN(n1321) );
NAND2_X1 U1119 ( .A1(G237), .A2(n1430), .ZN(n1124) );
NOR2_X1 U1120 ( .A1(n1166), .A2(n1142), .ZN(n1144) );
INV_X1 U1121 ( .A(n1165), .ZN(n1142) );
NAND2_X1 U1122 ( .A1(G221), .A2(n1376), .ZN(n1165) );
NAND2_X1 U1123 ( .A1(n1430), .A2(n1239), .ZN(n1376) );
XNOR2_X1 U1124 ( .A(G234), .B(KEYINPUT27), .ZN(n1430) );
INV_X1 U1125 ( .A(n1143), .ZN(n1166) );
XOR2_X1 U1126 ( .A(n1431), .B(n1273), .Z(n1143) );
INV_X1 U1127 ( .A(G469), .ZN(n1273) );
NAND2_X1 U1128 ( .A1(n1432), .A2(n1239), .ZN(n1431) );
INV_X1 U1129 ( .A(G902), .ZN(n1239) );
XOR2_X1 U1130 ( .A(n1433), .B(n1434), .Z(n1432) );
XNOR2_X1 U1131 ( .A(n1435), .B(n1274), .ZN(n1434) );
XOR2_X1 U1132 ( .A(n1436), .B(n1437), .Z(n1274) );
XNOR2_X1 U1133 ( .A(n1438), .B(G110), .ZN(n1437) );
INV_X1 U1134 ( .A(G140), .ZN(n1438) );
NAND2_X1 U1135 ( .A1(G227), .A2(n1385), .ZN(n1436) );
XOR2_X1 U1136 ( .A(G953), .B(KEYINPUT26), .Z(n1385) );
XNOR2_X1 U1137 ( .A(n1195), .B(n1439), .ZN(n1435) );
NOR2_X1 U1138 ( .A1(KEYINPUT36), .A2(n1262), .ZN(n1439) );
XOR2_X1 U1139 ( .A(n1440), .B(n1203), .Z(n1262) );
XOR2_X1 U1140 ( .A(G137), .B(KEYINPUT10), .Z(n1203) );
XNOR2_X1 U1141 ( .A(G131), .B(n1201), .ZN(n1440) );
XOR2_X1 U1142 ( .A(G134), .B(KEYINPUT47), .Z(n1201) );
XNOR2_X1 U1143 ( .A(n1366), .B(n1441), .ZN(n1195) );
NOR2_X1 U1144 ( .A1(KEYINPUT35), .A2(n1442), .ZN(n1441) );
XOR2_X1 U1145 ( .A(KEYINPUT53), .B(G128), .Z(n1442) );
XNOR2_X1 U1146 ( .A(G143), .B(G146), .ZN(n1366) );
XOR2_X1 U1147 ( .A(n1443), .B(n1444), .Z(n1433) );
NOR2_X1 U1148 ( .A1(n1269), .A2(n1445), .ZN(n1444) );
XOR2_X1 U1149 ( .A(KEYINPUT63), .B(KEYINPUT59), .Z(n1445) );
XNOR2_X1 U1150 ( .A(n1415), .B(n1446), .ZN(n1269) );
NOR2_X1 U1151 ( .A1(KEYINPUT49), .A2(n1447), .ZN(n1446) );
XNOR2_X1 U1152 ( .A(G101), .B(KEYINPUT41), .ZN(n1447) );
XOR2_X1 U1153 ( .A(G104), .B(G107), .Z(n1415) );
XNOR2_X1 U1154 ( .A(KEYINPUT56), .B(KEYINPUT33), .ZN(n1443) );
endmodule


