//Key = 0111011001011010010001100011010011011010111000111101010111111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U746 ( .A(G107), .B(n1016), .ZN(G9) );
NAND2_X1 U747 ( .A1(KEYINPUT11), .A2(n1017), .ZN(n1016) );
INV_X1 U748 ( .A(n1018), .ZN(n1017) );
NOR2_X1 U749 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U750 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
NOR2_X1 U751 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR4_X1 U752 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1025) );
XOR2_X1 U753 ( .A(KEYINPUT10), .B(n1031), .Z(n1030) );
AND3_X1 U754 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
XOR2_X1 U755 ( .A(n1035), .B(KEYINPUT40), .Z(n1029) );
NAND4_X1 U756 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1034), .ZN(n1035) );
NOR2_X1 U757 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
XNOR2_X1 U758 ( .A(n1041), .B(KEYINPUT30), .ZN(n1039) );
INV_X1 U759 ( .A(n1042), .ZN(n1037) );
NOR2_X1 U760 ( .A1(KEYINPUT36), .A2(n1043), .ZN(n1028) );
AND2_X1 U761 ( .A1(n1032), .A2(n1044), .ZN(n1043) );
NOR3_X1 U762 ( .A1(n1042), .A2(n1045), .A3(n1046), .ZN(n1027) );
INV_X1 U763 ( .A(n1047), .ZN(n1046) );
NOR2_X1 U764 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
NOR2_X1 U765 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
INV_X1 U766 ( .A(n1034), .ZN(n1051) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U768 ( .A1(n1054), .A2(n1055), .ZN(n1048) );
NOR2_X1 U769 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
AND2_X1 U770 ( .A1(n1058), .A2(KEYINPUT36), .ZN(n1056) );
NAND4_X1 U771 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1021) );
NAND4_X1 U772 ( .A1(n1032), .A2(n1034), .A3(n1047), .A4(n1063), .ZN(n1059) );
NAND2_X1 U773 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U774 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U775 ( .A1(n1042), .A2(n1055), .ZN(n1032) );
NOR3_X1 U776 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1019) );
INV_X1 U777 ( .A(n1061), .ZN(n1068) );
NAND4_X1 U778 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1061) );
NOR4_X1 U779 ( .A1(n1073), .A2(n1074), .A3(n1066), .A4(n1036), .ZN(n1072) );
NOR2_X1 U780 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
AND2_X1 U781 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND3_X1 U782 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1073) );
NAND2_X1 U783 ( .A1(G478), .A2(n1082), .ZN(n1081) );
NAND2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
INV_X1 U785 ( .A(KEYINPUT38), .ZN(n1084) );
NAND2_X1 U786 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
OR2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(n1079) );
NOR4_X1 U788 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1071) );
AND3_X1 U789 ( .A1(KEYINPUT42), .A2(n1093), .A3(G475), .ZN(n1092) );
NOR2_X1 U790 ( .A1(KEYINPUT42), .A2(G475), .ZN(n1091) );
AND2_X1 U791 ( .A1(n1094), .A2(KEYINPUT15), .ZN(n1090) );
NOR3_X1 U792 ( .A1(KEYINPUT15), .A2(n1095), .A3(n1094), .ZN(n1089) );
XOR2_X1 U793 ( .A(n1096), .B(KEYINPUT0), .Z(n1070) );
NOR2_X1 U794 ( .A1(n1097), .A2(n1098), .ZN(n1069) );
NOR2_X1 U795 ( .A1(n1085), .A2(n1086), .ZN(n1098) );
INV_X1 U796 ( .A(n1099), .ZN(n1085) );
NOR2_X1 U797 ( .A1(G902), .A2(n1100), .ZN(n1097) );
NOR3_X1 U798 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NOR2_X1 U799 ( .A1(G478), .A2(n1104), .ZN(n1103) );
NOR2_X1 U800 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND3_X1 U801 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1101) );
NAND2_X1 U802 ( .A1(n1110), .A2(n1087), .ZN(n1109) );
NAND3_X1 U803 ( .A1(n1111), .A2(n1086), .A3(KEYINPUT38), .ZN(n1108) );
NAND2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U805 ( .A1(KEYINPUT42), .A2(G475), .ZN(n1113) );
NAND2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(G72) );
NAND2_X1 U807 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U808 ( .A(KEYINPUT58), .B(n1118), .Z(n1114) );
NOR2_X1 U809 ( .A1(n1116), .A2(n1119), .ZN(n1118) );
XOR2_X1 U810 ( .A(n1117), .B(n1024), .Z(n1119) );
OR2_X1 U811 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XNOR2_X1 U812 ( .A(n1122), .B(n1123), .ZN(n1120) );
XNOR2_X1 U813 ( .A(n1124), .B(n1125), .ZN(n1123) );
NOR2_X1 U814 ( .A1(KEYINPUT31), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U815 ( .A(n1127), .B(n1128), .ZN(n1126) );
XNOR2_X1 U816 ( .A(n1129), .B(n1130), .ZN(n1122) );
NAND2_X1 U817 ( .A1(KEYINPUT46), .A2(n1131), .ZN(n1129) );
AND2_X1 U818 ( .A1(G953), .A2(n1132), .ZN(n1116) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1132) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(G69) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U822 ( .A(n1137), .B(KEYINPUT27), .Z(n1136) );
NAND3_X1 U823 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
NAND2_X1 U824 ( .A1(G953), .A2(n1141), .ZN(n1139) );
NAND2_X1 U825 ( .A1(n1142), .A2(n1062), .ZN(n1138) );
NOR3_X1 U826 ( .A1(n1140), .A2(G953), .A3(n1143), .ZN(n1135) );
INV_X1 U827 ( .A(n1142), .ZN(n1143) );
NAND3_X1 U828 ( .A1(n1144), .A2(n1060), .A3(n1145), .ZN(n1142) );
XNOR2_X1 U829 ( .A(n1146), .B(n1147), .ZN(n1140) );
XNOR2_X1 U830 ( .A(n1148), .B(n1149), .ZN(n1146) );
NAND3_X1 U831 ( .A1(G953), .A2(n1150), .A3(KEYINPUT26), .ZN(n1133) );
NAND2_X1 U832 ( .A1(G898), .A2(G224), .ZN(n1150) );
NOR2_X1 U833 ( .A1(n1151), .A2(n1152), .ZN(G66) );
XNOR2_X1 U834 ( .A(n1153), .B(n1110), .ZN(n1152) );
NOR3_X1 U835 ( .A1(n1154), .A2(KEYINPUT43), .A3(n1087), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1151), .A2(n1155), .ZN(G63) );
XNOR2_X1 U837 ( .A(n1156), .B(n1104), .ZN(n1155) );
NAND2_X1 U838 ( .A1(n1157), .A2(G478), .ZN(n1156) );
NOR2_X1 U839 ( .A1(n1151), .A2(n1158), .ZN(G60) );
XOR2_X1 U840 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U841 ( .A1(G475), .A2(n1157), .ZN(n1160) );
NAND2_X1 U842 ( .A1(KEYINPUT33), .A2(n1112), .ZN(n1159) );
XNOR2_X1 U843 ( .A(G104), .B(n1161), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1151), .A2(n1162), .ZN(G57) );
XOR2_X1 U845 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U846 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U847 ( .A1(n1157), .A2(G472), .ZN(n1165) );
XOR2_X1 U848 ( .A(n1167), .B(KEYINPUT13), .Z(n1163) );
NAND2_X1 U849 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U850 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U851 ( .A(n1172), .B(KEYINPUT4), .Z(n1168) );
NAND2_X1 U852 ( .A1(n1130), .A2(n1173), .ZN(n1172) );
NOR2_X1 U853 ( .A1(n1151), .A2(n1174), .ZN(G54) );
XOR2_X1 U854 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U855 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U856 ( .A(G140), .B(n1179), .ZN(n1178) );
NAND2_X1 U857 ( .A1(n1157), .A2(G469), .ZN(n1177) );
XOR2_X1 U858 ( .A(n1180), .B(n1181), .Z(n1175) );
XNOR2_X1 U859 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND2_X1 U860 ( .A1(KEYINPUT9), .A2(n1184), .ZN(n1182) );
NOR2_X1 U861 ( .A1(n1151), .A2(n1185), .ZN(G51) );
XOR2_X1 U862 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U863 ( .A(n1188), .B(n1189), .ZN(n1187) );
XNOR2_X1 U864 ( .A(n1190), .B(n1130), .ZN(n1186) );
XOR2_X1 U865 ( .A(n1191), .B(KEYINPUT24), .Z(n1190) );
NAND2_X1 U866 ( .A1(n1157), .A2(n1105), .ZN(n1191) );
INV_X1 U867 ( .A(n1094), .ZN(n1105) );
INV_X1 U868 ( .A(n1154), .ZN(n1157) );
NAND2_X1 U869 ( .A1(n1192), .A2(n1193), .ZN(n1154) );
NAND3_X1 U870 ( .A1(n1194), .A2(n1060), .A3(n1195), .ZN(n1193) );
XOR2_X1 U871 ( .A(n1024), .B(KEYINPUT53), .Z(n1195) );
NAND2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1024) );
AND4_X1 U873 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
AND4_X1 U874 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1196) );
OR3_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
INV_X1 U877 ( .A(KEYINPUT39), .ZN(n1210) );
NOR3_X1 U878 ( .A1(n1026), .A2(n1033), .A3(n1211), .ZN(n1209) );
NOR2_X1 U879 ( .A1(KEYINPUT39), .A2(n1212), .ZN(n1207) );
NAND4_X1 U880 ( .A1(n1213), .A2(n1214), .A3(n1047), .A4(n1215), .ZN(n1060) );
INV_X1 U881 ( .A(n1216), .ZN(n1214) );
XOR2_X1 U882 ( .A(n1217), .B(KEYINPUT45), .Z(n1213) );
INV_X1 U883 ( .A(n1022), .ZN(n1194) );
NAND2_X1 U884 ( .A1(n1218), .A2(n1145), .ZN(n1022) );
AND3_X1 U885 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1145) );
NAND3_X1 U886 ( .A1(n1052), .A2(n1058), .A3(n1222), .ZN(n1221) );
XNOR2_X1 U887 ( .A(n1144), .B(KEYINPUT35), .ZN(n1218) );
AND4_X1 U888 ( .A1(n1161), .A2(n1223), .A3(n1224), .A4(n1018), .ZN(n1144) );
NAND3_X1 U889 ( .A1(n1058), .A2(n1041), .A3(n1225), .ZN(n1018) );
NAND3_X1 U890 ( .A1(n1225), .A2(n1041), .A3(n1057), .ZN(n1161) );
XNOR2_X1 U891 ( .A(KEYINPUT44), .B(n1077), .ZN(n1192) );
NOR2_X1 U892 ( .A1(n1062), .A2(G952), .ZN(n1151) );
XNOR2_X1 U893 ( .A(G146), .B(n1203), .ZN(G48) );
NAND4_X1 U894 ( .A1(n1226), .A2(n1227), .A3(n1057), .A4(n1228), .ZN(n1203) );
XOR2_X1 U895 ( .A(n1202), .B(n1229), .Z(G45) );
NAND2_X1 U896 ( .A1(KEYINPUT41), .A2(G143), .ZN(n1229) );
NAND4_X1 U897 ( .A1(n1227), .A2(n1052), .A3(n1230), .A4(n1231), .ZN(n1202) );
XOR2_X1 U898 ( .A(n1201), .B(n1232), .Z(G42) );
XNOR2_X1 U899 ( .A(G140), .B(KEYINPUT25), .ZN(n1232) );
NAND3_X1 U900 ( .A1(n1053), .A2(n1057), .A3(n1212), .ZN(n1201) );
XOR2_X1 U901 ( .A(n1233), .B(n1234), .Z(G39) );
NAND2_X1 U902 ( .A1(n1212), .A2(n1235), .ZN(n1234) );
NAND2_X1 U903 ( .A1(KEYINPUT14), .A2(n1236), .ZN(n1233) );
XOR2_X1 U904 ( .A(KEYINPUT19), .B(G137), .Z(n1236) );
XNOR2_X1 U905 ( .A(G134), .B(n1200), .ZN(G36) );
NAND3_X1 U906 ( .A1(n1052), .A2(n1058), .A3(n1212), .ZN(n1200) );
XNOR2_X1 U907 ( .A(G131), .B(n1199), .ZN(G33) );
NAND3_X1 U908 ( .A1(n1057), .A2(n1052), .A3(n1212), .ZN(n1199) );
NOR3_X1 U909 ( .A1(n1237), .A2(n1211), .A3(n1026), .ZN(n1212) );
NAND2_X1 U910 ( .A1(n1067), .A2(n1238), .ZN(n1026) );
XNOR2_X1 U911 ( .A(G128), .B(n1198), .ZN(G30) );
NAND4_X1 U912 ( .A1(n1226), .A2(n1227), .A3(n1058), .A4(n1228), .ZN(n1198) );
NOR3_X1 U913 ( .A1(n1237), .A2(n1211), .A3(n1064), .ZN(n1227) );
XNOR2_X1 U914 ( .A(G101), .B(n1223), .ZN(G3) );
NAND3_X1 U915 ( .A1(n1052), .A2(n1225), .A3(n1034), .ZN(n1223) );
XNOR2_X1 U916 ( .A(G125), .B(n1204), .ZN(G27) );
NAND4_X1 U917 ( .A1(n1053), .A2(n1057), .A3(n1239), .A4(n1047), .ZN(n1204) );
NOR2_X1 U918 ( .A1(n1211), .A2(n1064), .ZN(n1239) );
INV_X1 U919 ( .A(n1215), .ZN(n1064) );
AND2_X1 U920 ( .A1(n1042), .A2(n1240), .ZN(n1211) );
NAND3_X1 U921 ( .A1(G902), .A2(n1241), .A3(n1121), .ZN(n1240) );
NOR2_X1 U922 ( .A1(n1062), .A2(G900), .ZN(n1121) );
XNOR2_X1 U923 ( .A(n1242), .B(n1243), .ZN(G24) );
NOR2_X1 U924 ( .A1(n1244), .A2(n1216), .ZN(n1243) );
NAND3_X1 U925 ( .A1(n1230), .A2(n1231), .A3(n1041), .ZN(n1216) );
INV_X1 U926 ( .A(n1055), .ZN(n1041) );
NAND2_X1 U927 ( .A1(n1245), .A2(n1246), .ZN(n1055) );
INV_X1 U928 ( .A(n1228), .ZN(n1246) );
XOR2_X1 U929 ( .A(n1219), .B(n1247), .Z(G21) );
NAND2_X1 U930 ( .A1(KEYINPUT22), .A2(G119), .ZN(n1247) );
NAND2_X1 U931 ( .A1(n1235), .A2(n1222), .ZN(n1219) );
INV_X1 U932 ( .A(n1206), .ZN(n1235) );
NAND3_X1 U933 ( .A1(n1226), .A2(n1228), .A3(n1034), .ZN(n1206) );
XNOR2_X1 U934 ( .A(G116), .B(n1248), .ZN(G18) );
NAND4_X1 U935 ( .A1(n1249), .A2(n1044), .A3(n1052), .A4(n1217), .ZN(n1248) );
AND2_X1 U936 ( .A1(n1047), .A2(n1058), .ZN(n1044) );
NOR2_X1 U937 ( .A1(n1231), .A2(n1250), .ZN(n1058) );
XNOR2_X1 U938 ( .A(n1215), .B(KEYINPUT48), .ZN(n1249) );
XOR2_X1 U939 ( .A(n1220), .B(n1251), .Z(G15) );
XOR2_X1 U940 ( .A(KEYINPUT12), .B(G113), .Z(n1251) );
NAND3_X1 U941 ( .A1(n1222), .A2(n1052), .A3(n1057), .ZN(n1220) );
AND2_X1 U942 ( .A1(n1250), .A2(n1231), .ZN(n1057) );
AND2_X1 U943 ( .A1(n1245), .A2(n1228), .ZN(n1052) );
XNOR2_X1 U944 ( .A(KEYINPUT5), .B(n1252), .ZN(n1245) );
INV_X1 U945 ( .A(n1244), .ZN(n1222) );
NAND3_X1 U946 ( .A1(n1215), .A2(n1217), .A3(n1047), .ZN(n1244) );
NOR2_X1 U947 ( .A1(n1040), .A2(n1036), .ZN(n1047) );
INV_X1 U948 ( .A(n1253), .ZN(n1036) );
NAND2_X1 U949 ( .A1(n1254), .A2(n1255), .ZN(G12) );
NAND2_X1 U950 ( .A1(G110), .A2(n1224), .ZN(n1255) );
XOR2_X1 U951 ( .A(n1256), .B(KEYINPUT54), .Z(n1254) );
OR2_X1 U952 ( .A1(n1224), .A2(G110), .ZN(n1256) );
NAND3_X1 U953 ( .A1(n1034), .A2(n1225), .A3(n1053), .ZN(n1224) );
AND2_X1 U954 ( .A1(n1257), .A2(n1226), .ZN(n1053) );
XNOR2_X1 U955 ( .A(n1252), .B(KEYINPUT28), .ZN(n1226) );
XNOR2_X1 U956 ( .A(n1087), .B(n1258), .ZN(n1252) );
NOR2_X1 U957 ( .A1(n1088), .A2(KEYINPUT52), .ZN(n1258) );
AND2_X1 U958 ( .A1(n1110), .A2(n1077), .ZN(n1088) );
XOR2_X1 U959 ( .A(n1259), .B(n1260), .Z(n1110) );
XNOR2_X1 U960 ( .A(n1261), .B(n1262), .ZN(n1260) );
NOR2_X1 U961 ( .A1(KEYINPUT37), .A2(n1263), .ZN(n1262) );
XOR2_X1 U962 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U963 ( .A(G110), .B(n1266), .ZN(n1265) );
NAND2_X1 U964 ( .A1(n1267), .A2(KEYINPUT51), .ZN(n1266) );
XNOR2_X1 U965 ( .A(G125), .B(n1268), .ZN(n1267) );
XNOR2_X1 U966 ( .A(KEYINPUT2), .B(n1124), .ZN(n1268) );
XNOR2_X1 U967 ( .A(G119), .B(n1269), .ZN(n1264) );
XOR2_X1 U968 ( .A(G146), .B(G128), .Z(n1269) );
NAND4_X1 U969 ( .A1(n1270), .A2(KEYINPUT1), .A3(G221), .A4(G234), .ZN(n1261) );
XNOR2_X1 U970 ( .A(G953), .B(KEYINPUT61), .ZN(n1270) );
XNOR2_X1 U971 ( .A(G137), .B(KEYINPUT62), .ZN(n1259) );
NAND2_X1 U972 ( .A1(G217), .A2(n1271), .ZN(n1087) );
XNOR2_X1 U973 ( .A(n1228), .B(KEYINPUT16), .ZN(n1257) );
XNOR2_X1 U974 ( .A(n1272), .B(n1273), .ZN(n1228) );
XNOR2_X1 U975 ( .A(KEYINPUT6), .B(n1086), .ZN(n1273) );
INV_X1 U976 ( .A(G472), .ZN(n1086) );
NAND2_X1 U977 ( .A1(KEYINPUT49), .A2(n1099), .ZN(n1272) );
NAND2_X1 U978 ( .A1(n1111), .A2(n1077), .ZN(n1099) );
XOR2_X1 U979 ( .A(n1166), .B(n1183), .Z(n1111) );
XOR2_X1 U980 ( .A(n1173), .B(n1171), .Z(n1183) );
XNOR2_X1 U981 ( .A(n1148), .B(n1274), .ZN(n1166) );
XNOR2_X1 U982 ( .A(G101), .B(n1275), .ZN(n1274) );
NAND2_X1 U983 ( .A1(n1276), .A2(G210), .ZN(n1275) );
AND3_X1 U984 ( .A1(n1033), .A2(n1217), .A3(n1215), .ZN(n1225) );
NOR2_X1 U985 ( .A1(n1067), .A2(n1066), .ZN(n1215) );
INV_X1 U986 ( .A(n1238), .ZN(n1066) );
NAND2_X1 U987 ( .A1(G214), .A2(n1277), .ZN(n1238) );
XOR2_X1 U988 ( .A(n1095), .B(n1094), .Z(n1067) );
NAND2_X1 U989 ( .A1(G210), .A2(n1277), .ZN(n1094) );
NAND2_X1 U990 ( .A1(n1278), .A2(n1077), .ZN(n1277) );
XOR2_X1 U991 ( .A(KEYINPUT63), .B(G237), .Z(n1278) );
NOR2_X1 U992 ( .A1(n1106), .A2(G902), .ZN(n1095) );
XOR2_X1 U993 ( .A(n1279), .B(n1189), .Z(n1106) );
XNOR2_X1 U994 ( .A(n1131), .B(n1280), .ZN(n1189) );
AND2_X1 U995 ( .A1(n1062), .A2(G224), .ZN(n1280) );
XNOR2_X1 U996 ( .A(n1281), .B(n1282), .ZN(n1279) );
NOR2_X1 U997 ( .A1(KEYINPUT23), .A2(n1130), .ZN(n1282) );
NOR2_X1 U998 ( .A1(KEYINPUT18), .A2(n1188), .ZN(n1281) );
XNOR2_X1 U999 ( .A(n1283), .B(n1149), .ZN(n1188) );
XNOR2_X1 U1000 ( .A(n1284), .B(G122), .ZN(n1149) );
NAND2_X1 U1001 ( .A1(KEYINPUT47), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1002 ( .A(KEYINPUT57), .B(n1184), .ZN(n1285) );
INV_X1 U1003 ( .A(G110), .ZN(n1184) );
NAND3_X1 U1004 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1283) );
NAND2_X1 U1005 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
INV_X1 U1006 ( .A(n1148), .ZN(n1290) );
INV_X1 U1007 ( .A(n1147), .ZN(n1289) );
NAND2_X1 U1008 ( .A1(n1291), .A2(n1292), .ZN(n1287) );
INV_X1 U1009 ( .A(KEYINPUT60), .ZN(n1292) );
NAND2_X1 U1010 ( .A1(n1293), .A2(n1148), .ZN(n1291) );
XNOR2_X1 U1011 ( .A(KEYINPUT56), .B(n1147), .ZN(n1293) );
NAND2_X1 U1012 ( .A1(KEYINPUT60), .A2(n1294), .ZN(n1286) );
NAND2_X1 U1013 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
OR2_X1 U1014 ( .A1(n1147), .A2(KEYINPUT56), .ZN(n1296) );
NAND3_X1 U1015 ( .A1(n1148), .A2(n1147), .A3(KEYINPUT56), .ZN(n1295) );
XOR2_X1 U1016 ( .A(n1297), .B(n1298), .Z(n1147) );
NAND2_X1 U1017 ( .A1(KEYINPUT29), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1018 ( .A(n1300), .B(G104), .ZN(n1299) );
INV_X1 U1019 ( .A(G107), .ZN(n1300) );
XOR2_X1 U1020 ( .A(G113), .B(n1301), .Z(n1148) );
XNOR2_X1 U1021 ( .A(G119), .B(n1302), .ZN(n1301) );
NAND2_X1 U1022 ( .A1(n1042), .A2(n1303), .ZN(n1217) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1141), .ZN(n1303) );
INV_X1 U1024 ( .A(G898), .ZN(n1141) );
NAND3_X1 U1025 ( .A1(n1241), .A2(n1062), .A3(G952), .ZN(n1042) );
NAND2_X1 U1026 ( .A1(G234), .A2(G237), .ZN(n1241) );
INV_X1 U1027 ( .A(n1237), .ZN(n1033) );
NAND2_X1 U1028 ( .A1(n1253), .A2(n1040), .ZN(n1237) );
NAND2_X1 U1029 ( .A1(n1304), .A2(n1096), .ZN(n1040) );
NAND3_X1 U1030 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1096) );
INV_X1 U1031 ( .A(G469), .ZN(n1076) );
NAND2_X1 U1032 ( .A1(G469), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1033 ( .A1(n1078), .A2(n1077), .ZN(n1305) );
XOR2_X1 U1034 ( .A(n1306), .B(n1307), .Z(n1078) );
XOR2_X1 U1035 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1036 ( .A(G110), .B(n1179), .ZN(n1309) );
AND2_X1 U1037 ( .A1(G227), .A2(n1062), .ZN(n1179) );
NAND2_X1 U1038 ( .A1(KEYINPUT55), .A2(n1124), .ZN(n1308) );
XNOR2_X1 U1039 ( .A(n1310), .B(n1170), .ZN(n1306) );
INV_X1 U1040 ( .A(n1173), .ZN(n1170) );
XNOR2_X1 U1041 ( .A(n1311), .B(n1128), .ZN(n1173) );
XOR2_X1 U1042 ( .A(G131), .B(G137), .Z(n1128) );
NAND2_X1 U1043 ( .A1(KEYINPUT3), .A2(n1127), .ZN(n1311) );
NAND2_X1 U1044 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
NAND2_X1 U1045 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
INV_X1 U1046 ( .A(KEYINPUT50), .ZN(n1315) );
XNOR2_X1 U1047 ( .A(n1171), .B(n1180), .ZN(n1314) );
NAND3_X1 U1048 ( .A1(n1180), .A2(n1130), .A3(KEYINPUT50), .ZN(n1312) );
INV_X1 U1049 ( .A(n1171), .ZN(n1130) );
XOR2_X1 U1050 ( .A(G146), .B(n1316), .Z(n1171) );
XNOR2_X1 U1051 ( .A(n1317), .B(n1298), .ZN(n1180) );
INV_X1 U1052 ( .A(G101), .ZN(n1298) );
NAND2_X1 U1053 ( .A1(n1318), .A2(KEYINPUT32), .ZN(n1317) );
XNOR2_X1 U1054 ( .A(G107), .B(n1319), .ZN(n1318) );
NOR2_X1 U1055 ( .A1(G104), .A2(KEYINPUT34), .ZN(n1319) );
NAND2_X1 U1056 ( .A1(G221), .A2(n1271), .ZN(n1253) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1077), .ZN(n1271) );
NOR2_X1 U1058 ( .A1(n1231), .A2(n1230), .ZN(n1034) );
INV_X1 U1059 ( .A(n1250), .ZN(n1230) );
XNOR2_X1 U1060 ( .A(n1320), .B(G478), .ZN(n1250) );
NAND2_X1 U1061 ( .A1(KEYINPUT59), .A2(n1082), .ZN(n1320) );
NAND2_X1 U1062 ( .A1(n1321), .A2(n1077), .ZN(n1082) );
INV_X1 U1063 ( .A(n1104), .ZN(n1321) );
XNOR2_X1 U1064 ( .A(n1322), .B(n1323), .ZN(n1104) );
XNOR2_X1 U1065 ( .A(n1324), .B(n1316), .ZN(n1323) );
XOR2_X1 U1066 ( .A(G128), .B(G143), .Z(n1316) );
NAND2_X1 U1067 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1068 ( .A1(G122), .A2(n1302), .ZN(n1326) );
INV_X1 U1069 ( .A(G116), .ZN(n1302) );
XOR2_X1 U1070 ( .A(n1327), .B(KEYINPUT20), .Z(n1325) );
NAND2_X1 U1071 ( .A1(G116), .A2(n1242), .ZN(n1327) );
XOR2_X1 U1072 ( .A(n1328), .B(n1329), .Z(n1322) );
XNOR2_X1 U1073 ( .A(n1127), .B(G107), .ZN(n1329) );
INV_X1 U1074 ( .A(G134), .ZN(n1127) );
NAND3_X1 U1075 ( .A1(G234), .A2(n1062), .A3(G217), .ZN(n1328) );
INV_X1 U1076 ( .A(G953), .ZN(n1062) );
XNOR2_X1 U1077 ( .A(n1093), .B(n1330), .ZN(n1231) );
XOR2_X1 U1078 ( .A(KEYINPUT8), .B(G475), .Z(n1330) );
NAND2_X1 U1079 ( .A1(n1112), .A2(n1077), .ZN(n1093) );
INV_X1 U1080 ( .A(G902), .ZN(n1077) );
XNOR2_X1 U1081 ( .A(n1331), .B(n1332), .ZN(n1112) );
XNOR2_X1 U1082 ( .A(G104), .B(n1333), .ZN(n1332) );
NAND2_X1 U1083 ( .A1(n1276), .A2(G214), .ZN(n1333) );
NOR2_X1 U1084 ( .A1(G953), .A2(G237), .ZN(n1276) );
XOR2_X1 U1085 ( .A(n1334), .B(n1335), .Z(n1331) );
XOR2_X1 U1086 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1087 ( .A(G143), .B(n1124), .ZN(n1337) );
INV_X1 U1088 ( .A(G140), .ZN(n1124) );
XOR2_X1 U1089 ( .A(KEYINPUT7), .B(G146), .Z(n1336) );
XOR2_X1 U1090 ( .A(n1338), .B(n1339), .Z(n1334) );
XOR2_X1 U1091 ( .A(G131), .B(G113), .Z(n1339) );
XNOR2_X1 U1092 ( .A(n1340), .B(n1341), .ZN(n1338) );
NAND2_X1 U1093 ( .A1(KEYINPUT21), .A2(n1131), .ZN(n1341) );
INV_X1 U1094 ( .A(G125), .ZN(n1131) );
NAND2_X1 U1095 ( .A1(KEYINPUT17), .A2(n1242), .ZN(n1340) );
INV_X1 U1096 ( .A(G122), .ZN(n1242) );
endmodule


