//Key = 0100010001101011011000110100001100010000000111110111100111010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385;

XNOR2_X1 U760 ( .A(G107), .B(n1040), .ZN(G9) );
NAND2_X1 U761 ( .A1(KEYINPUT51), .A2(n1041), .ZN(n1040) );
INV_X1 U762 ( .A(n1042), .ZN(n1041) );
NOR2_X1 U763 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR3_X1 U764 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NAND3_X1 U765 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1045) );
NAND2_X1 U766 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
NAND2_X1 U767 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND4_X1 U768 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND2_X1 U769 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XNOR2_X1 U770 ( .A(n1061), .B(KEYINPUT13), .ZN(n1059) );
NAND2_X1 U771 ( .A1(n1062), .A2(n1063), .ZN(n1053) );
NAND2_X1 U772 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U773 ( .A1(n1057), .A2(n1066), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U775 ( .A1(n1055), .A2(n1069), .ZN(n1068) );
NAND2_X1 U776 ( .A1(n1056), .A2(n1070), .ZN(n1064) );
NAND2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U778 ( .A1(n1057), .A2(n1073), .ZN(n1072) );
NAND2_X1 U779 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U780 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U781 ( .A(KEYINPUT24), .B(n1078), .Z(n1077) );
NAND2_X1 U782 ( .A1(n1055), .A2(n1079), .ZN(n1071) );
NAND2_X1 U783 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U784 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U785 ( .A(n1084), .ZN(n1051) );
AND3_X1 U786 ( .A1(n1050), .A2(n1085), .A3(n1049), .ZN(n1043) );
NAND4_X1 U787 ( .A1(n1056), .A2(n1057), .A3(n1086), .A4(n1087), .ZN(n1049) );
NOR3_X1 U788 ( .A1(n1088), .A2(n1078), .A3(n1089), .ZN(n1087) );
XOR2_X1 U789 ( .A(n1090), .B(G472), .Z(n1086) );
INV_X1 U790 ( .A(G952), .ZN(n1085) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(G72) );
NAND2_X1 U792 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U793 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
NAND2_X1 U794 ( .A1(n1097), .A2(n1094), .ZN(n1096) );
NAND2_X1 U795 ( .A1(G953), .A2(n1098), .ZN(n1094) );
INV_X1 U796 ( .A(n1093), .ZN(n1095) );
XNOR2_X1 U797 ( .A(n1099), .B(n1100), .ZN(n1093) );
NOR2_X1 U798 ( .A1(n1101), .A2(G953), .ZN(n1100) );
NAND2_X1 U799 ( .A1(n1102), .A2(n1097), .ZN(n1099) );
INV_X1 U800 ( .A(n1103), .ZN(n1097) );
XOR2_X1 U801 ( .A(n1104), .B(n1105), .Z(n1102) );
XNOR2_X1 U802 ( .A(n1106), .B(KEYINPUT35), .ZN(n1105) );
NAND2_X1 U803 ( .A1(KEYINPUT46), .A2(n1107), .ZN(n1106) );
NAND2_X1 U804 ( .A1(n1108), .A2(n1109), .ZN(G69) );
NAND2_X1 U805 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1112), .B(KEYINPUT11), .Z(n1108) );
NAND2_X1 U807 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U808 ( .A(n1111), .B(n1115), .ZN(n1114) );
NOR3_X1 U809 ( .A1(n1116), .A2(KEYINPUT41), .A3(G953), .ZN(n1115) );
NAND2_X1 U810 ( .A1(n1117), .A2(n1118), .ZN(n1111) );
XNOR2_X1 U811 ( .A(n1119), .B(n1120), .ZN(n1117) );
XNOR2_X1 U812 ( .A(KEYINPUT34), .B(n1110), .ZN(n1113) );
NAND2_X1 U813 ( .A1(n1118), .A2(n1121), .ZN(n1110) );
NAND2_X1 U814 ( .A1(G953), .A2(n1122), .ZN(n1121) );
INV_X1 U815 ( .A(n1123), .ZN(n1118) );
NOR2_X1 U816 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U817 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U818 ( .A(KEYINPUT43), .B(n1128), .Z(n1127) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U820 ( .A1(n1124), .A2(n1131), .ZN(G63) );
XOR2_X1 U821 ( .A(n1132), .B(n1133), .Z(n1131) );
AND2_X1 U822 ( .A1(G478), .A2(n1134), .ZN(n1132) );
NOR2_X1 U823 ( .A1(n1124), .A2(n1135), .ZN(G60) );
XOR2_X1 U824 ( .A(n1136), .B(n1137), .Z(n1135) );
AND2_X1 U825 ( .A1(G475), .A2(n1134), .ZN(n1137) );
XNOR2_X1 U826 ( .A(G104), .B(n1138), .ZN(G6) );
NAND4_X1 U827 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1062), .ZN(n1138) );
NOR2_X1 U828 ( .A1(KEYINPUT61), .A2(n1142), .ZN(n1141) );
NOR2_X1 U829 ( .A1(n1124), .A2(n1143), .ZN(G57) );
XOR2_X1 U830 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U831 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1144) );
AND2_X1 U833 ( .A1(G472), .A2(n1134), .ZN(n1149) );
NOR2_X1 U834 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
XOR2_X1 U835 ( .A(n1152), .B(KEYINPUT62), .Z(n1151) );
NAND2_X1 U836 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U837 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NOR2_X1 U838 ( .A1(n1124), .A2(n1155), .ZN(G54) );
XOR2_X1 U839 ( .A(n1156), .B(n1157), .Z(n1155) );
AND2_X1 U840 ( .A1(G469), .A2(n1134), .ZN(n1157) );
INV_X1 U841 ( .A(n1130), .ZN(n1134) );
NOR3_X1 U842 ( .A1(n1158), .A2(KEYINPUT36), .A3(n1159), .ZN(n1156) );
NOR2_X1 U843 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U844 ( .A(n1162), .B(KEYINPUT44), .Z(n1158) );
NAND2_X1 U845 ( .A1(n1160), .A2(n1161), .ZN(n1162) );
XNOR2_X1 U846 ( .A(n1163), .B(n1164), .ZN(n1161) );
XNOR2_X1 U847 ( .A(n1165), .B(n1166), .ZN(n1160) );
XOR2_X1 U848 ( .A(n1153), .B(n1167), .Z(n1165) );
NOR2_X1 U849 ( .A1(KEYINPUT58), .A2(n1168), .ZN(n1167) );
NOR2_X1 U850 ( .A1(n1124), .A2(n1169), .ZN(G51) );
NOR2_X1 U851 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U852 ( .A(n1172), .B(KEYINPUT45), .Z(n1171) );
NAND2_X1 U853 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
OR3_X1 U854 ( .A1(n1175), .A2(KEYINPUT21), .A3(n1130), .ZN(n1174) );
NOR4_X1 U855 ( .A1(KEYINPUT21), .A2(n1173), .A3(n1175), .A4(n1130), .ZN(n1170) );
NAND2_X1 U856 ( .A1(G902), .A2(n1176), .ZN(n1130) );
NAND2_X1 U857 ( .A1(n1116), .A2(n1101), .ZN(n1176) );
INV_X1 U858 ( .A(n1046), .ZN(n1101) );
NAND4_X1 U859 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1046) );
NOR3_X1 U860 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NOR3_X1 U861 ( .A1(n1080), .A2(n1184), .A3(n1185), .ZN(n1183) );
NOR2_X1 U862 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR3_X1 U863 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
INV_X1 U864 ( .A(n1069), .ZN(n1190) );
NOR4_X1 U865 ( .A1(n1142), .A2(n1139), .A3(n1191), .A4(n1074), .ZN(n1186) );
NOR2_X1 U866 ( .A1(n1192), .A2(n1193), .ZN(n1181) );
NOR2_X1 U867 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
INV_X1 U868 ( .A(n1047), .ZN(n1116) );
NAND4_X1 U869 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1047) );
AND4_X1 U870 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1042), .ZN(n1199) );
NAND3_X1 U871 ( .A1(n1069), .A2(n1062), .A3(n1140), .ZN(n1042) );
NOR2_X1 U872 ( .A1(n1203), .A2(n1204), .ZN(n1198) );
NOR2_X1 U873 ( .A1(n1080), .A2(n1205), .ZN(n1204) );
NOR2_X1 U874 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
NAND4_X1 U875 ( .A1(n1062), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1197) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND4_X1 U877 ( .A1(n1055), .A2(n1213), .A3(n1080), .A4(n1207), .ZN(n1212) );
INV_X1 U878 ( .A(KEYINPUT23), .ZN(n1207) );
OR2_X1 U879 ( .A1(n1211), .A2(n1140), .ZN(n1209) );
NAND3_X1 U880 ( .A1(n1061), .A2(n1214), .A3(n1215), .ZN(n1196) );
INV_X1 U881 ( .A(G210), .ZN(n1175) );
XNOR2_X1 U882 ( .A(n1216), .B(G125), .ZN(n1173) );
NOR2_X1 U883 ( .A1(n1217), .A2(G952), .ZN(n1124) );
XNOR2_X1 U884 ( .A(G146), .B(n1178), .ZN(G48) );
NAND3_X1 U885 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1178) );
XOR2_X1 U886 ( .A(n1221), .B(n1222), .Z(G45) );
NOR2_X1 U887 ( .A1(KEYINPUT20), .A2(n1223), .ZN(n1222) );
NOR4_X1 U888 ( .A1(n1224), .A2(n1080), .A3(n1142), .A4(n1139), .ZN(n1221) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U890 ( .A(n1061), .B(KEYINPUT47), .ZN(n1225) );
XNOR2_X1 U891 ( .A(G140), .B(n1227), .ZN(G42) );
NAND2_X1 U892 ( .A1(n1228), .A2(n1057), .ZN(n1227) );
XNOR2_X1 U893 ( .A(n1195), .B(KEYINPUT9), .ZN(n1228) );
AND2_X1 U894 ( .A1(n1220), .A2(n1229), .ZN(n1195) );
XNOR2_X1 U895 ( .A(n1182), .B(n1230), .ZN(G39) );
XNOR2_X1 U896 ( .A(G137), .B(KEYINPUT16), .ZN(n1230) );
AND4_X1 U897 ( .A1(n1226), .A2(n1218), .A3(n1056), .A4(n1057), .ZN(n1182) );
XNOR2_X1 U898 ( .A(n1231), .B(n1179), .ZN(G36) );
NAND4_X1 U899 ( .A1(n1226), .A2(n1061), .A3(n1057), .A4(n1069), .ZN(n1179) );
NAND2_X1 U900 ( .A1(KEYINPUT57), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U901 ( .A(n1233), .B(n1234), .ZN(G33) );
NOR2_X1 U902 ( .A1(n1193), .A2(n1235), .ZN(n1234) );
XOR2_X1 U903 ( .A(KEYINPUT55), .B(n1194), .Z(n1235) );
AND2_X1 U904 ( .A1(n1220), .A2(n1061), .ZN(n1194) );
AND3_X1 U905 ( .A1(n1139), .A2(n1208), .A3(n1226), .ZN(n1220) );
NOR2_X1 U906 ( .A1(n1074), .A2(n1184), .ZN(n1226) );
XNOR2_X1 U907 ( .A(n1189), .B(KEYINPUT56), .ZN(n1074) );
INV_X1 U908 ( .A(n1057), .ZN(n1193) );
NOR2_X1 U909 ( .A1(n1236), .A2(n1082), .ZN(n1057) );
XNOR2_X1 U910 ( .A(G128), .B(n1237), .ZN(G30) );
NAND4_X1 U911 ( .A1(n1218), .A2(n1069), .A3(KEYINPUT15), .A4(n1238), .ZN(n1237) );
NOR3_X1 U912 ( .A1(n1189), .A2(n1184), .A3(n1080), .ZN(n1238) );
INV_X1 U913 ( .A(n1219), .ZN(n1080) );
INV_X1 U914 ( .A(n1239), .ZN(n1184) );
XNOR2_X1 U915 ( .A(n1240), .B(n1241), .ZN(G3) );
NAND2_X1 U916 ( .A1(KEYINPUT5), .A2(n1202), .ZN(n1240) );
NAND3_X1 U917 ( .A1(n1056), .A2(n1140), .A3(n1061), .ZN(n1202) );
XNOR2_X1 U918 ( .A(G125), .B(n1177), .ZN(G27) );
NAND4_X1 U919 ( .A1(n1215), .A2(n1229), .A3(n1219), .A4(n1239), .ZN(n1177) );
NAND2_X1 U920 ( .A1(n1084), .A2(n1242), .ZN(n1239) );
NAND3_X1 U921 ( .A1(G902), .A2(n1243), .A3(n1103), .ZN(n1242) );
NOR2_X1 U922 ( .A1(G900), .A2(n1217), .ZN(n1103) );
XNOR2_X1 U923 ( .A(G122), .B(n1206), .ZN(G24) );
NAND3_X1 U924 ( .A1(n1055), .A2(n1062), .A3(n1244), .ZN(n1206) );
NOR3_X1 U925 ( .A1(n1245), .A2(n1142), .A3(n1139), .ZN(n1244) );
INV_X1 U926 ( .A(n1208), .ZN(n1142) );
NOR2_X1 U927 ( .A1(n1246), .A2(n1247), .ZN(n1062) );
XNOR2_X1 U928 ( .A(G119), .B(n1248), .ZN(G21) );
NAND2_X1 U929 ( .A1(n1249), .A2(n1219), .ZN(n1248) );
XOR2_X1 U930 ( .A(n1205), .B(KEYINPUT25), .Z(n1249) );
NAND4_X1 U931 ( .A1(n1218), .A2(n1055), .A3(n1056), .A4(n1213), .ZN(n1205) );
INV_X1 U932 ( .A(n1188), .ZN(n1218) );
NAND2_X1 U933 ( .A1(n1247), .A2(n1246), .ZN(n1188) );
XNOR2_X1 U934 ( .A(G116), .B(n1201), .ZN(G18) );
NAND4_X1 U935 ( .A1(n1061), .A2(n1055), .A3(n1069), .A4(n1214), .ZN(n1201) );
NOR2_X1 U936 ( .A1(n1208), .A2(n1139), .ZN(n1069) );
NAND2_X1 U937 ( .A1(n1250), .A2(n1251), .ZN(G15) );
NAND2_X1 U938 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U939 ( .A1(n1254), .A2(n1255), .ZN(n1252) );
NAND2_X1 U940 ( .A1(KEYINPUT32), .A2(n1256), .ZN(n1255) );
OR2_X1 U941 ( .A1(n1257), .A2(KEYINPUT32), .ZN(n1254) );
NAND2_X1 U942 ( .A1(G113), .A2(n1257), .ZN(n1250) );
NOR2_X1 U943 ( .A1(n1258), .A2(KEYINPUT54), .ZN(n1257) );
INV_X1 U944 ( .A(n1256), .ZN(n1258) );
NAND3_X1 U945 ( .A1(n1214), .A2(n1259), .A3(n1215), .ZN(n1256) );
INV_X1 U946 ( .A(n1067), .ZN(n1215) );
NAND3_X1 U947 ( .A1(n1139), .A2(n1208), .A3(n1055), .ZN(n1067) );
AND2_X1 U948 ( .A1(n1076), .A2(n1260), .ZN(n1055) );
INV_X1 U949 ( .A(n1088), .ZN(n1076) );
INV_X1 U950 ( .A(n1211), .ZN(n1139) );
XNOR2_X1 U951 ( .A(KEYINPUT7), .B(n1191), .ZN(n1259) );
INV_X1 U952 ( .A(n1061), .ZN(n1191) );
NOR2_X1 U953 ( .A1(n1247), .A2(n1261), .ZN(n1061) );
INV_X1 U954 ( .A(n1245), .ZN(n1214) );
XNOR2_X1 U955 ( .A(G110), .B(n1200), .ZN(G12) );
NAND3_X1 U956 ( .A1(n1056), .A2(n1140), .A3(n1229), .ZN(n1200) );
INV_X1 U957 ( .A(n1060), .ZN(n1229) );
NAND2_X1 U958 ( .A1(n1261), .A2(n1247), .ZN(n1060) );
XOR2_X1 U959 ( .A(n1089), .B(KEYINPUT42), .Z(n1247) );
XNOR2_X1 U960 ( .A(n1129), .B(n1262), .ZN(n1089) );
AND2_X1 U961 ( .A1(n1263), .A2(n1126), .ZN(n1262) );
XNOR2_X1 U962 ( .A(n1264), .B(n1265), .ZN(n1126) );
XOR2_X1 U963 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U964 ( .A1(KEYINPUT3), .A2(n1104), .ZN(n1266) );
XOR2_X1 U965 ( .A(n1268), .B(n1269), .Z(n1264) );
NOR2_X1 U966 ( .A1(KEYINPUT33), .A2(n1270), .ZN(n1269) );
XOR2_X1 U967 ( .A(n1271), .B(G137), .Z(n1270) );
NAND3_X1 U968 ( .A1(n1272), .A2(n1217), .A3(G221), .ZN(n1271) );
XOR2_X1 U969 ( .A(KEYINPUT48), .B(G234), .Z(n1272) );
XNOR2_X1 U970 ( .A(G119), .B(G110), .ZN(n1268) );
NAND2_X1 U971 ( .A1(G217), .A2(n1273), .ZN(n1129) );
INV_X1 U972 ( .A(n1246), .ZN(n1261) );
NAND2_X1 U973 ( .A1(n1274), .A2(n1275), .ZN(n1246) );
OR2_X1 U974 ( .A1(n1090), .A2(G472), .ZN(n1275) );
XOR2_X1 U975 ( .A(n1276), .B(KEYINPUT19), .Z(n1274) );
NAND2_X1 U976 ( .A1(G472), .A2(n1090), .ZN(n1276) );
NAND3_X1 U977 ( .A1(n1277), .A2(n1278), .A3(n1263), .ZN(n1090) );
NAND2_X1 U978 ( .A1(KEYINPUT12), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U979 ( .A(n1280), .B(n1281), .ZN(n1279) );
NAND2_X1 U980 ( .A1(n1282), .A2(n1283), .ZN(n1277) );
INV_X1 U981 ( .A(KEYINPUT12), .ZN(n1283) );
NAND2_X1 U982 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND2_X1 U983 ( .A1(n1281), .A2(n1286), .ZN(n1285) );
INV_X1 U984 ( .A(n1280), .ZN(n1286) );
NOR2_X1 U985 ( .A1(n1287), .A2(KEYINPUT29), .ZN(n1281) );
NAND3_X1 U986 ( .A1(KEYINPUT29), .A2(n1147), .A3(n1280), .ZN(n1284) );
XNOR2_X1 U987 ( .A(n1288), .B(KEYINPUT49), .ZN(n1280) );
NAND2_X1 U988 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U989 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U990 ( .A(n1293), .B(n1154), .ZN(n1292) );
XNOR2_X1 U991 ( .A(KEYINPUT6), .B(n1146), .ZN(n1291) );
XOR2_X1 U992 ( .A(n1294), .B(KEYINPUT8), .Z(n1289) );
NAND2_X1 U993 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U994 ( .A(n1154), .B(n1293), .Z(n1296) );
NOR2_X1 U995 ( .A1(KEYINPUT60), .A2(n1153), .ZN(n1293) );
XNOR2_X1 U996 ( .A(n1297), .B(KEYINPUT26), .ZN(n1154) );
XOR2_X1 U997 ( .A(KEYINPUT6), .B(n1146), .Z(n1295) );
XNOR2_X1 U998 ( .A(n1298), .B(G113), .ZN(n1146) );
NAND2_X1 U999 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U1000 ( .A1(G116), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1001 ( .A(n1302), .B(KEYINPUT28), .Z(n1299) );
OR2_X1 U1002 ( .A1(n1301), .A2(G116), .ZN(n1302) );
INV_X1 U1003 ( .A(n1287), .ZN(n1147) );
XOR2_X1 U1004 ( .A(n1303), .B(n1241), .Z(n1287) );
NAND3_X1 U1005 ( .A1(n1304), .A2(n1217), .A3(G210), .ZN(n1303) );
NOR2_X1 U1006 ( .A1(n1245), .A2(n1189), .ZN(n1140) );
NAND2_X1 U1007 ( .A1(n1260), .A2(n1088), .ZN(n1189) );
XNOR2_X1 U1008 ( .A(n1305), .B(G469), .ZN(n1088) );
NAND2_X1 U1009 ( .A1(n1306), .A2(n1263), .ZN(n1305) );
XOR2_X1 U1010 ( .A(n1307), .B(KEYINPUT0), .Z(n1306) );
NAND2_X1 U1011 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
OR2_X1 U1012 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1013 ( .A(n1312), .B(KEYINPUT53), .Z(n1308) );
NAND2_X1 U1014 ( .A1(n1311), .A2(n1310), .ZN(n1312) );
NAND2_X1 U1015 ( .A1(n1313), .A2(n1314), .ZN(n1310) );
NAND2_X1 U1016 ( .A1(n1164), .A2(G110), .ZN(n1314) );
NAND2_X1 U1017 ( .A1(n1315), .A2(n1163), .ZN(n1313) );
INV_X1 U1018 ( .A(G110), .ZN(n1163) );
XNOR2_X1 U1019 ( .A(n1164), .B(KEYINPUT2), .ZN(n1315) );
XOR2_X1 U1020 ( .A(G140), .B(n1316), .Z(n1164) );
NOR2_X1 U1021 ( .A1(G953), .A2(n1098), .ZN(n1316) );
INV_X1 U1022 ( .A(G227), .ZN(n1098) );
XOR2_X1 U1023 ( .A(n1166), .B(n1107), .Z(n1311) );
XNOR2_X1 U1024 ( .A(n1168), .B(n1153), .ZN(n1107) );
XNOR2_X1 U1025 ( .A(G131), .B(n1317), .ZN(n1153) );
XNOR2_X1 U1026 ( .A(G137), .B(n1232), .ZN(n1317) );
INV_X1 U1027 ( .A(G134), .ZN(n1232) );
XNOR2_X1 U1028 ( .A(G143), .B(n1267), .ZN(n1168) );
XNOR2_X1 U1029 ( .A(n1318), .B(G146), .ZN(n1267) );
INV_X1 U1030 ( .A(G128), .ZN(n1318) );
NAND2_X1 U1031 ( .A1(n1319), .A2(n1320), .ZN(n1166) );
NAND2_X1 U1032 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
INV_X1 U1033 ( .A(n1323), .ZN(n1322) );
NAND2_X1 U1034 ( .A1(n1324), .A2(n1325), .ZN(n1321) );
NAND2_X1 U1035 ( .A1(G107), .A2(n1241), .ZN(n1325) );
NAND2_X1 U1036 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
NAND2_X1 U1037 ( .A1(n1323), .A2(n1328), .ZN(n1319) );
NAND2_X1 U1038 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1039 ( .A1(n1241), .A2(n1327), .ZN(n1330) );
NAND2_X1 U1040 ( .A1(n1326), .A2(G107), .ZN(n1329) );
XNOR2_X1 U1041 ( .A(n1331), .B(G101), .ZN(n1326) );
XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(KEYINPUT1), .ZN(n1331) );
NOR2_X1 U1043 ( .A1(n1332), .A2(G104), .ZN(n1323) );
INV_X1 U1044 ( .A(KEYINPUT10), .ZN(n1332) );
XOR2_X1 U1045 ( .A(KEYINPUT14), .B(n1078), .Z(n1260) );
AND2_X1 U1046 ( .A1(G221), .A2(n1273), .ZN(n1078) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1263), .ZN(n1273) );
NAND2_X1 U1048 ( .A1(n1219), .A2(n1213), .ZN(n1245) );
NAND2_X1 U1049 ( .A1(n1084), .A2(n1333), .ZN(n1213) );
NAND3_X1 U1050 ( .A1(n1123), .A2(n1243), .A3(G902), .ZN(n1333) );
NOR2_X1 U1051 ( .A1(G898), .A2(n1217), .ZN(n1123) );
NAND3_X1 U1052 ( .A1(n1050), .A2(n1243), .A3(G952), .ZN(n1084) );
NAND2_X1 U1053 ( .A1(G234), .A2(G237), .ZN(n1243) );
XOR2_X1 U1054 ( .A(G953), .B(KEYINPUT18), .Z(n1050) );
NOR2_X1 U1055 ( .A1(n1083), .A2(n1082), .ZN(n1219) );
AND2_X1 U1056 ( .A1(G214), .A2(n1334), .ZN(n1082) );
NAND2_X1 U1057 ( .A1(n1263), .A2(n1304), .ZN(n1334) );
INV_X1 U1058 ( .A(n1236), .ZN(n1083) );
NAND2_X1 U1059 ( .A1(n1335), .A2(n1336), .ZN(n1236) );
NAND2_X1 U1060 ( .A1(G210), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1061 ( .A1(n1263), .A2(n1338), .ZN(n1337) );
OR2_X1 U1062 ( .A1(n1304), .A2(n1339), .ZN(n1338) );
NAND3_X1 U1063 ( .A1(n1340), .A2(n1263), .A3(n1339), .ZN(n1335) );
XOR2_X1 U1064 ( .A(n1216), .B(n1341), .Z(n1339) );
NOR2_X1 U1065 ( .A1(G125), .A2(KEYINPUT38), .ZN(n1341) );
XOR2_X1 U1066 ( .A(n1342), .B(n1343), .Z(n1216) );
XOR2_X1 U1067 ( .A(n1344), .B(n1345), .Z(n1343) );
NOR2_X1 U1068 ( .A1(KEYINPUT39), .A2(n1120), .ZN(n1345) );
NAND2_X1 U1069 ( .A1(n1346), .A2(n1347), .ZN(n1120) );
NAND2_X1 U1070 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XNOR2_X1 U1071 ( .A(G110), .B(KEYINPUT22), .ZN(n1348) );
XOR2_X1 U1072 ( .A(n1350), .B(KEYINPUT63), .Z(n1346) );
NAND2_X1 U1073 ( .A1(n1351), .A2(G122), .ZN(n1350) );
XNOR2_X1 U1074 ( .A(G110), .B(KEYINPUT27), .ZN(n1351) );
NOR2_X1 U1075 ( .A1(G953), .A2(n1122), .ZN(n1344) );
INV_X1 U1076 ( .A(G224), .ZN(n1122) );
XOR2_X1 U1077 ( .A(n1119), .B(n1297), .Z(n1342) );
XOR2_X1 U1078 ( .A(G128), .B(n1352), .Z(n1297) );
NOR2_X1 U1079 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NOR3_X1 U1080 ( .A1(KEYINPUT31), .A2(G146), .A3(n1223), .ZN(n1354) );
NOR2_X1 U1081 ( .A1(n1355), .A2(n1356), .ZN(n1353) );
INV_X1 U1082 ( .A(KEYINPUT31), .ZN(n1356) );
XNOR2_X1 U1083 ( .A(G146), .B(n1223), .ZN(n1355) );
XOR2_X1 U1084 ( .A(n1357), .B(n1358), .Z(n1119) );
XOR2_X1 U1085 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1086 ( .A(G104), .B(n1241), .ZN(n1360) );
INV_X1 U1087 ( .A(G101), .ZN(n1241) );
XNOR2_X1 U1088 ( .A(G113), .B(n1361), .ZN(n1357) );
XNOR2_X1 U1089 ( .A(KEYINPUT17), .B(n1301), .ZN(n1361) );
INV_X1 U1090 ( .A(G119), .ZN(n1301) );
INV_X1 U1091 ( .A(G902), .ZN(n1263) );
NAND2_X1 U1092 ( .A1(G210), .A2(G237), .ZN(n1340) );
NOR2_X1 U1093 ( .A1(n1211), .A2(n1208), .ZN(n1056) );
XOR2_X1 U1094 ( .A(G475), .B(n1362), .Z(n1208) );
NOR2_X1 U1095 ( .A1(n1136), .A2(G902), .ZN(n1362) );
AND2_X1 U1096 ( .A1(n1363), .A2(n1364), .ZN(n1136) );
NAND2_X1 U1097 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1098 ( .A(KEYINPUT59), .B(n1367), .Z(n1363) );
NOR2_X1 U1099 ( .A1(n1365), .A2(n1366), .ZN(n1367) );
XNOR2_X1 U1100 ( .A(n1368), .B(n1369), .ZN(n1366) );
XNOR2_X1 U1101 ( .A(n1349), .B(G104), .ZN(n1369) );
INV_X1 U1102 ( .A(G122), .ZN(n1349) );
NAND2_X1 U1103 ( .A1(KEYINPUT30), .A2(n1253), .ZN(n1368) );
INV_X1 U1104 ( .A(G113), .ZN(n1253) );
XNOR2_X1 U1105 ( .A(n1370), .B(n1371), .ZN(n1365) );
XNOR2_X1 U1106 ( .A(G146), .B(n1233), .ZN(n1371) );
INV_X1 U1107 ( .A(G131), .ZN(n1233) );
XNOR2_X1 U1108 ( .A(n1372), .B(n1104), .ZN(n1370) );
XNOR2_X1 U1109 ( .A(G140), .B(G125), .ZN(n1104) );
NAND2_X1 U1110 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND4_X1 U1111 ( .A1(G214), .A2(n1375), .A3(n1304), .A4(n1217), .ZN(n1374) );
NAND2_X1 U1112 ( .A1(n1376), .A2(n1377), .ZN(n1373) );
NAND3_X1 U1113 ( .A1(n1304), .A2(n1217), .A3(G214), .ZN(n1377) );
INV_X1 U1114 ( .A(G237), .ZN(n1304) );
XOR2_X1 U1115 ( .A(KEYINPUT50), .B(n1375), .Z(n1376) );
XNOR2_X1 U1116 ( .A(n1223), .B(KEYINPUT4), .ZN(n1375) );
XNOR2_X1 U1117 ( .A(n1378), .B(G478), .ZN(n1211) );
OR2_X1 U1118 ( .A1(n1133), .A2(G902), .ZN(n1378) );
XNOR2_X1 U1119 ( .A(n1379), .B(n1380), .ZN(n1133) );
XOR2_X1 U1120 ( .A(n1359), .B(n1381), .Z(n1380) );
XOR2_X1 U1121 ( .A(n1382), .B(n1383), .Z(n1381) );
NOR2_X1 U1122 ( .A1(G122), .A2(KEYINPUT37), .ZN(n1383) );
AND3_X1 U1123 ( .A1(G217), .A2(n1217), .A3(G234), .ZN(n1382) );
INV_X1 U1124 ( .A(G953), .ZN(n1217) );
XNOR2_X1 U1125 ( .A(G116), .B(n1327), .ZN(n1359) );
INV_X1 U1126 ( .A(G107), .ZN(n1327) );
XOR2_X1 U1127 ( .A(n1384), .B(n1385), .Z(n1379) );
NOR2_X1 U1128 ( .A1(KEYINPUT40), .A2(n1223), .ZN(n1385) );
INV_X1 U1129 ( .A(G143), .ZN(n1223) );
XNOR2_X1 U1130 ( .A(G134), .B(G128), .ZN(n1384) );
endmodule


