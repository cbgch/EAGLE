//Key = 0111100100100010111101100000111111110010001010011100101110110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314;

XNOR2_X1 U721 ( .A(n1005), .B(n1006), .ZN(G9) );
NOR3_X1 U722 ( .A1(n1007), .A2(KEYINPUT53), .A3(n1008), .ZN(n1006) );
NAND3_X1 U723 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(G75) );
NAND2_X1 U724 ( .A1(G952), .A2(n1012), .ZN(n1011) );
NAND4_X1 U725 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR2_X1 U726 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U727 ( .A1(KEYINPUT6), .A2(n1019), .ZN(n1015) );
NAND4_X1 U728 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1014) );
NAND2_X1 U729 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND3_X1 U730 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
INV_X1 U731 ( .A(KEYINPUT3), .ZN(n1027) );
NAND2_X1 U732 ( .A1(n1029), .A2(n1030), .ZN(n1022) );
NAND3_X1 U733 ( .A1(n1031), .A2(n1032), .A3(KEYINPUT46), .ZN(n1029) );
NAND2_X1 U734 ( .A1(n1024), .A2(n1033), .ZN(n1013) );
NAND2_X1 U735 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U736 ( .A1(n1036), .A2(n1037), .A3(n1031), .ZN(n1035) );
NAND2_X1 U737 ( .A1(n1020), .A2(n1038), .ZN(n1036) );
NAND2_X1 U738 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U739 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
OR2_X1 U740 ( .A1(n1007), .A2(KEYINPUT45), .ZN(n1042) );
NAND2_X1 U741 ( .A1(n1021), .A2(n1043), .ZN(n1034) );
NAND2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U743 ( .A1(n1039), .A2(n1046), .A3(n1020), .ZN(n1045) );
NAND2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U746 ( .A1(n1031), .A2(n1051), .ZN(n1044) );
NAND2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U748 ( .A1(n1054), .A2(n1037), .ZN(n1053) );
NAND2_X1 U749 ( .A1(n1055), .A2(n1056), .ZN(n1037) );
NAND3_X1 U750 ( .A1(n1057), .A2(n1039), .A3(KEYINPUT45), .ZN(n1055) );
NAND2_X1 U751 ( .A1(n1058), .A2(n1059), .ZN(n1054) );
NAND2_X1 U752 ( .A1(n1032), .A2(n1060), .ZN(n1059) );
INV_X1 U753 ( .A(KEYINPUT46), .ZN(n1060) );
NAND2_X1 U754 ( .A1(KEYINPUT3), .A2(n1028), .ZN(n1058) );
NAND2_X1 U755 ( .A1(n1039), .A2(n1061), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U758 ( .A(n1030), .ZN(n1024) );
NAND2_X1 U759 ( .A1(n1066), .A2(n1067), .ZN(n1009) );
NAND2_X1 U760 ( .A1(KEYINPUT6), .A2(G952), .ZN(n1067) );
INV_X1 U761 ( .A(n1019), .ZN(n1066) );
NAND4_X1 U762 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1019) );
NOR4_X1 U763 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
XOR2_X1 U764 ( .A(n1076), .B(n1077), .Z(n1075) );
XNOR2_X1 U765 ( .A(n1078), .B(n1079), .ZN(n1074) );
XOR2_X1 U766 ( .A(KEYINPUT43), .B(KEYINPUT12), .Z(n1079) );
XOR2_X1 U767 ( .A(n1080), .B(KEYINPUT2), .Z(n1072) );
NOR3_X1 U768 ( .A1(n1049), .A2(n1081), .A3(n1064), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1069) );
XNOR2_X1 U770 ( .A(G475), .B(KEYINPUT28), .ZN(n1082) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(n1068) );
XOR2_X1 U772 ( .A(n1086), .B(KEYINPUT27), .Z(n1085) );
NAND2_X1 U773 ( .A1(KEYINPUT32), .A2(n1087), .ZN(n1084) );
XOR2_X1 U774 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U775 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U777 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U778 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U779 ( .A1(KEYINPUT22), .A2(n1098), .ZN(n1097) );
NAND3_X1 U780 ( .A1(n1099), .A2(n1100), .A3(KEYINPUT30), .ZN(n1096) );
NAND2_X1 U781 ( .A1(KEYINPUT34), .A2(n1101), .ZN(n1100) );
NAND3_X1 U782 ( .A1(G134), .A2(n1102), .A3(n1103), .ZN(n1099) );
INV_X1 U783 ( .A(KEYINPUT34), .ZN(n1103) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(n1094) );
NOR2_X1 U785 ( .A1(G900), .A2(n1010), .ZN(n1092) );
NOR2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1090) );
XNOR2_X1 U787 ( .A(G953), .B(KEYINPUT33), .ZN(n1107) );
NOR2_X1 U788 ( .A1(n1108), .A2(n1010), .ZN(n1088) );
NOR2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U790 ( .A1(n1111), .A2(n1112), .ZN(G69) );
NAND3_X1 U791 ( .A1(n1113), .A2(n1114), .A3(KEYINPUT14), .ZN(n1112) );
OR2_X1 U792 ( .A1(n1010), .A2(G224), .ZN(n1114) );
XNOR2_X1 U793 ( .A(n1115), .B(n1116), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1117), .A2(n1118), .ZN(n1111) );
NAND2_X1 U795 ( .A1(KEYINPUT14), .A2(n1119), .ZN(n1118) );
NAND2_X1 U796 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1116), .B(n1115), .Z(n1117) );
NOR2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1115) );
XNOR2_X1 U800 ( .A(n1123), .B(KEYINPUT57), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U803 ( .A(n1128), .B(KEYINPUT17), .ZN(n1126) );
OR2_X1 U804 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
NAND3_X1 U805 ( .A1(n1129), .A2(n1130), .A3(n1010), .ZN(n1116) );
OR2_X1 U806 ( .A1(n1018), .A2(KEYINPUT51), .ZN(n1130) );
NAND2_X1 U807 ( .A1(n1131), .A2(KEYINPUT51), .ZN(n1129) );
NOR2_X1 U808 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U810 ( .A1(KEYINPUT15), .A2(n1136), .ZN(n1135) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U812 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1141), .ZN(G63) );
XOR2_X1 U814 ( .A(n1142), .B(n1143), .Z(n1141) );
AND2_X1 U815 ( .A1(G478), .A2(n1139), .ZN(n1142) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1144), .ZN(G60) );
XNOR2_X1 U817 ( .A(n1145), .B(n1146), .ZN(n1144) );
AND2_X1 U818 ( .A1(G475), .A2(n1139), .ZN(n1146) );
XOR2_X1 U819 ( .A(G104), .B(n1147), .Z(G6) );
NOR3_X1 U820 ( .A1(n1041), .A2(KEYINPUT40), .A3(n1008), .ZN(n1147) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(G57) );
XNOR2_X1 U822 ( .A(n1150), .B(n1151), .ZN(n1149) );
AND2_X1 U823 ( .A1(G472), .A2(n1139), .ZN(n1151) );
INV_X1 U824 ( .A(n1152), .ZN(n1139) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1010), .ZN(n1148) );
XNOR2_X1 U826 ( .A(G952), .B(KEYINPUT54), .ZN(n1153) );
NOR2_X1 U827 ( .A1(n1132), .A2(n1154), .ZN(G54) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U830 ( .A1(KEYINPUT35), .A2(n1159), .ZN(n1158) );
NAND3_X1 U831 ( .A1(G902), .A2(G469), .A3(n1160), .ZN(n1157) );
XOR2_X1 U832 ( .A(n1161), .B(KEYINPUT8), .Z(n1160) );
NOR2_X1 U833 ( .A1(n1132), .A2(n1162), .ZN(G51) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1163) );
NOR2_X1 U837 ( .A1(n1077), .A2(n1152), .ZN(n1168) );
NAND2_X1 U838 ( .A1(G902), .A2(n1161), .ZN(n1152) );
NAND2_X1 U839 ( .A1(n1169), .A2(n1106), .ZN(n1161) );
INV_X1 U840 ( .A(n1017), .ZN(n1106) );
NAND4_X1 U841 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1017) );
AND4_X1 U842 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
AND2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
NAND3_X1 U844 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1170) );
XOR2_X1 U845 ( .A(KEYINPUT5), .B(n1028), .Z(n1181) );
XOR2_X1 U846 ( .A(n1018), .B(KEYINPUT7), .Z(n1169) );
NAND4_X1 U847 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1018) );
NOR4_X1 U848 ( .A1(n1187), .A2(n1131), .A3(n1188), .A4(n1189), .ZN(n1186) );
AND2_X1 U849 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NAND2_X1 U850 ( .A1(n1192), .A2(n1193), .ZN(n1185) );
NAND2_X1 U851 ( .A1(n1007), .A2(n1041), .ZN(n1193) );
INV_X1 U852 ( .A(n1057), .ZN(n1007) );
INV_X1 U853 ( .A(n1008), .ZN(n1192) );
NAND2_X1 U854 ( .A1(n1194), .A2(n1039), .ZN(n1008) );
XNOR2_X1 U855 ( .A(n1195), .B(n1098), .ZN(n1167) );
NAND3_X1 U856 ( .A1(G224), .A2(n1010), .A3(n1196), .ZN(n1195) );
XNOR2_X1 U857 ( .A(KEYINPUT62), .B(KEYINPUT1), .ZN(n1196) );
NOR2_X1 U858 ( .A1(n1010), .A2(G952), .ZN(n1132) );
XNOR2_X1 U859 ( .A(G146), .B(n1171), .ZN(G48) );
NAND4_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1171) );
XOR2_X1 U861 ( .A(G143), .B(n1201), .Z(G45) );
NOR2_X1 U862 ( .A1(KEYINPUT11), .A2(n1179), .ZN(n1201) );
NAND4_X1 U863 ( .A1(n1202), .A2(n1032), .A3(n1203), .A4(n1199), .ZN(n1179) );
NOR2_X1 U864 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U865 ( .A(G140), .B(n1206), .ZN(G42) );
NOR2_X1 U866 ( .A1(KEYINPUT23), .A2(n1207), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1208), .A2(n1056), .ZN(n1207) );
XOR2_X1 U868 ( .A(n1209), .B(KEYINPUT0), .Z(n1208) );
NAND2_X1 U869 ( .A1(n1198), .A2(n1028), .ZN(n1209) );
AND2_X1 U870 ( .A1(n1202), .A2(n1180), .ZN(n1198) );
XNOR2_X1 U871 ( .A(G137), .B(n1178), .ZN(G39) );
NAND2_X1 U872 ( .A1(n1182), .A2(n1210), .ZN(n1178) );
XNOR2_X1 U873 ( .A(G134), .B(n1177), .ZN(G36) );
NAND3_X1 U874 ( .A1(n1032), .A2(n1057), .A3(n1182), .ZN(n1177) );
XNOR2_X1 U875 ( .A(G131), .B(n1176), .ZN(G33) );
NAND3_X1 U876 ( .A1(n1180), .A2(n1032), .A3(n1182), .ZN(n1176) );
AND2_X1 U877 ( .A1(n1020), .A2(n1202), .ZN(n1182) );
NOR2_X1 U878 ( .A1(n1047), .A2(n1211), .ZN(n1202) );
XNOR2_X1 U879 ( .A(n1212), .B(KEYINPUT47), .ZN(n1047) );
INV_X1 U880 ( .A(n1056), .ZN(n1020) );
NAND2_X1 U881 ( .A1(n1065), .A2(n1213), .ZN(n1056) );
XNOR2_X1 U882 ( .A(G128), .B(n1175), .ZN(G30) );
NAND4_X1 U883 ( .A1(n1197), .A2(n1199), .A3(n1057), .A4(n1214), .ZN(n1175) );
NOR3_X1 U884 ( .A1(n1212), .A2(n1211), .A3(n1078), .ZN(n1214) );
INV_X1 U885 ( .A(n1215), .ZN(n1211) );
XOR2_X1 U886 ( .A(G101), .B(n1187), .Z(G3) );
AND3_X1 U887 ( .A1(n1032), .A2(n1194), .A3(n1021), .ZN(n1187) );
XNOR2_X1 U888 ( .A(G125), .B(n1174), .ZN(G27) );
NAND4_X1 U889 ( .A1(n1199), .A2(n1215), .A3(n1028), .A4(n1216), .ZN(n1174) );
NOR2_X1 U890 ( .A1(n1026), .A2(n1041), .ZN(n1216) );
NAND2_X1 U891 ( .A1(n1030), .A2(n1217), .ZN(n1215) );
NAND4_X1 U892 ( .A1(G902), .A2(G953), .A3(n1218), .A4(n1110), .ZN(n1217) );
INV_X1 U893 ( .A(G900), .ZN(n1110) );
XOR2_X1 U894 ( .A(n1219), .B(G122), .Z(G24) );
NAND2_X1 U895 ( .A1(KEYINPUT10), .A2(n1220), .ZN(n1219) );
NAND2_X1 U896 ( .A1(n1221), .A2(n1199), .ZN(n1220) );
XOR2_X1 U897 ( .A(n1222), .B(KEYINPUT63), .Z(n1221) );
NAND3_X1 U898 ( .A1(n1031), .A2(n1223), .A3(n1191), .ZN(n1222) );
AND3_X1 U899 ( .A1(n1073), .A2(n1224), .A3(n1039), .ZN(n1191) );
NAND2_X1 U900 ( .A1(n1225), .A2(n1226), .ZN(n1039) );
NAND2_X1 U901 ( .A1(n1028), .A2(n1227), .ZN(n1226) );
INV_X1 U902 ( .A(KEYINPUT49), .ZN(n1227) );
NAND3_X1 U903 ( .A1(n1228), .A2(n1078), .A3(KEYINPUT49), .ZN(n1225) );
XOR2_X1 U904 ( .A(KEYINPUT42), .B(n1229), .Z(n1223) );
INV_X1 U905 ( .A(n1026), .ZN(n1031) );
XNOR2_X1 U906 ( .A(n1230), .B(n1131), .ZN(G21) );
AND2_X1 U907 ( .A1(n1210), .A2(n1190), .ZN(n1131) );
AND3_X1 U908 ( .A1(n1197), .A2(n1200), .A3(n1021), .ZN(n1210) );
XOR2_X1 U909 ( .A(n1183), .B(n1231), .Z(G18) );
NAND2_X1 U910 ( .A1(KEYINPUT48), .A2(G116), .ZN(n1231) );
NAND3_X1 U911 ( .A1(n1032), .A2(n1057), .A3(n1190), .ZN(n1183) );
NOR2_X1 U912 ( .A1(n1224), .A2(n1205), .ZN(n1057) );
INV_X1 U913 ( .A(n1073), .ZN(n1205) );
XNOR2_X1 U914 ( .A(G113), .B(n1232), .ZN(G15) );
NAND2_X1 U915 ( .A1(KEYINPUT19), .A2(n1233), .ZN(n1232) );
INV_X1 U916 ( .A(n1184), .ZN(n1233) );
NAND3_X1 U917 ( .A1(n1180), .A2(n1032), .A3(n1190), .ZN(n1184) );
NOR3_X1 U918 ( .A1(n1062), .A2(n1229), .A3(n1026), .ZN(n1190) );
NAND2_X1 U919 ( .A1(n1050), .A2(n1234), .ZN(n1026) );
XNOR2_X1 U920 ( .A(n1235), .B(KEYINPUT59), .ZN(n1050) );
NOR2_X1 U921 ( .A1(n1197), .A2(n1078), .ZN(n1032) );
INV_X1 U922 ( .A(n1200), .ZN(n1078) );
INV_X1 U923 ( .A(n1228), .ZN(n1197) );
INV_X1 U924 ( .A(n1041), .ZN(n1180) );
NAND2_X1 U925 ( .A1(n1236), .A2(n1224), .ZN(n1041) );
XNOR2_X1 U926 ( .A(n1073), .B(KEYINPUT41), .ZN(n1236) );
XNOR2_X1 U927 ( .A(n1189), .B(n1237), .ZN(G12) );
XOR2_X1 U928 ( .A(KEYINPUT61), .B(G110), .Z(n1237) );
AND3_X1 U929 ( .A1(n1194), .A2(n1028), .A3(n1021), .ZN(n1189) );
NOR2_X1 U930 ( .A1(n1073), .A2(n1224), .ZN(n1021) );
INV_X1 U931 ( .A(n1204), .ZN(n1224) );
NOR2_X1 U932 ( .A1(n1238), .A2(n1081), .ZN(n1204) );
NOR2_X1 U933 ( .A1(n1083), .A2(G475), .ZN(n1081) );
AND2_X1 U934 ( .A1(G475), .A2(n1083), .ZN(n1238) );
NAND2_X1 U935 ( .A1(n1145), .A2(n1239), .ZN(n1083) );
XNOR2_X1 U936 ( .A(n1240), .B(n1241), .ZN(n1145) );
XOR2_X1 U937 ( .A(n1105), .B(n1242), .Z(n1241) );
XOR2_X1 U938 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR2_X1 U939 ( .A1(G122), .A2(KEYINPUT25), .ZN(n1243) );
XOR2_X1 U940 ( .A(n1245), .B(n1246), .Z(n1240) );
XOR2_X1 U941 ( .A(G143), .B(G113), .Z(n1246) );
XNOR2_X1 U942 ( .A(G104), .B(n1247), .ZN(n1245) );
NOR2_X1 U943 ( .A1(n1248), .A2(KEYINPUT9), .ZN(n1247) );
AND2_X1 U944 ( .A1(n1249), .A2(G214), .ZN(n1248) );
XNOR2_X1 U945 ( .A(n1250), .B(G478), .ZN(n1073) );
OR2_X1 U946 ( .A1(n1143), .A2(G902), .ZN(n1250) );
XNOR2_X1 U947 ( .A(n1251), .B(n1252), .ZN(n1143) );
XOR2_X1 U948 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U949 ( .A(n1255), .B(n1256), .Z(n1254) );
AND3_X1 U950 ( .A1(G234), .A2(n1010), .A3(G217), .ZN(n1256) );
NAND2_X1 U951 ( .A1(KEYINPUT29), .A2(n1257), .ZN(n1255) );
NAND2_X1 U952 ( .A1(KEYINPUT44), .A2(n1005), .ZN(n1253) );
INV_X1 U953 ( .A(G107), .ZN(n1005) );
XNOR2_X1 U954 ( .A(G116), .B(n1258), .ZN(n1251) );
XOR2_X1 U955 ( .A(G134), .B(G122), .Z(n1258) );
NOR2_X1 U956 ( .A1(n1228), .A2(n1200), .ZN(n1028) );
XNOR2_X1 U957 ( .A(n1259), .B(G472), .ZN(n1200) );
NAND2_X1 U958 ( .A1(n1150), .A2(n1239), .ZN(n1259) );
XNOR2_X1 U959 ( .A(n1260), .B(n1261), .ZN(n1150) );
XOR2_X1 U960 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U961 ( .A(n1264), .B(G101), .Z(n1263) );
NAND2_X1 U962 ( .A1(G210), .A2(n1249), .ZN(n1264) );
NOR2_X1 U963 ( .A1(G953), .A2(G237), .ZN(n1249) );
XNOR2_X1 U964 ( .A(G131), .B(G113), .ZN(n1262) );
XNOR2_X1 U965 ( .A(n1265), .B(n1101), .ZN(n1260) );
XNOR2_X1 U966 ( .A(n1165), .B(n1266), .ZN(n1265) );
XNOR2_X1 U967 ( .A(n1080), .B(KEYINPUT38), .ZN(n1228) );
XOR2_X1 U968 ( .A(n1267), .B(n1140), .Z(n1080) );
AND2_X1 U969 ( .A1(G217), .A2(n1268), .ZN(n1140) );
NAND2_X1 U970 ( .A1(n1269), .A2(n1239), .ZN(n1267) );
XNOR2_X1 U971 ( .A(n1137), .B(n1138), .ZN(n1269) );
XOR2_X1 U972 ( .A(G119), .B(n1270), .Z(n1138) );
XOR2_X1 U973 ( .A(G140), .B(G128), .Z(n1270) );
XOR2_X1 U974 ( .A(n1271), .B(n1272), .Z(n1137) );
XOR2_X1 U975 ( .A(n1273), .B(n1244), .Z(n1271) );
XNOR2_X1 U976 ( .A(n1098), .B(G146), .ZN(n1244) );
NAND3_X1 U977 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
OR2_X1 U978 ( .A1(n1277), .A2(KEYINPUT4), .ZN(n1276) );
NAND3_X1 U979 ( .A1(KEYINPUT4), .A2(n1277), .A3(n1102), .ZN(n1275) );
INV_X1 U980 ( .A(G137), .ZN(n1102) );
NAND2_X1 U981 ( .A1(G137), .A2(n1278), .ZN(n1274) );
NAND2_X1 U982 ( .A1(KEYINPUT4), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U983 ( .A(KEYINPUT55), .B(n1277), .ZN(n1279) );
NAND3_X1 U984 ( .A1(G221), .A2(G234), .A3(n1280), .ZN(n1277) );
XNOR2_X1 U985 ( .A(G953), .B(KEYINPUT20), .ZN(n1280) );
NOR3_X1 U986 ( .A1(n1212), .A2(n1229), .A3(n1062), .ZN(n1194) );
INV_X1 U987 ( .A(n1199), .ZN(n1062) );
NOR2_X1 U988 ( .A1(n1065), .A2(n1064), .ZN(n1199) );
INV_X1 U989 ( .A(n1213), .ZN(n1064) );
NAND2_X1 U990 ( .A1(G214), .A2(n1281), .ZN(n1213) );
XOR2_X1 U991 ( .A(n1282), .B(n1076), .Z(n1065) );
NAND2_X1 U992 ( .A1(n1283), .A2(n1239), .ZN(n1076) );
XOR2_X1 U993 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U994 ( .A(n1166), .B(n1286), .ZN(n1285) );
NOR2_X1 U995 ( .A1(KEYINPUT24), .A2(n1165), .ZN(n1286) );
XOR2_X1 U996 ( .A(G146), .B(n1257), .Z(n1165) );
XNOR2_X1 U997 ( .A(n1127), .B(n1287), .ZN(n1166) );
XNOR2_X1 U998 ( .A(n1288), .B(KEYINPUT58), .ZN(n1287) );
NAND2_X1 U999 ( .A1(KEYINPUT31), .A2(n1128), .ZN(n1288) );
XNOR2_X1 U1000 ( .A(n1289), .B(n1290), .ZN(n1128) );
XOR2_X1 U1001 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U1002 ( .A(G104), .B(n1293), .Z(n1292) );
NOR2_X1 U1003 ( .A1(G101), .A2(KEYINPUT13), .ZN(n1293) );
NOR2_X1 U1004 ( .A1(n1294), .A2(n1295), .ZN(n1291) );
AND3_X1 U1005 ( .A1(KEYINPUT36), .A2(n1230), .A3(G116), .ZN(n1295) );
NOR2_X1 U1006 ( .A1(KEYINPUT36), .A2(n1266), .ZN(n1294) );
XNOR2_X1 U1007 ( .A(G116), .B(n1230), .ZN(n1266) );
INV_X1 U1008 ( .A(G119), .ZN(n1230) );
XNOR2_X1 U1009 ( .A(G107), .B(n1296), .ZN(n1289) );
XOR2_X1 U1010 ( .A(KEYINPUT50), .B(G113), .Z(n1296) );
XNOR2_X1 U1011 ( .A(G122), .B(n1272), .ZN(n1127) );
XOR2_X1 U1012 ( .A(n1297), .B(n1298), .Z(n1284) );
XNOR2_X1 U1013 ( .A(KEYINPUT18), .B(n1098), .ZN(n1298) );
INV_X1 U1014 ( .A(G125), .ZN(n1098) );
NAND2_X1 U1015 ( .A1(G224), .A2(n1010), .ZN(n1297) );
NAND2_X1 U1016 ( .A1(KEYINPUT21), .A2(n1077), .ZN(n1282) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1281), .ZN(n1077) );
NAND2_X1 U1018 ( .A1(n1299), .A2(n1239), .ZN(n1281) );
INV_X1 U1019 ( .A(G237), .ZN(n1299) );
AND2_X1 U1020 ( .A1(n1030), .A2(n1300), .ZN(n1229) );
NAND3_X1 U1021 ( .A1(n1122), .A2(n1218), .A3(G902), .ZN(n1300) );
NOR2_X1 U1022 ( .A1(n1010), .A2(G898), .ZN(n1122) );
NAND3_X1 U1023 ( .A1(n1218), .A2(n1010), .A3(G952), .ZN(n1030) );
INV_X1 U1024 ( .A(G953), .ZN(n1010) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1218) );
OR2_X1 U1026 ( .A1(n1235), .A2(n1049), .ZN(n1212) );
INV_X1 U1027 ( .A(n1234), .ZN(n1049) );
NAND2_X1 U1028 ( .A1(G221), .A2(n1268), .ZN(n1234) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1239), .ZN(n1268) );
XNOR2_X1 U1030 ( .A(n1086), .B(n1087), .ZN(n1235) );
XNOR2_X1 U1031 ( .A(G469), .B(KEYINPUT60), .ZN(n1087) );
NAND2_X1 U1032 ( .A1(n1301), .A2(n1239), .ZN(n1086) );
INV_X1 U1033 ( .A(G902), .ZN(n1239) );
XOR2_X1 U1034 ( .A(n1302), .B(n1155), .Z(n1301) );
XNOR2_X1 U1035 ( .A(n1303), .B(n1304), .ZN(n1155) );
XNOR2_X1 U1036 ( .A(n1101), .B(n1105), .ZN(n1304) );
XOR2_X1 U1037 ( .A(G131), .B(G140), .Z(n1105) );
XNOR2_X1 U1038 ( .A(G134), .B(G137), .ZN(n1101) );
XNOR2_X1 U1039 ( .A(n1272), .B(n1305), .ZN(n1303) );
XOR2_X1 U1040 ( .A(KEYINPUT16), .B(n1306), .Z(n1305) );
NOR2_X1 U1041 ( .A1(G953), .A2(n1109), .ZN(n1306) );
INV_X1 U1042 ( .A(G227), .ZN(n1109) );
XOR2_X1 U1043 ( .A(G110), .B(KEYINPUT26), .Z(n1272) );
NOR2_X1 U1044 ( .A1(KEYINPUT39), .A2(n1159), .ZN(n1302) );
XOR2_X1 U1045 ( .A(n1307), .B(n1308), .Z(n1159) );
XOR2_X1 U1046 ( .A(n1309), .B(n1104), .Z(n1308) );
NAND2_X1 U1047 ( .A1(n1310), .A2(n1311), .ZN(n1104) );
NAND2_X1 U1048 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
INV_X1 U1049 ( .A(G146), .ZN(n1313) );
XOR2_X1 U1050 ( .A(KEYINPUT52), .B(n1257), .Z(n1312) );
NAND2_X1 U1051 ( .A1(G146), .A2(n1257), .ZN(n1310) );
XOR2_X1 U1052 ( .A(G128), .B(G143), .Z(n1257) );
NAND2_X1 U1053 ( .A1(KEYINPUT56), .A2(G107), .ZN(n1309) );
XNOR2_X1 U1054 ( .A(G104), .B(n1314), .ZN(n1307) );
NOR2_X1 U1055 ( .A1(G101), .A2(KEYINPUT37), .ZN(n1314) );
endmodule


