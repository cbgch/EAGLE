//Key = 0010100000100001000100111101100010011110110011000011010101010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297;

XNOR2_X1 U715 ( .A(n978), .B(n979), .ZN(G9) );
XNOR2_X1 U716 ( .A(G107), .B(KEYINPUT12), .ZN(n979) );
NOR2_X1 U717 ( .A1(n980), .A2(n981), .ZN(G75) );
NOR3_X1 U718 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n981) );
XOR2_X1 U719 ( .A(KEYINPUT60), .B(n985), .Z(n984) );
NAND3_X1 U720 ( .A1(n986), .A2(n987), .A3(G952), .ZN(n982) );
NAND2_X1 U721 ( .A1(n988), .A2(n989), .ZN(n986) );
NAND2_X1 U722 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND3_X1 U723 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND2_X1 U724 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND2_X1 U725 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U726 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U727 ( .A1(n1001), .A2(n1002), .ZN(n995) );
NAND2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U729 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND3_X1 U730 ( .A1(n997), .A2(n1007), .A3(n1001), .ZN(n990) );
NAND2_X1 U731 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U732 ( .A1(n994), .A2(n1010), .ZN(n1009) );
OR2_X1 U733 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U734 ( .A1(n992), .A2(n1013), .ZN(n1008) );
NAND2_X1 U735 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U736 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U737 ( .A(n1018), .ZN(n988) );
NOR3_X1 U738 ( .A1(n1019), .A2(G953), .A3(n985), .ZN(n980) );
AND3_X1 U739 ( .A1(n994), .A2(n1020), .A3(n997), .ZN(n985) );
INV_X1 U740 ( .A(n1021), .ZN(n997) );
XOR2_X1 U741 ( .A(KEYINPUT34), .B(n1022), .Z(n1020) );
NOR4_X1 U742 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
XNOR2_X1 U743 ( .A(G472), .B(n1027), .ZN(n1026) );
NAND2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U745 ( .A1(KEYINPUT23), .A2(n1030), .ZN(n1029) );
NAND2_X1 U746 ( .A1(KEYINPUT11), .A2(n1031), .ZN(n1028) );
XOR2_X1 U747 ( .A(KEYINPUT48), .B(n1032), .Z(n1024) );
NOR2_X1 U748 ( .A1(G475), .A2(n1033), .ZN(n1032) );
NAND3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1023) );
NAND2_X1 U750 ( .A1(G475), .A2(n1033), .ZN(n1036) );
NAND2_X1 U751 ( .A1(G478), .A2(n1037), .ZN(n1034) );
XOR2_X1 U752 ( .A(KEYINPUT17), .B(G952), .Z(n1019) );
XOR2_X1 U753 ( .A(n1038), .B(n1039), .Z(G72) );
XOR2_X1 U754 ( .A(n1040), .B(n1041), .Z(n1039) );
NAND2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1044), .A2(G953), .ZN(n1043) );
XNOR2_X1 U757 ( .A(G900), .B(KEYINPUT13), .ZN(n1044) );
XOR2_X1 U758 ( .A(n1045), .B(n1046), .Z(n1042) );
XNOR2_X1 U759 ( .A(n1047), .B(n1048), .ZN(n1046) );
NAND3_X1 U760 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1047) );
NAND2_X1 U761 ( .A1(KEYINPUT5), .A2(n1052), .ZN(n1050) );
NAND2_X1 U762 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XNOR2_X1 U763 ( .A(KEYINPUT6), .B(n1055), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1049) );
INV_X1 U765 ( .A(KEYINPUT5), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
OR3_X1 U767 ( .A1(n1055), .A2(G137), .A3(KEYINPUT6), .ZN(n1059) );
NAND2_X1 U768 ( .A1(KEYINPUT6), .A2(n1055), .ZN(n1058) );
NAND2_X1 U769 ( .A1(G953), .A2(n1060), .ZN(n1040) );
NAND2_X1 U770 ( .A1(n1061), .A2(G900), .ZN(n1060) );
XNOR2_X1 U771 ( .A(G227), .B(KEYINPUT27), .ZN(n1061) );
NOR2_X1 U772 ( .A1(n1062), .A2(G953), .ZN(n1038) );
NAND2_X1 U773 ( .A1(n1063), .A2(n1064), .ZN(G69) );
NAND2_X1 U774 ( .A1(n1065), .A2(n987), .ZN(n1064) );
XNOR2_X1 U775 ( .A(n1066), .B(n1067), .ZN(n1065) );
NOR2_X1 U776 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XNOR2_X1 U777 ( .A(KEYINPUT51), .B(KEYINPUT0), .ZN(n1069) );
NAND2_X1 U778 ( .A1(n1070), .A2(G953), .ZN(n1063) );
XOR2_X1 U779 ( .A(n1066), .B(n1071), .Z(n1070) );
AND2_X1 U780 ( .A1(G224), .A2(G898), .ZN(n1071) );
NAND2_X1 U781 ( .A1(n1072), .A2(n1073), .ZN(n1066) );
NAND2_X1 U782 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U783 ( .A(n1075), .B(n1076), .ZN(n1072) );
XOR2_X1 U784 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U785 ( .A1(n1079), .A2(KEYINPUT42), .ZN(n1077) );
NOR2_X1 U786 ( .A1(n1080), .A2(n1081), .ZN(G66) );
XOR2_X1 U787 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U788 ( .A(KEYINPUT53), .B(n1084), .Z(n1083) );
NOR2_X1 U789 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U790 ( .A1(n1080), .A2(n1087), .ZN(G63) );
NOR2_X1 U791 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U792 ( .A(n1090), .B(KEYINPUT59), .Z(n1089) );
NAND2_X1 U793 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U794 ( .A(KEYINPUT33), .B(n1093), .ZN(n1092) );
NOR2_X1 U795 ( .A1(n1094), .A2(n1091), .ZN(n1088) );
NOR2_X1 U796 ( .A1(n1086), .A2(n1095), .ZN(n1091) );
INV_X1 U797 ( .A(G478), .ZN(n1095) );
INV_X1 U798 ( .A(n1093), .ZN(n1094) );
NOR2_X1 U799 ( .A1(n1080), .A2(n1096), .ZN(G60) );
XOR2_X1 U800 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND3_X1 U801 ( .A1(G475), .A2(G902), .A3(n1099), .ZN(n1097) );
XOR2_X1 U802 ( .A(n983), .B(KEYINPUT3), .Z(n1099) );
XNOR2_X1 U803 ( .A(G104), .B(n1100), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1080), .A2(n1101), .ZN(G57) );
XOR2_X1 U805 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U806 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U807 ( .A1(n1106), .A2(n1086), .ZN(n1104) );
INV_X1 U808 ( .A(G472), .ZN(n1106) );
XOR2_X1 U809 ( .A(n1107), .B(n1108), .Z(n1102) );
NOR2_X1 U810 ( .A1(KEYINPUT47), .A2(n1109), .ZN(n1108) );
NOR2_X1 U811 ( .A1(KEYINPUT1), .A2(n1110), .ZN(n1107) );
XNOR2_X1 U812 ( .A(n1111), .B(n1112), .ZN(n1110) );
NAND2_X1 U813 ( .A1(n1113), .A2(KEYINPUT41), .ZN(n1111) );
XNOR2_X1 U814 ( .A(G131), .B(n1114), .ZN(n1113) );
NOR2_X1 U815 ( .A1(n1080), .A2(n1115), .ZN(G54) );
XOR2_X1 U816 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U817 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U818 ( .A1(n1120), .A2(n1086), .ZN(n1118) );
XOR2_X1 U819 ( .A(n1121), .B(n1122), .Z(n1116) );
NAND2_X1 U820 ( .A1(n1123), .A2(KEYINPUT35), .ZN(n1122) );
XNOR2_X1 U821 ( .A(n1124), .B(n1125), .ZN(n1123) );
NAND2_X1 U822 ( .A1(KEYINPUT45), .A2(G140), .ZN(n1124) );
NOR2_X1 U823 ( .A1(n1080), .A2(n1126), .ZN(G51) );
XOR2_X1 U824 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U825 ( .A1(n1129), .A2(n1086), .ZN(n1128) );
NAND2_X1 U826 ( .A1(G902), .A2(n983), .ZN(n1086) );
NAND2_X1 U827 ( .A1(n1062), .A2(n1068), .ZN(n983) );
AND2_X1 U828 ( .A1(n1130), .A2(n1131), .ZN(n1068) );
NOR4_X1 U829 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n978), .ZN(n1131) );
AND3_X1 U830 ( .A1(n992), .A2(n1135), .A3(n1136), .ZN(n978) );
NOR4_X1 U831 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1130) );
NOR2_X1 U832 ( .A1(n1141), .A2(n1014), .ZN(n1140) );
XOR2_X1 U833 ( .A(n1142), .B(KEYINPUT58), .Z(n1141) );
AND3_X1 U834 ( .A1(n1001), .A2(n1136), .A3(n1011), .ZN(n1139) );
INV_X1 U835 ( .A(n1100), .ZN(n1138) );
NAND3_X1 U836 ( .A1(n1136), .A2(n992), .A3(n1143), .ZN(n1100) );
INV_X1 U837 ( .A(n1144), .ZN(n1137) );
AND4_X1 U838 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1062) );
NOR4_X1 U839 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NOR3_X1 U840 ( .A1(n1153), .A2(n1014), .A3(n1000), .ZN(n1152) );
NOR4_X1 U841 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n999), .ZN(n1151) );
XNOR2_X1 U842 ( .A(n994), .B(KEYINPUT16), .ZN(n1154) );
INV_X1 U843 ( .A(n1157), .ZN(n1150) );
NOR2_X1 U844 ( .A1(n1158), .A2(n1159), .ZN(n1147) );
INV_X1 U845 ( .A(n1160), .ZN(n1159) );
NAND2_X1 U846 ( .A1(n1161), .A2(n1162), .ZN(n1127) );
XNOR2_X1 U847 ( .A(KEYINPUT40), .B(KEYINPUT19), .ZN(n1161) );
NOR2_X1 U848 ( .A1(n987), .A2(G952), .ZN(n1080) );
XOR2_X1 U849 ( .A(G146), .B(n1158), .Z(G48) );
NOR3_X1 U850 ( .A1(n1153), .A2(n1014), .A3(n999), .ZN(n1158) );
XNOR2_X1 U851 ( .A(G143), .B(n1157), .ZN(G45) );
NAND3_X1 U852 ( .A1(n1163), .A2(n1011), .A3(n1164), .ZN(n1157) );
NOR3_X1 U853 ( .A1(n1014), .A2(n1165), .A3(n1166), .ZN(n1164) );
XOR2_X1 U854 ( .A(G140), .B(n1149), .Z(G42) );
AND2_X1 U855 ( .A1(n1167), .A2(n1012), .ZN(n1149) );
XNOR2_X1 U856 ( .A(G137), .B(n1145), .ZN(G39) );
NAND3_X1 U857 ( .A1(n1001), .A2(n994), .A3(n1168), .ZN(n1145) );
INV_X1 U858 ( .A(n1153), .ZN(n1168) );
XNOR2_X1 U859 ( .A(G134), .B(n1146), .ZN(G36) );
NAND4_X1 U860 ( .A1(n1163), .A2(n1011), .A3(n994), .A4(n1135), .ZN(n1146) );
INV_X1 U861 ( .A(n1169), .ZN(n994) );
XNOR2_X1 U862 ( .A(n1170), .B(n1171), .ZN(G33) );
AND2_X1 U863 ( .A1(n1011), .A2(n1167), .ZN(n1171) );
NOR3_X1 U864 ( .A1(n1156), .A2(n1169), .A3(n999), .ZN(n1167) );
INV_X1 U865 ( .A(n1143), .ZN(n999) );
NAND2_X1 U866 ( .A1(n1017), .A2(n1172), .ZN(n1169) );
INV_X1 U867 ( .A(n1163), .ZN(n1156) );
XOR2_X1 U868 ( .A(G128), .B(n1173), .Z(G30) );
NOR4_X1 U869 ( .A1(KEYINPUT14), .A2(n1014), .A3(n1000), .A4(n1153), .ZN(n1173) );
NAND3_X1 U870 ( .A1(n1174), .A2(n1025), .A3(n1163), .ZN(n1153) );
NOR2_X1 U871 ( .A1(n1003), .A2(n1175), .ZN(n1163) );
INV_X1 U872 ( .A(n1135), .ZN(n1000) );
XOR2_X1 U873 ( .A(n1176), .B(n1177), .Z(G3) );
XNOR2_X1 U874 ( .A(KEYINPUT22), .B(n1178), .ZN(n1177) );
NAND4_X1 U875 ( .A1(KEYINPUT36), .A2(n1001), .A3(n1011), .A4(n1136), .ZN(n1176) );
XNOR2_X1 U876 ( .A(G125), .B(n1160), .ZN(G27) );
NAND3_X1 U877 ( .A1(n1012), .A2(n1143), .A3(n1179), .ZN(n1160) );
NOR3_X1 U878 ( .A1(n1021), .A2(n1175), .A3(n1014), .ZN(n1179) );
AND2_X1 U879 ( .A1(n1180), .A2(n1018), .ZN(n1175) );
NAND2_X1 U880 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
INV_X1 U881 ( .A(G900), .ZN(n1182) );
XOR2_X1 U882 ( .A(n1134), .B(n1183), .Z(G24) );
NOR2_X1 U883 ( .A1(KEYINPUT63), .A2(n1184), .ZN(n1183) );
AND4_X1 U884 ( .A1(n1185), .A2(n992), .A3(n1186), .A4(n1187), .ZN(n1134) );
NOR2_X1 U885 ( .A1(n1025), .A2(n1174), .ZN(n992) );
XOR2_X1 U886 ( .A(G119), .B(n1188), .Z(G21) );
NOR2_X1 U887 ( .A1(n1189), .A2(n1142), .ZN(n1188) );
NAND3_X1 U888 ( .A1(n1174), .A2(n1001), .A3(n1190), .ZN(n1142) );
NOR3_X1 U889 ( .A1(n1021), .A2(n1191), .A3(n1192), .ZN(n1190) );
XOR2_X1 U890 ( .A(n1014), .B(KEYINPUT54), .Z(n1189) );
XOR2_X1 U891 ( .A(n1133), .B(n1193), .Z(G18) );
NOR2_X1 U892 ( .A1(KEYINPUT8), .A2(n1194), .ZN(n1193) );
AND3_X1 U893 ( .A1(n1011), .A2(n1135), .A3(n1185), .ZN(n1133) );
NOR2_X1 U894 ( .A1(n1186), .A2(n1165), .ZN(n1135) );
INV_X1 U895 ( .A(n1187), .ZN(n1165) );
XOR2_X1 U896 ( .A(G113), .B(n1132), .Z(G15) );
AND3_X1 U897 ( .A1(n1143), .A2(n1011), .A3(n1185), .ZN(n1132) );
NOR3_X1 U898 ( .A1(n1014), .A2(n1191), .A3(n1021), .ZN(n1185) );
NAND2_X1 U899 ( .A1(n1006), .A2(n1195), .ZN(n1021) );
INV_X1 U900 ( .A(n1155), .ZN(n1011) );
NAND2_X1 U901 ( .A1(n1174), .A2(n1192), .ZN(n1155) );
NOR2_X1 U902 ( .A1(n1187), .A2(n1166), .ZN(n1143) );
INV_X1 U903 ( .A(n1186), .ZN(n1166) );
XNOR2_X1 U904 ( .A(G110), .B(n1144), .ZN(G12) );
NAND3_X1 U905 ( .A1(n1001), .A2(n1136), .A3(n1012), .ZN(n1144) );
NOR2_X1 U906 ( .A1(n1192), .A2(n1174), .ZN(n1012) );
XNOR2_X1 U907 ( .A(G472), .B(n1196), .ZN(n1174) );
NOR2_X1 U908 ( .A1(n1031), .A2(KEYINPUT43), .ZN(n1196) );
INV_X1 U909 ( .A(n1030), .ZN(n1031) );
NAND2_X1 U910 ( .A1(n1197), .A2(n1198), .ZN(n1030) );
XNOR2_X1 U911 ( .A(n1199), .B(n1200), .ZN(n1197) );
XOR2_X1 U912 ( .A(n1105), .B(n1109), .Z(n1200) );
NAND3_X1 U913 ( .A1(n1201), .A2(n987), .A3(G210), .ZN(n1109) );
XOR2_X1 U914 ( .A(G101), .B(n1078), .Z(n1105) );
INV_X1 U915 ( .A(n1025), .ZN(n1192) );
XOR2_X1 U916 ( .A(n1202), .B(n1085), .Z(n1025) );
NAND2_X1 U917 ( .A1(G217), .A2(n1203), .ZN(n1085) );
NAND2_X1 U918 ( .A1(n1082), .A2(n1204), .ZN(n1202) );
XOR2_X1 U919 ( .A(KEYINPUT29), .B(n1198), .Z(n1204) );
XOR2_X1 U920 ( .A(n1205), .B(n1206), .Z(n1082) );
XOR2_X1 U921 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U922 ( .A(n1054), .B(G119), .ZN(n1208) );
XOR2_X1 U923 ( .A(KEYINPUT9), .B(KEYINPUT38), .Z(n1207) );
XOR2_X1 U924 ( .A(n1209), .B(n1210), .Z(n1205) );
XNOR2_X1 U925 ( .A(n1211), .B(n1212), .ZN(n1210) );
XNOR2_X1 U926 ( .A(G110), .B(n1213), .ZN(n1209) );
AND3_X1 U927 ( .A1(G221), .A2(n987), .A3(G234), .ZN(n1213) );
NOR3_X1 U928 ( .A1(n1003), .A2(n1191), .A3(n1014), .ZN(n1136) );
OR2_X1 U929 ( .A1(n1017), .A2(n1016), .ZN(n1014) );
INV_X1 U930 ( .A(n1172), .ZN(n1016) );
NAND2_X1 U931 ( .A1(G214), .A2(n1214), .ZN(n1172) );
XNOR2_X1 U932 ( .A(n1215), .B(n1129), .ZN(n1017) );
NAND2_X1 U933 ( .A1(G210), .A2(n1214), .ZN(n1129) );
NAND2_X1 U934 ( .A1(n1201), .A2(n1216), .ZN(n1214) );
NAND2_X1 U935 ( .A1(n1162), .A2(n1198), .ZN(n1215) );
XNOR2_X1 U936 ( .A(n1217), .B(n1218), .ZN(n1162) );
XNOR2_X1 U937 ( .A(n1219), .B(n1075), .ZN(n1218) );
XOR2_X1 U938 ( .A(n1220), .B(n1184), .Z(n1075) );
NAND2_X1 U939 ( .A1(KEYINPUT55), .A2(n1125), .ZN(n1220) );
INV_X1 U940 ( .A(n1112), .ZN(n1219) );
XOR2_X1 U941 ( .A(n1221), .B(n1222), .Z(n1217) );
AND2_X1 U942 ( .A1(n987), .A2(G224), .ZN(n1222) );
XNOR2_X1 U943 ( .A(n1223), .B(n1224), .ZN(n1221) );
INV_X1 U944 ( .A(G125), .ZN(n1224) );
NAND2_X1 U945 ( .A1(n1225), .A2(KEYINPUT44), .ZN(n1223) );
XNOR2_X1 U946 ( .A(n1079), .B(n1078), .ZN(n1225) );
XNOR2_X1 U947 ( .A(n1226), .B(n1227), .ZN(n1078) );
XNOR2_X1 U948 ( .A(G116), .B(G119), .ZN(n1226) );
AND2_X1 U949 ( .A1(n1228), .A2(n1229), .ZN(n1079) );
NAND2_X1 U950 ( .A1(n1230), .A2(G101), .ZN(n1229) );
XNOR2_X1 U951 ( .A(n1231), .B(n1232), .ZN(n1230) );
XOR2_X1 U952 ( .A(n1233), .B(KEYINPUT31), .Z(n1228) );
NAND2_X1 U953 ( .A1(n1234), .A2(n1178), .ZN(n1233) );
XNOR2_X1 U954 ( .A(G104), .B(n1231), .ZN(n1234) );
NAND2_X1 U955 ( .A1(KEYINPUT10), .A2(n1235), .ZN(n1231) );
XNOR2_X1 U956 ( .A(KEYINPUT32), .B(n1236), .ZN(n1235) );
AND2_X1 U957 ( .A1(n1237), .A2(n1018), .ZN(n1191) );
NAND3_X1 U958 ( .A1(n1238), .A2(n987), .A3(G952), .ZN(n1018) );
NAND2_X1 U959 ( .A1(n1181), .A2(n1074), .ZN(n1237) );
XOR2_X1 U960 ( .A(KEYINPUT37), .B(G898), .Z(n1074) );
AND3_X1 U961 ( .A1(G902), .A2(n1238), .A3(G953), .ZN(n1181) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1238) );
OR2_X1 U963 ( .A1(n1006), .A2(n1005), .ZN(n1003) );
INV_X1 U964 ( .A(n1195), .ZN(n1005) );
NAND2_X1 U965 ( .A1(G221), .A2(n1203), .ZN(n1195) );
NAND2_X1 U966 ( .A1(G234), .A2(n1216), .ZN(n1203) );
XNOR2_X1 U967 ( .A(n1239), .B(n1120), .ZN(n1006) );
INV_X1 U968 ( .A(G469), .ZN(n1120) );
NAND3_X1 U969 ( .A1(n1240), .A2(n1241), .A3(n1198), .ZN(n1239) );
NAND2_X1 U970 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
INV_X1 U971 ( .A(KEYINPUT7), .ZN(n1243) );
XNOR2_X1 U972 ( .A(n1244), .B(n1245), .ZN(n1242) );
NOR2_X1 U973 ( .A1(KEYINPUT26), .A2(n1246), .ZN(n1244) );
NAND3_X1 U974 ( .A1(n1246), .A2(n1245), .A3(KEYINPUT7), .ZN(n1240) );
XOR2_X1 U975 ( .A(n1247), .B(KEYINPUT56), .Z(n1245) );
NAND2_X1 U976 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U977 ( .A1(KEYINPUT50), .A2(n1119), .ZN(n1249) );
XOR2_X1 U978 ( .A(n1250), .B(n1199), .Z(n1119) );
XNOR2_X1 U979 ( .A(n1114), .B(n1045), .ZN(n1199) );
XNOR2_X1 U980 ( .A(n1170), .B(n1112), .ZN(n1045) );
NAND3_X1 U981 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1248) );
INV_X1 U982 ( .A(KEYINPUT50), .ZN(n1253) );
XNOR2_X1 U983 ( .A(n1114), .B(n1170), .ZN(n1252) );
NAND2_X1 U984 ( .A1(n1254), .A2(n1255), .ZN(n1114) );
NAND2_X1 U985 ( .A1(KEYINPUT46), .A2(n1256), .ZN(n1255) );
NAND2_X1 U986 ( .A1(n1051), .A2(n1257), .ZN(n1256) );
NAND2_X1 U987 ( .A1(G134), .A2(n1054), .ZN(n1257) );
INV_X1 U988 ( .A(G137), .ZN(n1054) );
NAND2_X1 U989 ( .A1(G137), .A2(n1055), .ZN(n1051) );
INV_X1 U990 ( .A(G134), .ZN(n1055) );
NAND2_X1 U991 ( .A1(n1258), .A2(n1259), .ZN(n1254) );
INV_X1 U992 ( .A(KEYINPUT46), .ZN(n1259) );
XNOR2_X1 U993 ( .A(G137), .B(G134), .ZN(n1258) );
XNOR2_X1 U994 ( .A(n1112), .B(n1250), .ZN(n1251) );
XNOR2_X1 U995 ( .A(n1260), .B(n1261), .ZN(n1250) );
XNOR2_X1 U996 ( .A(KEYINPUT25), .B(n1178), .ZN(n1261) );
INV_X1 U997 ( .A(G101), .ZN(n1178) );
NAND3_X1 U998 ( .A1(KEYINPUT2), .A2(n1262), .A3(n1263), .ZN(n1260) );
XOR2_X1 U999 ( .A(n1264), .B(KEYINPUT20), .Z(n1263) );
NAND2_X1 U1000 ( .A1(G104), .A2(n1236), .ZN(n1264) );
NAND2_X1 U1001 ( .A1(G107), .A2(n1232), .ZN(n1262) );
XOR2_X1 U1002 ( .A(G143), .B(n1212), .Z(n1112) );
XOR2_X1 U1003 ( .A(G128), .B(G146), .Z(n1212) );
XOR2_X1 U1004 ( .A(n1121), .B(n1265), .Z(n1246) );
XNOR2_X1 U1005 ( .A(G140), .B(n1125), .ZN(n1265) );
INV_X1 U1006 ( .A(G110), .ZN(n1125) );
NAND2_X1 U1007 ( .A1(G227), .A2(n987), .ZN(n1121) );
NOR2_X1 U1008 ( .A1(n1187), .A2(n1186), .ZN(n1001) );
XNOR2_X1 U1009 ( .A(n1033), .B(n1266), .ZN(n1186) );
XOR2_X1 U1010 ( .A(KEYINPUT30), .B(G475), .Z(n1266) );
NAND2_X1 U1011 ( .A1(n1098), .A2(n1198), .ZN(n1033) );
XOR2_X1 U1012 ( .A(n1267), .B(n1268), .Z(n1098) );
XOR2_X1 U1013 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U1014 ( .A(n1184), .B(n1271), .ZN(n1270) );
AND3_X1 U1015 ( .A1(G214), .A2(n987), .A3(n1201), .ZN(n1271) );
INV_X1 U1016 ( .A(G237), .ZN(n1201) );
XNOR2_X1 U1017 ( .A(G146), .B(n1170), .ZN(n1269) );
INV_X1 U1018 ( .A(G131), .ZN(n1170) );
XOR2_X1 U1019 ( .A(n1272), .B(n1273), .Z(n1267) );
XNOR2_X1 U1020 ( .A(n1227), .B(n1211), .ZN(n1273) );
INV_X1 U1021 ( .A(n1048), .ZN(n1211) );
XOR2_X1 U1022 ( .A(G125), .B(G140), .Z(n1048) );
XOR2_X1 U1023 ( .A(G113), .B(KEYINPUT18), .Z(n1227) );
XOR2_X1 U1024 ( .A(n1274), .B(n1275), .Z(n1272) );
NOR2_X1 U1025 ( .A1(KEYINPUT21), .A2(n1232), .ZN(n1275) );
INV_X1 U1026 ( .A(G104), .ZN(n1232) );
NAND2_X1 U1027 ( .A1(KEYINPUT61), .A2(n1276), .ZN(n1274) );
INV_X1 U1028 ( .A(G143), .ZN(n1276) );
NAND3_X1 U1029 ( .A1(n1277), .A2(n1278), .A3(n1035), .ZN(n1187) );
OR2_X1 U1030 ( .A1(n1037), .A2(G478), .ZN(n1035) );
OR2_X1 U1031 ( .A1(G478), .A2(KEYINPUT15), .ZN(n1278) );
NAND3_X1 U1032 ( .A1(G478), .A2(n1037), .A3(KEYINPUT15), .ZN(n1277) );
NAND2_X1 U1033 ( .A1(n1198), .A2(n1093), .ZN(n1037) );
NAND2_X1 U1034 ( .A1(n1279), .A2(n1280), .ZN(n1093) );
NAND4_X1 U1035 ( .A1(n1281), .A2(n987), .A3(n1282), .A4(n1283), .ZN(n1280) );
AND2_X1 U1036 ( .A1(G234), .A2(G217), .ZN(n1283) );
NAND2_X1 U1037 ( .A1(n1284), .A2(n1285), .ZN(n1279) );
NAND3_X1 U1038 ( .A1(G234), .A2(n987), .A3(G217), .ZN(n1285) );
INV_X1 U1039 ( .A(G953), .ZN(n987) );
NAND2_X1 U1040 ( .A1(n1282), .A2(n1281), .ZN(n1284) );
NAND2_X1 U1041 ( .A1(n1286), .A2(n1287), .ZN(n1281) );
INV_X1 U1042 ( .A(n1288), .ZN(n1287) );
XOR2_X1 U1043 ( .A(n1289), .B(KEYINPUT24), .Z(n1286) );
XNOR2_X1 U1044 ( .A(n1290), .B(KEYINPUT28), .ZN(n1282) );
NAND2_X1 U1045 ( .A1(n1289), .A2(n1288), .ZN(n1290) );
XNOR2_X1 U1046 ( .A(n1291), .B(n1292), .ZN(n1288) );
XNOR2_X1 U1047 ( .A(KEYINPUT4), .B(n1194), .ZN(n1292) );
INV_X1 U1048 ( .A(G116), .ZN(n1194) );
XNOR2_X1 U1049 ( .A(n1293), .B(n1236), .ZN(n1291) );
INV_X1 U1050 ( .A(G107), .ZN(n1236) );
NAND2_X1 U1051 ( .A1(KEYINPUT57), .A2(n1184), .ZN(n1293) );
INV_X1 U1052 ( .A(G122), .ZN(n1184) );
XOR2_X1 U1053 ( .A(n1294), .B(n1295), .Z(n1289) );
XOR2_X1 U1054 ( .A(G128), .B(n1296), .Z(n1295) );
NOR2_X1 U1055 ( .A1(KEYINPUT39), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1056 ( .A(G143), .B(KEYINPUT52), .ZN(n1297) );
XNOR2_X1 U1057 ( .A(G134), .B(KEYINPUT49), .ZN(n1294) );
XNOR2_X1 U1058 ( .A(n1216), .B(KEYINPUT62), .ZN(n1198) );
INV_X1 U1059 ( .A(G902), .ZN(n1216) );
endmodule


