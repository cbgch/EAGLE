//Key = 0000110100101000110000110101011010101011011101000001101100110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335;

XOR2_X1 U732 ( .A(n1016), .B(n1017), .Z(G9) );
XOR2_X1 U733 ( .A(KEYINPUT21), .B(G107), .Z(n1017) );
NOR2_X1 U734 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR4_X1 U737 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1023) );
NAND3_X1 U738 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1020) );
NAND2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U741 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1034) );
NAND2_X1 U743 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U744 ( .A1(n1043), .A2(n1044), .A3(n1038), .ZN(n1042) );
NAND2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
INV_X1 U746 ( .A(n1047), .ZN(n1046) );
XNOR2_X1 U747 ( .A(n1048), .B(KEYINPUT47), .ZN(n1045) );
NAND2_X1 U748 ( .A1(n1036), .A2(n1049), .ZN(n1041) );
NAND3_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1024), .ZN(n1052) );
INV_X1 U751 ( .A(KEYINPUT56), .ZN(n1024) );
NAND3_X1 U752 ( .A1(n1037), .A2(n1054), .A3(n1055), .ZN(n1051) );
INV_X1 U753 ( .A(KEYINPUT10), .ZN(n1054) );
NAND3_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1038), .ZN(n1037) );
NAND2_X1 U755 ( .A1(n1043), .A2(n1058), .ZN(n1057) );
OR2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1039), .A2(n1061), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U759 ( .A1(KEYINPUT10), .A2(n1055), .ZN(n1063) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND3_X1 U761 ( .A1(n1066), .A2(n1043), .A3(n1067), .ZN(n1050) );
INV_X1 U762 ( .A(n1028), .ZN(n1032) );
AND3_X1 U763 ( .A1(n1029), .A2(n1030), .A3(n1068), .ZN(n1018) );
NAND4_X1 U764 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1029) );
NOR4_X1 U765 ( .A1(n1064), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XNOR2_X1 U766 ( .A(n1076), .B(n1077), .ZN(n1073) );
NAND2_X1 U767 ( .A1(KEYINPUT45), .A2(n1078), .ZN(n1076) );
XOR2_X1 U768 ( .A(n1079), .B(G478), .Z(n1071) );
XOR2_X1 U769 ( .A(n1080), .B(KEYINPUT62), .Z(n1070) );
XOR2_X1 U770 ( .A(n1081), .B(n1082), .Z(n1069) );
NAND2_X1 U771 ( .A1(KEYINPUT38), .A2(G475), .ZN(n1081) );
XOR2_X1 U772 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U774 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U775 ( .A1(n1030), .A2(n1089), .ZN(n1088) );
NAND2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U777 ( .A(KEYINPUT7), .B(n1092), .Z(n1091) );
OR3_X1 U778 ( .A1(n1093), .A2(KEYINPUT13), .A3(n1094), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1095), .A2(n1096), .ZN(n1085) );
INV_X1 U780 ( .A(KEYINPUT13), .ZN(n1096) );
NOR2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1095) );
XNOR2_X1 U782 ( .A(n1097), .B(n1098), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U784 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U785 ( .A(n1103), .B(KEYINPUT14), .Z(n1099) );
OR2_X1 U786 ( .A1(n1102), .A2(n1101), .ZN(n1103) );
XNOR2_X1 U787 ( .A(n1104), .B(n1105), .ZN(n1101) );
XOR2_X1 U788 ( .A(G134), .B(n1106), .Z(n1105) );
NOR2_X1 U789 ( .A1(G137), .A2(KEYINPUT1), .ZN(n1106) );
NAND2_X1 U790 ( .A1(KEYINPUT5), .A2(n1107), .ZN(n1104) );
NOR2_X1 U791 ( .A1(n1030), .A2(G900), .ZN(n1093) );
NAND2_X1 U792 ( .A1(G953), .A2(n1108), .ZN(n1083) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1109), .B(n1110), .Z(G69) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1030), .ZN(n1112) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
NAND2_X1 U799 ( .A1(G953), .A2(n1115), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1118), .B(n1119), .Z(n1116) );
XOR2_X1 U801 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U802 ( .A(KEYINPUT27), .B(n1122), .Z(n1118) );
NAND2_X1 U803 ( .A1(n1030), .A2(n1123), .ZN(n1109) );
NAND3_X1 U804 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
XNOR2_X1 U805 ( .A(n1127), .B(KEYINPUT28), .ZN(n1126) );
XOR2_X1 U806 ( .A(KEYINPUT52), .B(n1128), .Z(n1125) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(G66) );
XOR2_X1 U808 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND4_X1 U809 ( .A1(G217), .A2(n1022), .A3(n1133), .A4(n1134), .ZN(n1131) );
NAND2_X1 U810 ( .A1(G902), .A2(n1135), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1138), .ZN(n1136) );
INV_X1 U813 ( .A(KEYINPUT42), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1139), .ZN(G63) );
NOR3_X1 U815 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
NOR2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
AND2_X1 U817 ( .A1(n1022), .A2(G478), .ZN(n1144) );
INV_X1 U818 ( .A(n1145), .ZN(n1143) );
INV_X1 U819 ( .A(n1079), .ZN(n1141) );
XOR2_X1 U820 ( .A(KEYINPUT35), .B(n1146), .Z(n1140) );
NOR3_X1 U821 ( .A1(n1145), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR2_X1 U822 ( .A1(n1129), .A2(n1149), .ZN(G60) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1148), .ZN(n1150) );
XNOR2_X1 U825 ( .A(G475), .B(KEYINPUT44), .ZN(n1152) );
XOR2_X1 U826 ( .A(G104), .B(n1153), .Z(G6) );
NOR2_X1 U827 ( .A1(n1129), .A2(n1154), .ZN(G57) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U829 ( .A(KEYINPUT11), .B(n1157), .Z(n1156) );
NOR2_X1 U830 ( .A1(n1078), .A2(n1148), .ZN(n1157) );
INV_X1 U831 ( .A(G472), .ZN(n1078) );
XOR2_X1 U832 ( .A(n1158), .B(n1159), .Z(n1155) );
NOR2_X1 U833 ( .A1(n1129), .A2(n1160), .ZN(G54) );
XOR2_X1 U834 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U835 ( .A(n1163), .B(n1102), .Z(n1162) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1102) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1161) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1148), .ZN(n1167) );
INV_X1 U839 ( .A(G469), .ZN(n1168) );
NOR2_X1 U840 ( .A1(KEYINPUT53), .A2(n1169), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U842 ( .A1(KEYINPUT37), .A2(n1172), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1173), .B(G140), .Z(n1172) );
NAND2_X1 U844 ( .A1(KEYINPUT12), .A2(n1174), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1129), .A2(n1175), .ZN(G51) );
XNOR2_X1 U846 ( .A(n1176), .B(n1177), .ZN(n1175) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1148), .ZN(n1178) );
NAND2_X1 U849 ( .A1(G902), .A2(n1022), .ZN(n1148) );
NAND3_X1 U850 ( .A1(n1090), .A2(n1124), .A3(n1181), .ZN(n1022) );
NOR3_X1 U851 ( .A1(n1092), .A2(n1127), .A3(n1128), .ZN(n1181) );
AND3_X1 U852 ( .A1(n1038), .A2(n1059), .A3(n1182), .ZN(n1092) );
AND4_X1 U853 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1124) );
NOR3_X1 U854 ( .A1(n1187), .A2(n1153), .A3(n1016), .ZN(n1186) );
AND3_X1 U855 ( .A1(n1188), .A2(n1059), .A3(n1036), .ZN(n1016) );
AND3_X1 U856 ( .A1(n1036), .A2(n1188), .A3(n1060), .ZN(n1153) );
NAND3_X1 U857 ( .A1(n1039), .A2(n1047), .A3(n1188), .ZN(n1185) );
AND4_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1090) );
AND4_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
AND2_X1 U860 ( .A1(n1197), .A2(n1068), .ZN(n1129) );
INV_X1 U861 ( .A(G952), .ZN(n1068) );
XOR2_X1 U862 ( .A(n1030), .B(KEYINPUT54), .Z(n1197) );
XNOR2_X1 U863 ( .A(G146), .B(n1189), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1060), .A2(n1198), .A3(n1199), .ZN(n1189) );
XOR2_X1 U865 ( .A(G143), .B(n1200), .Z(G45) );
NOR2_X1 U866 ( .A1(KEYINPUT48), .A2(n1190), .ZN(n1200) );
NAND3_X1 U867 ( .A1(n1182), .A2(n1198), .A3(n1201), .ZN(n1190) );
XNOR2_X1 U868 ( .A(G140), .B(n1196), .ZN(G42) );
NAND3_X1 U869 ( .A1(n1038), .A2(n1055), .A3(n1202), .ZN(n1196) );
XNOR2_X1 U870 ( .A(G137), .B(n1195), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1038), .A2(n1039), .A3(n1199), .ZN(n1195) );
XOR2_X1 U872 ( .A(n1203), .B(n1204), .Z(G36) );
NAND4_X1 U873 ( .A1(n1205), .A2(n1038), .A3(n1206), .A4(n1047), .ZN(n1204) );
AND2_X1 U874 ( .A1(n1207), .A2(n1059), .ZN(n1206) );
XOR2_X1 U875 ( .A(n1208), .B(KEYINPUT34), .Z(n1205) );
NAND2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(G33) );
NAND2_X1 U877 ( .A1(n1211), .A2(n1107), .ZN(n1210) );
XOR2_X1 U878 ( .A(KEYINPUT17), .B(n1212), .Z(n1209) );
NOR2_X1 U879 ( .A1(n1107), .A2(n1211), .ZN(n1212) );
NAND2_X1 U880 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
OR2_X1 U881 ( .A1(n1191), .A2(KEYINPUT49), .ZN(n1214) );
NAND3_X1 U882 ( .A1(n1060), .A2(n1038), .A3(n1182), .ZN(n1191) );
INV_X1 U883 ( .A(n1075), .ZN(n1038) );
NAND4_X1 U884 ( .A1(n1060), .A2(n1075), .A3(n1182), .A4(KEYINPUT49), .ZN(n1213) );
NOR2_X1 U885 ( .A1(n1215), .A2(n1216), .ZN(n1182) );
NAND2_X1 U886 ( .A1(n1066), .A2(n1217), .ZN(n1075) );
INV_X1 U887 ( .A(G131), .ZN(n1107) );
NAND2_X1 U888 ( .A1(n1218), .A2(n1219), .ZN(G30) );
NAND2_X1 U889 ( .A1(G128), .A2(n1194), .ZN(n1219) );
XOR2_X1 U890 ( .A(n1220), .B(KEYINPUT46), .Z(n1218) );
OR2_X1 U891 ( .A1(n1194), .A2(G128), .ZN(n1220) );
NAND3_X1 U892 ( .A1(n1198), .A2(n1059), .A3(n1199), .ZN(n1194) );
NOR4_X1 U893 ( .A1(n1221), .A2(n1208), .A3(n1216), .A4(n1222), .ZN(n1199) );
INV_X1 U894 ( .A(n1207), .ZN(n1216) );
XOR2_X1 U895 ( .A(G101), .B(n1223), .Z(G3) );
NOR4_X1 U896 ( .A1(n1224), .A2(n1225), .A3(n1025), .A4(n1215), .ZN(n1223) );
NAND2_X1 U897 ( .A1(n1055), .A2(n1047), .ZN(n1215) );
XNOR2_X1 U898 ( .A(n1198), .B(KEYINPUT61), .ZN(n1225) );
AND2_X1 U899 ( .A1(n1226), .A2(n1028), .ZN(n1224) );
XNOR2_X1 U900 ( .A(G125), .B(n1193), .ZN(G27) );
NAND2_X1 U901 ( .A1(n1202), .A2(n1053), .ZN(n1193) );
AND3_X1 U902 ( .A1(n1048), .A2(n1207), .A3(n1060), .ZN(n1202) );
NAND2_X1 U903 ( .A1(n1028), .A2(n1227), .ZN(n1207) );
NAND2_X1 U904 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U905 ( .A(G900), .ZN(n1229) );
XNOR2_X1 U906 ( .A(G122), .B(n1183), .ZN(G24) );
NAND3_X1 U907 ( .A1(n1230), .A2(n1036), .A3(n1201), .ZN(n1183) );
AND2_X1 U908 ( .A1(n1231), .A2(n1232), .ZN(n1201) );
XOR2_X1 U909 ( .A(KEYINPUT31), .B(n1233), .Z(n1231) );
INV_X1 U910 ( .A(n1026), .ZN(n1036) );
XOR2_X1 U911 ( .A(n1234), .B(G119), .Z(G21) );
NAND2_X1 U912 ( .A1(KEYINPUT63), .A2(n1184), .ZN(n1234) );
NAND4_X1 U913 ( .A1(n1235), .A2(n1230), .A3(n1039), .A4(n1074), .ZN(n1184) );
XOR2_X1 U914 ( .A(G116), .B(n1187), .Z(G18) );
AND3_X1 U915 ( .A1(n1047), .A2(n1059), .A3(n1230), .ZN(n1187) );
NAND2_X1 U916 ( .A1(n1236), .A2(n1237), .ZN(n1059) );
OR2_X1 U917 ( .A1(n1025), .A2(KEYINPUT16), .ZN(n1237) );
NAND3_X1 U918 ( .A1(n1233), .A2(n1238), .A3(KEYINPUT16), .ZN(n1236) );
XOR2_X1 U919 ( .A(G113), .B(n1128), .Z(G15) );
AND3_X1 U920 ( .A1(n1060), .A2(n1047), .A3(n1230), .ZN(n1128) );
AND2_X1 U921 ( .A1(n1053), .A2(n1239), .ZN(n1230) );
INV_X1 U922 ( .A(n1027), .ZN(n1053) );
NAND2_X1 U923 ( .A1(n1198), .A2(n1043), .ZN(n1027) );
NAND2_X1 U924 ( .A1(n1240), .A2(n1241), .ZN(n1043) );
OR2_X1 U925 ( .A1(n1208), .A2(KEYINPUT30), .ZN(n1241) );
INV_X1 U926 ( .A(n1055), .ZN(n1208) );
NAND3_X1 U927 ( .A1(n1065), .A2(n1242), .A3(KEYINPUT30), .ZN(n1240) );
NAND2_X1 U928 ( .A1(n1243), .A2(n1244), .ZN(n1047) );
OR2_X1 U929 ( .A1(n1026), .A2(KEYINPUT55), .ZN(n1244) );
NAND2_X1 U930 ( .A1(n1222), .A2(n1221), .ZN(n1026) );
INV_X1 U931 ( .A(n1235), .ZN(n1221) );
NAND3_X1 U932 ( .A1(n1222), .A2(n1235), .A3(KEYINPUT55), .ZN(n1243) );
NOR2_X1 U933 ( .A1(n1238), .A2(n1233), .ZN(n1060) );
INV_X1 U934 ( .A(n1245), .ZN(n1233) );
XOR2_X1 U935 ( .A(G110), .B(n1127), .Z(G12) );
AND3_X1 U936 ( .A1(n1188), .A2(n1039), .A3(n1048), .ZN(n1127) );
NOR2_X1 U937 ( .A1(n1235), .A2(n1222), .ZN(n1048) );
INV_X1 U938 ( .A(n1074), .ZN(n1222) );
NAND3_X1 U939 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1074) );
OR2_X1 U940 ( .A1(n1249), .A2(n1132), .ZN(n1248) );
NAND3_X1 U941 ( .A1(n1132), .A2(n1249), .A3(n1137), .ZN(n1247) );
NAND2_X1 U942 ( .A1(G217), .A2(n1138), .ZN(n1249) );
INV_X1 U943 ( .A(G234), .ZN(n1138) );
XNOR2_X1 U944 ( .A(n1250), .B(n1251), .ZN(n1132) );
XOR2_X1 U945 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U946 ( .A(G146), .B(G119), .Z(n1253) );
XOR2_X1 U947 ( .A(KEYINPUT57), .B(KEYINPUT4), .Z(n1252) );
XOR2_X1 U948 ( .A(n1254), .B(n1255), .Z(n1250) );
XOR2_X1 U949 ( .A(n1256), .B(n1257), .Z(n1255) );
AND3_X1 U950 ( .A1(G234), .A2(n1030), .A3(G221), .ZN(n1257) );
NOR2_X1 U951 ( .A1(KEYINPUT3), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U952 ( .A(G137), .B(KEYINPUT6), .ZN(n1258) );
XNOR2_X1 U953 ( .A(n1259), .B(n1260), .ZN(n1254) );
NOR2_X1 U954 ( .A1(G125), .A2(KEYINPUT33), .ZN(n1260) );
NAND2_X1 U955 ( .A1(G902), .A2(G217), .ZN(n1246) );
XOR2_X1 U956 ( .A(n1077), .B(n1261), .Z(n1235) );
NOR2_X1 U957 ( .A1(KEYINPUT9), .A2(n1262), .ZN(n1261) );
XOR2_X1 U958 ( .A(KEYINPUT50), .B(G472), .Z(n1262) );
NAND2_X1 U959 ( .A1(n1263), .A2(n1137), .ZN(n1077) );
XOR2_X1 U960 ( .A(n1264), .B(n1158), .Z(n1263) );
XOR2_X1 U961 ( .A(n1265), .B(n1266), .Z(n1158) );
XOR2_X1 U962 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U963 ( .A1(G210), .A2(n1269), .ZN(n1268) );
NAND2_X1 U964 ( .A1(KEYINPUT58), .A2(n1270), .ZN(n1267) );
XOR2_X1 U965 ( .A(n1271), .B(n1272), .Z(n1265) );
NAND2_X1 U966 ( .A1(KEYINPUT32), .A2(n1273), .ZN(n1264) );
XOR2_X1 U967 ( .A(KEYINPUT60), .B(n1159), .Z(n1273) );
INV_X1 U968 ( .A(n1025), .ZN(n1039) );
NAND2_X1 U969 ( .A1(n1238), .A2(n1245), .ZN(n1025) );
NAND3_X1 U970 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1245) );
OR2_X1 U971 ( .A1(n1079), .A2(KEYINPUT59), .ZN(n1276) );
NAND4_X1 U972 ( .A1(KEYINPUT25), .A2(n1079), .A3(KEYINPUT59), .A4(n1147), .ZN(n1275) );
INV_X1 U973 ( .A(G478), .ZN(n1147) );
NAND2_X1 U974 ( .A1(G478), .A2(n1277), .ZN(n1274) );
NAND2_X1 U975 ( .A1(KEYINPUT25), .A2(n1079), .ZN(n1277) );
NAND2_X1 U976 ( .A1(n1137), .A2(n1145), .ZN(n1079) );
NAND2_X1 U977 ( .A1(n1278), .A2(n1279), .ZN(n1145) );
NAND2_X1 U978 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U979 ( .A(n1282), .B(KEYINPUT24), .Z(n1278) );
OR2_X1 U980 ( .A1(n1281), .A2(n1280), .ZN(n1282) );
XNOR2_X1 U981 ( .A(n1283), .B(n1284), .ZN(n1280) );
XOR2_X1 U982 ( .A(G143), .B(G134), .Z(n1284) );
XOR2_X1 U983 ( .A(n1285), .B(G128), .Z(n1283) );
NAND2_X1 U984 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
OR2_X1 U985 ( .A1(n1288), .A2(G107), .ZN(n1287) );
XOR2_X1 U986 ( .A(n1289), .B(KEYINPUT15), .Z(n1286) );
NAND2_X1 U987 ( .A1(G107), .A2(n1288), .ZN(n1289) );
XNOR2_X1 U988 ( .A(n1290), .B(n1291), .ZN(n1288) );
XOR2_X1 U989 ( .A(KEYINPUT2), .B(G122), .Z(n1291) );
INV_X1 U990 ( .A(G116), .ZN(n1290) );
NAND3_X1 U991 ( .A1(G217), .A2(n1030), .A3(G234), .ZN(n1281) );
INV_X1 U992 ( .A(n1232), .ZN(n1238) );
XOR2_X1 U993 ( .A(n1082), .B(G475), .Z(n1232) );
NOR2_X1 U994 ( .A1(n1151), .A2(G902), .ZN(n1082) );
XNOR2_X1 U995 ( .A(n1292), .B(n1293), .ZN(n1151) );
XOR2_X1 U996 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U997 ( .A(G122), .B(G113), .Z(n1295) );
XOR2_X1 U998 ( .A(KEYINPUT29), .B(G131), .Z(n1294) );
XOR2_X1 U999 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U1000 ( .A(G104), .B(n1298), .Z(n1297) );
AND3_X1 U1001 ( .A1(G214), .A2(n1299), .A3(n1269), .ZN(n1298) );
NOR2_X1 U1002 ( .A1(G953), .A2(G237), .ZN(n1269) );
INV_X1 U1003 ( .A(KEYINPUT19), .ZN(n1299) );
XOR2_X1 U1004 ( .A(n1098), .B(n1165), .Z(n1296) );
XOR2_X1 U1005 ( .A(G125), .B(G140), .Z(n1098) );
AND3_X1 U1006 ( .A1(n1055), .A2(n1239), .A3(n1198), .ZN(n1188) );
NOR2_X1 U1007 ( .A1(n1066), .A2(n1067), .ZN(n1198) );
INV_X1 U1008 ( .A(n1217), .ZN(n1067) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1300), .ZN(n1217) );
XNOR2_X1 U1010 ( .A(n1301), .B(n1180), .ZN(n1066) );
NAND2_X1 U1011 ( .A1(G210), .A2(n1300), .ZN(n1180) );
NAND2_X1 U1012 ( .A1(n1137), .A2(n1302), .ZN(n1300) );
INV_X1 U1013 ( .A(G237), .ZN(n1302) );
NAND2_X1 U1014 ( .A1(n1303), .A2(n1137), .ZN(n1301) );
XNOR2_X1 U1015 ( .A(n1304), .B(n1179), .ZN(n1303) );
XNOR2_X1 U1016 ( .A(n1305), .B(n1122), .ZN(n1179) );
XOR2_X1 U1017 ( .A(G110), .B(G122), .Z(n1122) );
NAND3_X1 U1018 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1305) );
NAND2_X1 U1019 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1020 ( .A1(n1311), .A2(KEYINPUT41), .ZN(n1310) );
XNOR2_X1 U1021 ( .A(n1120), .B(KEYINPUT43), .ZN(n1311) );
NAND3_X1 U1022 ( .A1(KEYINPUT41), .A2(n1121), .A3(n1120), .ZN(n1307) );
INV_X1 U1023 ( .A(n1309), .ZN(n1121) );
XOR2_X1 U1024 ( .A(n1312), .B(n1313), .Z(n1309) );
XOR2_X1 U1025 ( .A(G107), .B(G101), .Z(n1313) );
NAND2_X1 U1026 ( .A1(KEYINPUT39), .A2(n1314), .ZN(n1312) );
INV_X1 U1027 ( .A(G104), .ZN(n1314) );
OR2_X1 U1028 ( .A1(n1120), .A2(KEYINPUT41), .ZN(n1306) );
XNOR2_X1 U1029 ( .A(n1315), .B(n1272), .ZN(n1120) );
XOR2_X1 U1030 ( .A(G113), .B(n1316), .Z(n1272) );
XOR2_X1 U1031 ( .A(KEYINPUT40), .B(G116), .Z(n1316) );
NAND2_X1 U1032 ( .A1(KEYINPUT36), .A2(n1270), .ZN(n1315) );
INV_X1 U1033 ( .A(G119), .ZN(n1270) );
NAND2_X1 U1034 ( .A1(KEYINPUT51), .A2(n1176), .ZN(n1304) );
XOR2_X1 U1035 ( .A(n1159), .B(n1317), .Z(n1176) );
XOR2_X1 U1036 ( .A(G125), .B(n1318), .Z(n1317) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1114), .ZN(n1318) );
INV_X1 U1038 ( .A(G224), .ZN(n1114) );
XNOR2_X1 U1039 ( .A(n1164), .B(n1319), .ZN(n1159) );
NOR2_X1 U1040 ( .A1(KEYINPUT18), .A2(n1165), .ZN(n1319) );
INV_X1 U1041 ( .A(G128), .ZN(n1164) );
NAND2_X1 U1042 ( .A1(n1226), .A2(n1028), .ZN(n1239) );
NAND3_X1 U1043 ( .A1(n1320), .A2(n1030), .A3(G952), .ZN(n1028) );
NAND2_X1 U1044 ( .A1(n1228), .A2(n1115), .ZN(n1226) );
INV_X1 U1045 ( .A(G898), .ZN(n1115) );
AND3_X1 U1046 ( .A1(n1321), .A2(n1320), .A3(G953), .ZN(n1228) );
NAND2_X1 U1047 ( .A1(G237), .A2(G234), .ZN(n1320) );
XOR2_X1 U1048 ( .A(KEYINPUT26), .B(G902), .Z(n1321) );
NOR2_X1 U1049 ( .A1(n1065), .A2(n1064), .ZN(n1055) );
INV_X1 U1050 ( .A(n1242), .ZN(n1064) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1322), .ZN(n1242) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1137), .ZN(n1322) );
XOR2_X1 U1053 ( .A(n1080), .B(KEYINPUT20), .Z(n1065) );
XOR2_X1 U1054 ( .A(n1323), .B(G469), .Z(n1080) );
NAND2_X1 U1055 ( .A1(n1324), .A2(n1137), .ZN(n1323) );
INV_X1 U1056 ( .A(G902), .ZN(n1137) );
XOR2_X1 U1057 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1058 ( .A(n1163), .B(n1259), .ZN(n1326) );
XNOR2_X1 U1059 ( .A(n1174), .B(n1327), .ZN(n1259) );
XOR2_X1 U1060 ( .A(G140), .B(G128), .Z(n1327) );
INV_X1 U1061 ( .A(G110), .ZN(n1174) );
XNOR2_X1 U1062 ( .A(n1271), .B(n1328), .ZN(n1163) );
XOR2_X1 U1063 ( .A(G107), .B(n1329), .Z(n1328) );
NOR2_X1 U1064 ( .A1(G104), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1065 ( .A(KEYINPUT22), .B(KEYINPUT0), .ZN(n1330) );
XOR2_X1 U1066 ( .A(n1331), .B(n1332), .Z(n1271) );
XOR2_X1 U1067 ( .A(G137), .B(G131), .Z(n1332) );
XOR2_X1 U1068 ( .A(n1333), .B(G101), .Z(n1331) );
NAND2_X1 U1069 ( .A1(KEYINPUT23), .A2(n1203), .ZN(n1333) );
INV_X1 U1070 ( .A(G134), .ZN(n1203) );
XOR2_X1 U1071 ( .A(n1334), .B(n1170), .Z(n1325) );
NAND2_X1 U1072 ( .A1(n1335), .A2(G227), .ZN(n1170) );
XOR2_X1 U1073 ( .A(n1030), .B(KEYINPUT8), .Z(n1335) );
INV_X1 U1074 ( .A(G953), .ZN(n1030) );
INV_X1 U1075 ( .A(n1165), .ZN(n1334) );
XNOR2_X1 U1076 ( .A(G143), .B(G146), .ZN(n1165) );
endmodule


