//Key = 1010110111100101010111011000111010110110111001000010000010111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;

XOR2_X1 U743 ( .A(n1016), .B(n1017), .Z(G9) );
NOR2_X1 U744 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR3_X1 U745 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NAND3_X1 U746 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1020) );
NAND2_X1 U747 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U748 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U749 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1035), .A2(n1036), .ZN(n1028) );
NAND3_X1 U752 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U753 ( .A1(n1030), .A2(n1040), .ZN(n1039) );
NAND2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U756 ( .A1(n1032), .A2(n1045), .ZN(n1038) );
NAND2_X1 U757 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
OR2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1046) );
NAND2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U762 ( .A1(KEYINPUT7), .A2(n1056), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NAND4_X1 U764 ( .A1(n1056), .A2(n1059), .A3(n1052), .A4(n1060), .ZN(n1037) );
INV_X1 U765 ( .A(KEYINPUT7), .ZN(n1059) );
INV_X1 U766 ( .A(n1061), .ZN(n1026) );
NOR3_X1 U767 ( .A1(n1062), .A2(G953), .A3(n1063), .ZN(n1018) );
INV_X1 U768 ( .A(n1023), .ZN(n1063) );
NAND4_X1 U769 ( .A1(n1043), .A2(n1048), .A3(n1064), .A4(n1065), .ZN(n1023) );
NOR4_X1 U770 ( .A1(n1066), .A2(n1044), .A3(n1067), .A4(n1068), .ZN(n1065) );
XOR2_X1 U771 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U772 ( .A1(KEYINPUT3), .A2(n1071), .ZN(n1070) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1067) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1064) );
XOR2_X1 U775 ( .A(n1076), .B(n1077), .Z(n1074) );
XOR2_X1 U776 ( .A(KEYINPUT31), .B(n1078), .Z(n1077) );
NOR2_X1 U777 ( .A1(G478), .A2(n1079), .ZN(n1078) );
XOR2_X1 U778 ( .A(KEYINPUT37), .B(KEYINPUT0), .Z(n1079) );
XOR2_X1 U779 ( .A(n1021), .B(KEYINPUT58), .Z(n1062) );
INV_X1 U780 ( .A(G952), .ZN(n1021) );
XOR2_X1 U781 ( .A(n1080), .B(n1081), .Z(G72) );
NOR3_X1 U782 ( .A1(n1024), .A2(KEYINPUT62), .A3(n1082), .ZN(n1081) );
AND2_X1 U783 ( .A1(G227), .A2(G900), .ZN(n1082) );
NAND2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1085), .A2(n1024), .ZN(n1084) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND3_X1 U787 ( .A1(n1087), .A2(G900), .A3(G953), .ZN(n1083) );
AND2_X1 U788 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U789 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U790 ( .A(KEYINPUT13), .B(n1092), .Z(n1088) );
NOR2_X1 U791 ( .A1(n1090), .A2(n1091), .ZN(n1092) );
XNOR2_X1 U792 ( .A(n1093), .B(n1094), .ZN(n1091) );
XNOR2_X1 U793 ( .A(n1095), .B(KEYINPUT46), .ZN(n1094) );
NAND2_X1 U794 ( .A1(KEYINPUT4), .A2(n1096), .ZN(n1095) );
XOR2_X1 U795 ( .A(n1097), .B(n1098), .Z(n1093) );
AND2_X1 U796 ( .A1(n1099), .A2(n1100), .ZN(n1090) );
NAND2_X1 U797 ( .A1(G140), .A2(G125), .ZN(n1100) );
NAND2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
INV_X1 U799 ( .A(G140), .ZN(n1102) );
XOR2_X1 U800 ( .A(n1103), .B(KEYINPUT47), .Z(n1101) );
NAND2_X1 U801 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND2_X1 U802 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U803 ( .A1(G953), .A2(n1108), .ZN(n1107) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1108) );
NAND2_X1 U805 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
INV_X1 U806 ( .A(n1106), .ZN(n1110) );
NOR2_X1 U807 ( .A1(KEYINPUT33), .A2(n1111), .ZN(n1106) );
XOR2_X1 U808 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U809 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U810 ( .A(KEYINPUT36), .B(G953), .Z(n1115) );
INV_X1 U811 ( .A(n1116), .ZN(n1114) );
NAND2_X1 U812 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
XOR2_X1 U813 ( .A(n1119), .B(n1120), .Z(n1117) );
NAND3_X1 U814 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1119) );
NAND2_X1 U815 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
INV_X1 U816 ( .A(KEYINPUT18), .ZN(n1125) );
NAND2_X1 U817 ( .A1(KEYINPUT18), .A2(n1126), .ZN(n1121) );
NAND2_X1 U818 ( .A1(n1118), .A2(n1127), .ZN(n1109) );
OR2_X1 U819 ( .A1(n1024), .A2(G224), .ZN(n1127) );
NOR2_X1 U820 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U821 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U822 ( .A1(n1132), .A2(n1072), .ZN(n1130) );
INV_X1 U823 ( .A(n1133), .ZN(n1072) );
NOR2_X1 U824 ( .A1(n1128), .A2(n1134), .ZN(G63) );
XOR2_X1 U825 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U826 ( .A1(KEYINPUT21), .A2(n1137), .ZN(n1136) );
NAND2_X1 U827 ( .A1(n1132), .A2(G478), .ZN(n1135) );
NOR2_X1 U828 ( .A1(n1128), .A2(n1138), .ZN(G60) );
XNOR2_X1 U829 ( .A(n1139), .B(n1140), .ZN(n1138) );
NAND2_X1 U830 ( .A1(n1132), .A2(G475), .ZN(n1139) );
NAND2_X1 U831 ( .A1(n1141), .A2(n1142), .ZN(G6) );
NAND2_X1 U832 ( .A1(G104), .A2(n1143), .ZN(n1142) );
XOR2_X1 U833 ( .A(n1144), .B(KEYINPUT26), .Z(n1141) );
OR2_X1 U834 ( .A1(n1143), .A2(G104), .ZN(n1144) );
NAND3_X1 U835 ( .A1(n1145), .A2(n1035), .A3(n1050), .ZN(n1143) );
NOR2_X1 U836 ( .A1(n1128), .A2(n1146), .ZN(G57) );
XOR2_X1 U837 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U838 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U839 ( .A(n1151), .B(G101), .Z(n1147) );
NAND3_X1 U840 ( .A1(G902), .A2(n1152), .A3(G472), .ZN(n1151) );
XOR2_X1 U841 ( .A(KEYINPUT19), .B(n1153), .Z(n1152) );
NOR2_X1 U842 ( .A1(n1128), .A2(n1154), .ZN(G54) );
XOR2_X1 U843 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U844 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U845 ( .A1(KEYINPUT8), .A2(n1159), .ZN(n1158) );
NAND2_X1 U846 ( .A1(n1132), .A2(G469), .ZN(n1157) );
INV_X1 U847 ( .A(n1160), .ZN(n1132) );
NOR2_X1 U848 ( .A1(n1128), .A2(n1161), .ZN(G51) );
XOR2_X1 U849 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U850 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR3_X1 U851 ( .A1(n1160), .A2(KEYINPUT11), .A3(n1166), .ZN(n1164) );
NAND2_X1 U852 ( .A1(G902), .A2(n1022), .ZN(n1160) );
INV_X1 U853 ( .A(n1153), .ZN(n1022) );
NOR2_X1 U854 ( .A1(n1116), .A2(n1086), .ZN(n1153) );
NAND4_X1 U855 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1086) );
NOR4_X1 U856 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170) );
INV_X1 U857 ( .A(n1175), .ZN(n1173) );
NAND2_X1 U858 ( .A1(n1176), .A2(n1177), .ZN(n1169) );
XNOR2_X1 U859 ( .A(n1178), .B(KEYINPUT61), .ZN(n1176) );
NAND2_X1 U860 ( .A1(n1179), .A2(n1180), .ZN(n1167) );
NAND2_X1 U861 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U862 ( .A1(n1050), .A2(n1183), .ZN(n1182) );
NAND2_X1 U863 ( .A1(n1184), .A2(n1051), .ZN(n1181) );
INV_X1 U864 ( .A(n1185), .ZN(n1179) );
NAND2_X1 U865 ( .A1(n1186), .A2(n1187), .ZN(n1116) );
NOR4_X1 U866 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR4_X1 U867 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1186) );
NOR2_X1 U868 ( .A1(n1196), .A2(n1041), .ZN(n1195) );
INV_X1 U869 ( .A(n1177), .ZN(n1041) );
XNOR2_X1 U870 ( .A(n1197), .B(KEYINPUT6), .ZN(n1196) );
NOR4_X1 U871 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1194) );
NOR2_X1 U872 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
INV_X1 U873 ( .A(KEYINPUT63), .ZN(n1203) );
NOR3_X1 U874 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1202) );
NOR2_X1 U875 ( .A1(KEYINPUT63), .A2(n1145), .ZN(n1198) );
INV_X1 U876 ( .A(n1017), .ZN(n1193) );
NAND3_X1 U877 ( .A1(n1051), .A2(n1035), .A3(n1145), .ZN(n1017) );
INV_X1 U878 ( .A(n1200), .ZN(n1035) );
INV_X1 U879 ( .A(n1207), .ZN(n1192) );
NOR2_X1 U880 ( .A1(n1208), .A2(n1209), .ZN(n1162) );
NOR2_X1 U881 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U882 ( .A(n1212), .B(KEYINPUT59), .Z(n1211) );
NOR2_X1 U883 ( .A1(n1213), .A2(n1214), .ZN(n1208) );
XOR2_X1 U884 ( .A(n1212), .B(KEYINPUT1), .Z(n1214) );
NOR2_X1 U885 ( .A1(n1024), .A2(G952), .ZN(n1128) );
XOR2_X1 U886 ( .A(G146), .B(n1174), .Z(G48) );
AND3_X1 U887 ( .A1(n1177), .A2(n1050), .A3(n1215), .ZN(n1174) );
XOR2_X1 U888 ( .A(n1216), .B(n1175), .Z(G45) );
NAND4_X1 U889 ( .A1(n1217), .A2(n1184), .A3(n1177), .A4(n1218), .ZN(n1175) );
NOR3_X1 U890 ( .A1(n1206), .A2(n1219), .A3(n1220), .ZN(n1218) );
XOR2_X1 U891 ( .A(n1221), .B(n1222), .Z(G42) );
XOR2_X1 U892 ( .A(KEYINPUT55), .B(G140), .Z(n1222) );
NOR4_X1 U893 ( .A1(KEYINPUT53), .A2(n1034), .A3(n1201), .A4(n1185), .ZN(n1221) );
XOR2_X1 U894 ( .A(n1096), .B(n1223), .Z(G39) );
NAND2_X1 U895 ( .A1(KEYINPUT23), .A2(n1172), .ZN(n1223) );
AND3_X1 U896 ( .A1(n1032), .A2(n1052), .A3(n1215), .ZN(n1172) );
XNOR2_X1 U897 ( .A(G134), .B(n1224), .ZN(G36) );
NAND4_X1 U898 ( .A1(n1225), .A2(n1226), .A3(n1051), .A4(n1227), .ZN(n1224) );
NOR2_X1 U899 ( .A1(n1033), .A2(n1060), .ZN(n1227) );
INV_X1 U900 ( .A(n1032), .ZN(n1060) );
XOR2_X1 U901 ( .A(KEYINPUT43), .B(n1056), .Z(n1225) );
XNOR2_X1 U902 ( .A(n1171), .B(n1228), .ZN(G33) );
XOR2_X1 U903 ( .A(KEYINPUT56), .B(G131), .Z(n1228) );
NOR3_X1 U904 ( .A1(n1201), .A2(n1033), .A3(n1185), .ZN(n1171) );
NAND3_X1 U905 ( .A1(n1056), .A2(n1226), .A3(n1032), .ZN(n1185) );
NOR2_X1 U906 ( .A1(n1229), .A2(n1230), .ZN(n1032) );
XOR2_X1 U907 ( .A(KEYINPUT50), .B(n1043), .Z(n1230) );
XOR2_X1 U908 ( .A(n1231), .B(n1232), .Z(G30) );
NAND2_X1 U909 ( .A1(n1178), .A2(n1177), .ZN(n1232) );
AND2_X1 U910 ( .A1(n1215), .A2(n1051), .ZN(n1178) );
NOR4_X1 U911 ( .A1(n1206), .A2(n1233), .A3(n1219), .A4(n1234), .ZN(n1215) );
XOR2_X1 U912 ( .A(n1235), .B(n1207), .Z(G3) );
NAND3_X1 U913 ( .A1(n1052), .A2(n1145), .A3(n1184), .ZN(n1207) );
INV_X1 U914 ( .A(n1033), .ZN(n1184) );
XOR2_X1 U915 ( .A(n1103), .B(n1168), .Z(G27) );
NAND3_X1 U916 ( .A1(n1177), .A2(n1050), .A3(n1236), .ZN(n1168) );
NOR3_X1 U917 ( .A1(n1034), .A2(n1219), .A3(n1237), .ZN(n1236) );
INV_X1 U918 ( .A(n1226), .ZN(n1219) );
NAND2_X1 U919 ( .A1(n1238), .A2(n1061), .ZN(n1226) );
XOR2_X1 U920 ( .A(KEYINPUT9), .B(n1239), .Z(n1238) );
NOR3_X1 U921 ( .A1(n1240), .A2(G900), .A3(n1024), .ZN(n1239) );
INV_X1 U922 ( .A(n1183), .ZN(n1034) );
XNOR2_X1 U923 ( .A(G122), .B(n1241), .ZN(G24) );
NAND2_X1 U924 ( .A1(n1197), .A2(n1177), .ZN(n1241) );
AND3_X1 U925 ( .A1(n1217), .A2(n1048), .A3(n1242), .ZN(n1197) );
NOR3_X1 U926 ( .A1(n1200), .A2(n1243), .A3(n1220), .ZN(n1242) );
NAND2_X1 U927 ( .A1(n1234), .A2(n1233), .ZN(n1200) );
XOR2_X1 U928 ( .A(n1244), .B(n1245), .Z(G21) );
NAND2_X1 U929 ( .A1(KEYINPUT28), .A2(n1191), .ZN(n1245) );
AND3_X1 U930 ( .A1(n1177), .A2(n1030), .A3(n1246), .ZN(n1191) );
NOR3_X1 U931 ( .A1(n1233), .A2(n1243), .A3(n1234), .ZN(n1246) );
AND2_X1 U932 ( .A1(n1052), .A2(n1048), .ZN(n1030) );
INV_X1 U933 ( .A(n1237), .ZN(n1048) );
NAND2_X1 U934 ( .A1(n1247), .A2(n1248), .ZN(G18) );
NAND2_X1 U935 ( .A1(n1190), .A2(n1249), .ZN(n1248) );
XOR2_X1 U936 ( .A(KEYINPUT35), .B(n1250), .Z(n1247) );
NOR2_X1 U937 ( .A1(n1190), .A2(n1249), .ZN(n1250) );
INV_X1 U938 ( .A(G116), .ZN(n1249) );
AND3_X1 U939 ( .A1(n1251), .A2(n1051), .A3(n1177), .ZN(n1190) );
XOR2_X1 U940 ( .A(n1205), .B(KEYINPUT17), .Z(n1177) );
NOR2_X1 U941 ( .A1(n1217), .A2(n1220), .ZN(n1051) );
XNOR2_X1 U942 ( .A(n1189), .B(n1252), .ZN(G15) );
XNOR2_X1 U943 ( .A(G113), .B(KEYINPUT39), .ZN(n1252) );
AND3_X1 U944 ( .A1(n1050), .A2(n1253), .A3(n1251), .ZN(n1189) );
NOR3_X1 U945 ( .A1(n1237), .A2(n1243), .A3(n1033), .ZN(n1251) );
NAND2_X1 U946 ( .A1(n1234), .A2(n1254), .ZN(n1033) );
NAND2_X1 U947 ( .A1(n1058), .A2(n1255), .ZN(n1237) );
INV_X1 U948 ( .A(n1201), .ZN(n1050) );
NAND2_X1 U949 ( .A1(n1217), .A2(n1220), .ZN(n1201) );
XOR2_X1 U950 ( .A(G110), .B(n1188), .Z(G12) );
AND3_X1 U951 ( .A1(n1052), .A2(n1145), .A3(n1183), .ZN(n1188) );
NOR2_X1 U952 ( .A1(n1254), .A2(n1234), .ZN(n1183) );
NOR2_X1 U953 ( .A1(n1256), .A2(n1066), .ZN(n1234) );
NOR2_X1 U954 ( .A1(n1133), .A2(n1257), .ZN(n1066) );
AND2_X1 U955 ( .A1(n1258), .A2(n1257), .ZN(n1256) );
INV_X1 U956 ( .A(n1073), .ZN(n1257) );
NAND2_X1 U957 ( .A1(n1259), .A2(n1131), .ZN(n1073) );
XNOR2_X1 U958 ( .A(n1260), .B(n1261), .ZN(n1131) );
XNOR2_X1 U959 ( .A(n1262), .B(n1263), .ZN(n1261) );
NAND2_X1 U960 ( .A1(KEYINPUT20), .A2(n1264), .ZN(n1262) );
XOR2_X1 U961 ( .A(n1096), .B(n1265), .Z(n1264) );
NAND2_X1 U962 ( .A1(n1266), .A2(G221), .ZN(n1265) );
XOR2_X1 U963 ( .A(n1267), .B(n1268), .Z(n1260) );
NOR2_X1 U964 ( .A1(KEYINPUT27), .A2(n1103), .ZN(n1268) );
XOR2_X1 U965 ( .A(n1244), .B(G146), .Z(n1267) );
XOR2_X1 U966 ( .A(KEYINPUT10), .B(G902), .Z(n1259) );
XOR2_X1 U967 ( .A(n1133), .B(KEYINPUT57), .Z(n1258) );
NAND2_X1 U968 ( .A1(G217), .A2(n1269), .ZN(n1133) );
INV_X1 U969 ( .A(n1233), .ZN(n1254) );
XOR2_X1 U970 ( .A(n1069), .B(n1071), .Z(n1233) );
XOR2_X1 U971 ( .A(G472), .B(KEYINPUT16), .Z(n1071) );
NAND2_X1 U972 ( .A1(n1270), .A2(n1271), .ZN(n1069) );
XOR2_X1 U973 ( .A(n1149), .B(n1272), .Z(n1270) );
XNOR2_X1 U974 ( .A(n1273), .B(n1274), .ZN(n1272) );
NOR2_X1 U975 ( .A1(KEYINPUT22), .A2(n1150), .ZN(n1274) );
XOR2_X1 U976 ( .A(n1275), .B(n1276), .Z(n1150) );
NAND2_X1 U977 ( .A1(KEYINPUT29), .A2(n1235), .ZN(n1273) );
INV_X1 U978 ( .A(G101), .ZN(n1235) );
XNOR2_X1 U979 ( .A(n1277), .B(n1278), .ZN(n1149) );
XOR2_X1 U980 ( .A(G113), .B(n1279), .Z(n1278) );
NOR2_X1 U981 ( .A1(KEYINPUT48), .A2(n1280), .ZN(n1279) );
NOR2_X1 U982 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NOR2_X1 U983 ( .A1(G119), .A2(n1283), .ZN(n1281) );
XOR2_X1 U984 ( .A(KEYINPUT38), .B(G116), .Z(n1283) );
NAND2_X1 U985 ( .A1(n1284), .A2(G210), .ZN(n1277) );
NOR3_X1 U986 ( .A1(n1205), .A2(n1243), .A3(n1206), .ZN(n1145) );
INV_X1 U987 ( .A(n1056), .ZN(n1206) );
NOR2_X1 U988 ( .A1(n1058), .A2(n1057), .ZN(n1056) );
INV_X1 U989 ( .A(n1255), .ZN(n1057) );
NAND2_X1 U990 ( .A1(G221), .A2(n1269), .ZN(n1255) );
NAND2_X1 U991 ( .A1(G234), .A2(n1271), .ZN(n1269) );
XOR2_X1 U992 ( .A(n1285), .B(G469), .Z(n1058) );
NAND2_X1 U993 ( .A1(n1286), .A2(n1271), .ZN(n1285) );
XOR2_X1 U994 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U995 ( .A(n1155), .B(n1159), .Z(n1288) );
NAND2_X1 U996 ( .A1(n1289), .A2(n1290), .ZN(n1159) );
NAND2_X1 U997 ( .A1(n1291), .A2(n1016), .ZN(n1290) );
XOR2_X1 U998 ( .A(KEYINPUT34), .B(n1292), .Z(n1291) );
NAND2_X1 U999 ( .A1(n1292), .A2(G107), .ZN(n1289) );
XOR2_X1 U1000 ( .A(n1293), .B(n1263), .Z(n1155) );
XOR2_X1 U1001 ( .A(G110), .B(n1294), .Z(n1263) );
XOR2_X1 U1002 ( .A(G140), .B(G128), .Z(n1294) );
XOR2_X1 U1003 ( .A(n1275), .B(n1295), .Z(n1293) );
AND2_X1 U1004 ( .A1(n1024), .A2(G227), .ZN(n1295) );
XOR2_X1 U1005 ( .A(n1097), .B(n1296), .Z(n1275) );
NOR2_X1 U1006 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U1007 ( .A(n1299), .B(KEYINPUT40), .Z(n1298) );
NAND2_X1 U1008 ( .A1(G134), .A2(n1096), .ZN(n1299) );
NOR2_X1 U1009 ( .A1(G134), .A2(n1096), .ZN(n1297) );
INV_X1 U1010 ( .A(G137), .ZN(n1096) );
XNOR2_X1 U1011 ( .A(G131), .B(n1300), .ZN(n1097) );
XOR2_X1 U1012 ( .A(KEYINPUT51), .B(KEYINPUT15), .Z(n1287) );
INV_X1 U1013 ( .A(n1204), .ZN(n1243) );
NAND2_X1 U1014 ( .A1(n1301), .A2(n1061), .ZN(n1204) );
NAND3_X1 U1015 ( .A1(n1302), .A2(n1024), .A3(G952), .ZN(n1061) );
OR2_X1 U1016 ( .A1(n1118), .A2(n1240), .ZN(n1301) );
NAND2_X1 U1017 ( .A1(G902), .A2(n1302), .ZN(n1240) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1019 ( .A(KEYINPUT12), .B(G237), .Z(n1303) );
OR2_X1 U1020 ( .A1(n1024), .A2(G898), .ZN(n1118) );
INV_X1 U1021 ( .A(n1253), .ZN(n1205) );
NOR2_X1 U1022 ( .A1(n1229), .A2(n1043), .ZN(n1253) );
XOR2_X1 U1023 ( .A(n1304), .B(n1305), .Z(n1043) );
NOR2_X1 U1024 ( .A1(n1306), .A2(n1166), .ZN(n1305) );
INV_X1 U1025 ( .A(G210), .ZN(n1166) );
XOR2_X1 U1026 ( .A(n1307), .B(KEYINPUT42), .Z(n1306) );
NAND2_X1 U1027 ( .A1(n1308), .A2(n1271), .ZN(n1304) );
INV_X1 U1028 ( .A(G902), .ZN(n1271) );
XOR2_X1 U1029 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U1030 ( .A(n1213), .B(n1165), .Z(n1310) );
XNOR2_X1 U1031 ( .A(n1120), .B(n1311), .ZN(n1165) );
NOR3_X1 U1032 ( .A1(n1124), .A2(KEYINPUT54), .A3(n1312), .ZN(n1311) );
INV_X1 U1033 ( .A(n1123), .ZN(n1312) );
NAND2_X1 U1034 ( .A1(n1313), .A2(n1126), .ZN(n1123) );
NOR2_X1 U1035 ( .A1(n1126), .A2(n1313), .ZN(n1124) );
XNOR2_X1 U1036 ( .A(G107), .B(n1292), .ZN(n1313) );
XOR2_X1 U1037 ( .A(G101), .B(G104), .Z(n1292) );
XOR2_X1 U1038 ( .A(G113), .B(n1314), .Z(n1126) );
NOR2_X1 U1039 ( .A1(n1282), .A2(n1315), .ZN(n1314) );
NOR2_X1 U1040 ( .A1(G119), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1041 ( .A(KEYINPUT24), .B(G116), .Z(n1316) );
NOR2_X1 U1042 ( .A1(n1244), .A2(G116), .ZN(n1282) );
INV_X1 U1043 ( .A(G119), .ZN(n1244) );
XNOR2_X1 U1044 ( .A(G110), .B(n1317), .ZN(n1120) );
NOR2_X1 U1045 ( .A1(G122), .A2(KEYINPUT25), .ZN(n1317) );
INV_X1 U1046 ( .A(n1210), .ZN(n1213) );
XOR2_X1 U1047 ( .A(n1318), .B(n1319), .Z(n1210) );
XOR2_X1 U1048 ( .A(KEYINPUT52), .B(G125), .Z(n1319) );
XOR2_X1 U1049 ( .A(n1276), .B(n1300), .Z(n1318) );
XOR2_X1 U1050 ( .A(G143), .B(G146), .Z(n1300) );
NAND2_X1 U1051 ( .A1(n1320), .A2(n1231), .ZN(n1276) );
INV_X1 U1052 ( .A(G128), .ZN(n1231) );
XNOR2_X1 U1053 ( .A(KEYINPUT5), .B(KEYINPUT2), .ZN(n1320) );
XOR2_X1 U1054 ( .A(n1212), .B(KEYINPUT60), .Z(n1309) );
NAND2_X1 U1055 ( .A1(G224), .A2(n1321), .ZN(n1212) );
XOR2_X1 U1056 ( .A(KEYINPUT30), .B(G953), .Z(n1321) );
XOR2_X1 U1057 ( .A(n1044), .B(KEYINPUT49), .Z(n1229) );
AND2_X1 U1058 ( .A1(G214), .A2(n1307), .ZN(n1044) );
OR2_X1 U1059 ( .A1(G902), .A2(G237), .ZN(n1307) );
NOR2_X1 U1060 ( .A1(n1322), .A2(n1217), .ZN(n1052) );
XNOR2_X1 U1061 ( .A(n1075), .B(KEYINPUT41), .ZN(n1217) );
XOR2_X1 U1062 ( .A(G475), .B(n1323), .Z(n1075) );
NOR2_X1 U1063 ( .A1(G902), .A2(n1140), .ZN(n1323) );
XNOR2_X1 U1064 ( .A(n1324), .B(n1325), .ZN(n1140) );
XOR2_X1 U1065 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1066 ( .A(G104), .B(n1328), .Z(n1327) );
NOR2_X1 U1067 ( .A1(KEYINPUT44), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1068 ( .A(n1216), .B(n1330), .Z(n1329) );
NAND2_X1 U1069 ( .A1(n1284), .A2(G214), .ZN(n1330) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1284) );
XOR2_X1 U1071 ( .A(G122), .B(G113), .Z(n1326) );
XOR2_X1 U1072 ( .A(n1331), .B(n1332), .Z(n1324) );
XOR2_X1 U1073 ( .A(G146), .B(G140), .Z(n1332) );
XOR2_X1 U1074 ( .A(G131), .B(n1103), .Z(n1331) );
INV_X1 U1075 ( .A(G125), .ZN(n1103) );
INV_X1 U1076 ( .A(n1220), .ZN(n1322) );
XOR2_X1 U1077 ( .A(n1076), .B(G478), .Z(n1220) );
OR2_X1 U1078 ( .A1(n1137), .A2(G902), .ZN(n1076) );
XNOR2_X1 U1079 ( .A(n1333), .B(n1334), .ZN(n1137) );
AND2_X1 U1080 ( .A1(n1266), .A2(G217), .ZN(n1334) );
AND2_X1 U1081 ( .A1(G234), .A2(n1024), .ZN(n1266) );
INV_X1 U1082 ( .A(G953), .ZN(n1024) );
NAND2_X1 U1083 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
NAND2_X1 U1084 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1085 ( .A(n1016), .B(n1339), .Z(n1338) );
INV_X1 U1086 ( .A(G107), .ZN(n1016) );
XOR2_X1 U1087 ( .A(n1216), .B(n1098), .Z(n1337) );
INV_X1 U1088 ( .A(G143), .ZN(n1216) );
XOR2_X1 U1089 ( .A(n1340), .B(KEYINPUT14), .Z(n1335) );
NAND2_X1 U1090 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1091 ( .A(G143), .B(n1098), .Z(n1342) );
XOR2_X1 U1092 ( .A(G128), .B(G134), .Z(n1098) );
XOR2_X1 U1093 ( .A(n1339), .B(G107), .Z(n1341) );
NAND2_X1 U1094 ( .A1(KEYINPUT45), .A2(n1343), .ZN(n1339) );
XNOR2_X1 U1095 ( .A(G122), .B(n1344), .ZN(n1343) );
NAND2_X1 U1096 ( .A1(KEYINPUT32), .A2(G116), .ZN(n1344) );
endmodule


