//Key = 0000001110100110011000101111010111000000000111011111111100000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337;

XNOR2_X1 U729 ( .A(n1017), .B(n1018), .ZN(G9) );
NAND2_X1 U730 ( .A1(KEYINPUT51), .A2(G107), .ZN(n1018) );
NAND4_X1 U731 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(G75) );
NAND4_X1 U732 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1021) );
NOR4_X1 U733 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U734 ( .A(n1031), .B(n1032), .Z(n1029) );
XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT43), .Z(n1032) );
XOR2_X1 U736 ( .A(n1033), .B(n1034), .Z(n1031) );
NOR2_X1 U737 ( .A1(KEYINPUT15), .A2(n1035), .ZN(n1034) );
XOR2_X1 U738 ( .A(n1036), .B(G472), .Z(n1028) );
NAND2_X1 U739 ( .A1(KEYINPUT63), .A2(n1037), .ZN(n1036) );
XNOR2_X1 U740 ( .A(n1038), .B(n1039), .ZN(n1025) );
NOR2_X1 U741 ( .A1(KEYINPUT42), .A2(n1040), .ZN(n1039) );
XOR2_X1 U742 ( .A(n1041), .B(n1042), .Z(n1023) );
XOR2_X1 U743 ( .A(KEYINPUT7), .B(KEYINPUT3), .Z(n1042) );
XNOR2_X1 U744 ( .A(G475), .B(n1043), .ZN(n1041) );
NOR2_X1 U745 ( .A1(n1044), .A2(KEYINPUT60), .ZN(n1043) );
NAND2_X1 U746 ( .A1(n1045), .A2(n1046), .ZN(n1020) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND4_X1 U748 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NAND2_X1 U749 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U750 ( .A1(n1024), .A2(n1055), .ZN(n1054) );
NAND2_X1 U751 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U752 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U753 ( .A1(n1060), .A2(n1061), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U755 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND4_X1 U756 ( .A1(n1024), .A2(n1060), .A3(n1066), .A4(n1067), .ZN(n1047) );
NAND2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U758 ( .A1(n1050), .A2(n1052), .ZN(n1069) );
NAND2_X1 U759 ( .A1(n1070), .A2(n1049), .ZN(n1066) );
NAND2_X1 U760 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
OR2_X1 U761 ( .A1(n1052), .A2(n1050), .ZN(n1072) );
OR3_X1 U762 ( .A1(n1073), .A2(n1074), .A3(n1027), .ZN(n1071) );
INV_X1 U763 ( .A(n1075), .ZN(n1045) );
XOR2_X1 U764 ( .A(n1076), .B(n1077), .Z(G72) );
NOR2_X1 U765 ( .A1(n1078), .A2(n1022), .ZN(n1077) );
AND2_X1 U766 ( .A1(G227), .A2(G900), .ZN(n1078) );
NOR3_X1 U767 ( .A1(KEYINPUT0), .A2(n1079), .A3(n1080), .ZN(n1076) );
NOR2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U769 ( .A(n1083), .B(KEYINPUT53), .Z(n1082) );
NAND2_X1 U770 ( .A1(n1022), .A2(n1084), .ZN(n1083) );
INV_X1 U771 ( .A(n1085), .ZN(n1081) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1085), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XOR2_X1 U774 ( .A(KEYINPUT46), .B(n1089), .Z(n1087) );
NOR2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U776 ( .A(n1092), .B(KEYINPUT6), .Z(n1091) );
NAND2_X1 U777 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U778 ( .A(KEYINPUT44), .B(n1095), .ZN(n1094) );
NOR2_X1 U779 ( .A1(n1095), .A2(n1093), .ZN(n1090) );
XNOR2_X1 U780 ( .A(n1096), .B(n1097), .ZN(n1093) );
XOR2_X1 U781 ( .A(n1098), .B(G140), .Z(n1095) );
NAND2_X1 U782 ( .A1(KEYINPUT18), .A2(n1099), .ZN(n1098) );
NAND2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(G69) );
NAND2_X1 U784 ( .A1(G953), .A2(n1102), .ZN(n1101) );
NAND2_X1 U785 ( .A1(G898), .A2(n1103), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U787 ( .A(n1106), .B(KEYINPUT30), .Z(n1100) );
NAND2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U789 ( .A1(G953), .A2(n1105), .ZN(n1108) );
INV_X1 U790 ( .A(G224), .ZN(n1105) );
XOR2_X1 U791 ( .A(n1104), .B(n1109), .Z(n1107) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(n1104) );
XNOR2_X1 U793 ( .A(KEYINPUT45), .B(n1112), .ZN(n1111) );
INV_X1 U794 ( .A(n1113), .ZN(n1112) );
XNOR2_X1 U795 ( .A(n1114), .B(n1115), .ZN(n1110) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XOR2_X1 U797 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND3_X1 U798 ( .A1(n1120), .A2(n1038), .A3(KEYINPUT27), .ZN(n1118) );
INV_X1 U799 ( .A(n1121), .ZN(n1038) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1122), .ZN(G63) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U802 ( .A1(n1120), .A2(G478), .ZN(n1123) );
NOR2_X1 U803 ( .A1(n1116), .A2(n1125), .ZN(G60) );
NOR3_X1 U804 ( .A1(n1044), .A2(n1126), .A3(n1127), .ZN(n1125) );
AND3_X1 U805 ( .A1(n1128), .A2(G475), .A3(n1120), .ZN(n1127) );
NOR2_X1 U806 ( .A1(n1129), .A2(n1128), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1019), .A2(n1130), .ZN(n1129) );
XOR2_X1 U808 ( .A(G104), .B(n1131), .Z(G6) );
NOR2_X1 U809 ( .A1(n1116), .A2(n1132), .ZN(G57) );
XOR2_X1 U810 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U811 ( .A(n1135), .B(n1136), .ZN(n1134) );
AND2_X1 U812 ( .A1(G472), .A2(n1120), .ZN(n1136) );
XNOR2_X1 U813 ( .A(n1137), .B(n1138), .ZN(n1133) );
NOR2_X1 U814 ( .A1(G101), .A2(KEYINPUT19), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1116), .A2(n1139), .ZN(G54) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U817 ( .A(n1113), .B(n1142), .ZN(n1141) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1140) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U820 ( .A1(KEYINPUT28), .A2(n1147), .ZN(n1146) );
AND2_X1 U821 ( .A1(G469), .A2(n1120), .ZN(n1145) );
NAND2_X1 U822 ( .A1(KEYINPUT25), .A2(n1097), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1116), .A2(n1148), .ZN(G51) );
XNOR2_X1 U824 ( .A(n1149), .B(n1150), .ZN(n1148) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
INV_X1 U827 ( .A(n1120), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1019), .ZN(n1120) );
AND2_X1 U829 ( .A1(n1109), .A2(n1086), .ZN(n1019) );
INV_X1 U830 ( .A(n1084), .ZN(n1086) );
NAND2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1084) );
NOR4_X1 U832 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1157) );
INV_X1 U833 ( .A(n1162), .ZN(n1159) );
INV_X1 U834 ( .A(n1163), .ZN(n1158) );
NOR4_X1 U835 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U837 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
INV_X1 U838 ( .A(KEYINPUT29), .ZN(n1171) );
NOR3_X1 U839 ( .A1(n1172), .A2(n1173), .A3(n1056), .ZN(n1165) );
NOR2_X1 U840 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U841 ( .A1(n1176), .A2(n1168), .ZN(n1175) );
NOR3_X1 U842 ( .A1(n1062), .A2(KEYINPUT29), .A3(n1177), .ZN(n1174) );
AND4_X1 U843 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1109) );
NOR4_X1 U844 ( .A1(n1182), .A2(n1017), .A3(n1131), .A4(n1183), .ZN(n1181) );
NOR3_X1 U845 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U847 ( .A(KEYINPUT57), .ZN(n1188) );
NOR4_X1 U848 ( .A1(n1189), .A2(n1027), .A3(n1190), .A4(n1068), .ZN(n1187) );
NOR2_X1 U849 ( .A1(KEYINPUT57), .A2(n1191), .ZN(n1185) );
AND3_X1 U850 ( .A1(n1192), .A2(n1060), .A3(n1073), .ZN(n1131) );
AND3_X1 U851 ( .A1(n1074), .A2(n1060), .A3(n1192), .ZN(n1017) );
AND2_X1 U852 ( .A1(n1193), .A2(n1194), .ZN(n1180) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1151) );
XOR2_X1 U854 ( .A(n1197), .B(KEYINPUT10), .Z(n1196) );
NOR2_X1 U855 ( .A1(n1022), .A2(G952), .ZN(n1116) );
XNOR2_X1 U856 ( .A(n1164), .B(n1198), .ZN(G48) );
NOR2_X1 U857 ( .A1(G146), .A2(KEYINPUT11), .ZN(n1198) );
AND2_X1 U858 ( .A1(n1199), .A2(n1073), .ZN(n1164) );
XNOR2_X1 U859 ( .A(G143), .B(n1170), .ZN(G45) );
NAND4_X1 U860 ( .A1(n1200), .A2(n1177), .A3(n1201), .A4(n1189), .ZN(n1170) );
XOR2_X1 U861 ( .A(G140), .B(n1161), .Z(G42) );
AND3_X1 U862 ( .A1(n1202), .A2(n1024), .A3(n1200), .ZN(n1161) );
XOR2_X1 U863 ( .A(G137), .B(n1160), .Z(G39) );
NOR3_X1 U864 ( .A1(n1184), .A2(n1168), .A3(n1172), .ZN(n1160) );
XNOR2_X1 U865 ( .A(G134), .B(n1203), .ZN(G36) );
NAND4_X1 U866 ( .A1(n1068), .A2(n1052), .A3(n1204), .A4(n1205), .ZN(n1203) );
NOR3_X1 U867 ( .A1(n1056), .A2(n1176), .A3(n1168), .ZN(n1205) );
INV_X1 U868 ( .A(n1074), .ZN(n1176) );
XNOR2_X1 U869 ( .A(KEYINPUT32), .B(n1206), .ZN(n1204) );
XNOR2_X1 U870 ( .A(G131), .B(n1207), .ZN(G33) );
NAND2_X1 U871 ( .A1(n1208), .A2(n1024), .ZN(n1207) );
INV_X1 U872 ( .A(n1168), .ZN(n1024) );
NAND2_X1 U873 ( .A1(n1065), .A2(n1209), .ZN(n1168) );
XOR2_X1 U874 ( .A(n1169), .B(KEYINPUT47), .Z(n1208) );
NAND3_X1 U875 ( .A1(n1073), .A2(n1201), .A3(n1200), .ZN(n1169) );
NAND2_X1 U876 ( .A1(n1210), .A2(n1211), .ZN(G30) );
NAND2_X1 U877 ( .A1(G128), .A2(n1162), .ZN(n1211) );
XOR2_X1 U878 ( .A(n1212), .B(KEYINPUT23), .Z(n1210) );
OR2_X1 U879 ( .A1(n1162), .A2(G128), .ZN(n1212) );
NAND2_X1 U880 ( .A1(n1199), .A2(n1074), .ZN(n1162) );
AND4_X1 U881 ( .A1(n1213), .A2(n1200), .A3(n1189), .A4(n1059), .ZN(n1199) );
INV_X1 U882 ( .A(n1172), .ZN(n1200) );
NAND3_X1 U883 ( .A1(n1052), .A2(n1206), .A3(n1068), .ZN(n1172) );
XNOR2_X1 U884 ( .A(n1214), .B(n1182), .ZN(G3) );
AND3_X1 U885 ( .A1(n1050), .A2(n1192), .A3(n1201), .ZN(n1182) );
XNOR2_X1 U886 ( .A(G125), .B(n1163), .ZN(G27) );
NAND3_X1 U887 ( .A1(n1215), .A2(n1206), .A3(n1202), .ZN(n1163) );
AND3_X1 U888 ( .A1(n1058), .A2(n1059), .A3(n1073), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1216), .A2(n1075), .ZN(n1206) );
NAND3_X1 U890 ( .A1(G902), .A2(n1217), .A3(n1218), .ZN(n1216) );
INV_X1 U891 ( .A(n1088), .ZN(n1218) );
NAND2_X1 U892 ( .A1(G953), .A2(n1219), .ZN(n1088) );
XOR2_X1 U893 ( .A(KEYINPUT50), .B(G900), .Z(n1219) );
XNOR2_X1 U894 ( .A(G122), .B(n1194), .ZN(G24) );
NAND3_X1 U895 ( .A1(n1191), .A2(n1060), .A3(n1177), .ZN(n1194) );
NOR2_X1 U896 ( .A1(n1220), .A2(n1221), .ZN(n1177) );
AND2_X1 U897 ( .A1(n1222), .A2(n1058), .ZN(n1060) );
XNOR2_X1 U898 ( .A(n1223), .B(n1224), .ZN(G21) );
NOR2_X1 U899 ( .A1(n1225), .A2(n1184), .ZN(n1224) );
NAND3_X1 U900 ( .A1(n1050), .A2(n1059), .A3(n1213), .ZN(n1184) );
XNOR2_X1 U901 ( .A(G116), .B(n1193), .ZN(G18) );
NAND3_X1 U902 ( .A1(n1191), .A2(n1074), .A3(n1201), .ZN(n1193) );
NOR2_X1 U903 ( .A1(n1226), .A2(n1221), .ZN(n1074) );
INV_X1 U904 ( .A(n1030), .ZN(n1221) );
XNOR2_X1 U905 ( .A(G113), .B(n1178), .ZN(G15) );
NAND3_X1 U906 ( .A1(n1201), .A2(n1191), .A3(n1073), .ZN(n1178) );
NOR2_X1 U907 ( .A1(n1030), .A2(n1220), .ZN(n1073) );
INV_X1 U908 ( .A(n1225), .ZN(n1191) );
NAND2_X1 U909 ( .A1(n1215), .A2(n1227), .ZN(n1225) );
NOR3_X1 U910 ( .A1(n1062), .A2(n1027), .A3(n1068), .ZN(n1215) );
INV_X1 U911 ( .A(n1056), .ZN(n1201) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1222), .ZN(n1056) );
INV_X1 U913 ( .A(n1059), .ZN(n1222) );
XOR2_X1 U914 ( .A(n1058), .B(KEYINPUT33), .Z(n1213) );
XNOR2_X1 U915 ( .A(G110), .B(n1179), .ZN(G12) );
NAND4_X1 U916 ( .A1(n1050), .A2(n1192), .A3(n1058), .A4(n1059), .ZN(n1179) );
XOR2_X1 U917 ( .A(n1228), .B(n1121), .Z(n1059) );
NAND2_X1 U918 ( .A1(G217), .A2(n1229), .ZN(n1121) );
XOR2_X1 U919 ( .A(n1040), .B(KEYINPUT35), .Z(n1228) );
NAND2_X1 U920 ( .A1(n1230), .A2(n1119), .ZN(n1040) );
XOR2_X1 U921 ( .A(n1231), .B(n1232), .Z(n1119) );
XNOR2_X1 U922 ( .A(n1233), .B(n1234), .ZN(n1232) );
NOR2_X1 U923 ( .A1(KEYINPUT21), .A2(n1235), .ZN(n1234) );
XOR2_X1 U924 ( .A(G110), .B(n1236), .Z(n1235) );
XNOR2_X1 U925 ( .A(G128), .B(n1223), .ZN(n1236) );
XOR2_X1 U926 ( .A(n1237), .B(n1238), .Z(n1231) );
NAND2_X1 U927 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
XNOR2_X1 U928 ( .A(G137), .B(n1241), .ZN(n1240) );
NAND2_X1 U929 ( .A1(n1242), .A2(G221), .ZN(n1241) );
XOR2_X1 U930 ( .A(KEYINPUT62), .B(KEYINPUT13), .Z(n1239) );
XNOR2_X1 U931 ( .A(G902), .B(KEYINPUT39), .ZN(n1230) );
XOR2_X1 U932 ( .A(n1037), .B(G472), .Z(n1058) );
NAND3_X1 U933 ( .A1(n1243), .A2(n1155), .A3(n1244), .ZN(n1037) );
NAND2_X1 U934 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U935 ( .A1(KEYINPUT26), .A2(n1247), .ZN(n1246) );
NAND2_X1 U936 ( .A1(KEYINPUT31), .A2(n1248), .ZN(n1247) );
INV_X1 U937 ( .A(n1137), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1249), .A2(n1250), .ZN(n1243) );
NAND2_X1 U939 ( .A1(KEYINPUT31), .A2(n1251), .ZN(n1250) );
NAND2_X1 U940 ( .A1(KEYINPUT26), .A2(n1137), .ZN(n1251) );
XNOR2_X1 U941 ( .A(n1252), .B(n1253), .ZN(n1137) );
XNOR2_X1 U942 ( .A(n1254), .B(n1255), .ZN(n1253) );
NOR2_X1 U943 ( .A1(KEYINPUT41), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U944 ( .A(G116), .B(G119), .ZN(n1256) );
XNOR2_X1 U945 ( .A(n1257), .B(n1258), .ZN(n1252) );
INV_X1 U946 ( .A(n1096), .ZN(n1258) );
INV_X1 U947 ( .A(n1248), .ZN(n1249) );
XOR2_X1 U948 ( .A(n1135), .B(n1214), .Z(n1248) );
INV_X1 U949 ( .A(G101), .ZN(n1214) );
NAND3_X1 U950 ( .A1(n1259), .A2(n1022), .A3(G210), .ZN(n1135) );
NOR4_X1 U951 ( .A1(n1062), .A2(n1049), .A3(n1190), .A4(n1027), .ZN(n1192) );
INV_X1 U952 ( .A(n1052), .ZN(n1027) );
NAND2_X1 U953 ( .A1(G221), .A2(n1229), .ZN(n1052) );
NAND2_X1 U954 ( .A1(n1260), .A2(n1155), .ZN(n1229) );
XNOR2_X1 U955 ( .A(G234), .B(KEYINPUT48), .ZN(n1260) );
INV_X1 U956 ( .A(n1227), .ZN(n1190) );
NAND2_X1 U957 ( .A1(n1075), .A2(n1261), .ZN(n1227) );
NAND4_X1 U958 ( .A1(G902), .A2(G953), .A3(n1217), .A4(n1262), .ZN(n1261) );
INV_X1 U959 ( .A(G898), .ZN(n1262) );
NAND3_X1 U960 ( .A1(n1217), .A2(n1022), .A3(G952), .ZN(n1075) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1217) );
INV_X1 U962 ( .A(n1068), .ZN(n1049) );
XNOR2_X1 U963 ( .A(n1033), .B(n1035), .ZN(n1068) );
XOR2_X1 U964 ( .A(G469), .B(KEYINPUT37), .Z(n1035) );
NAND2_X1 U965 ( .A1(n1263), .A2(n1155), .ZN(n1033) );
XOR2_X1 U966 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U967 ( .A(n1147), .B(n1142), .Z(n1265) );
XNOR2_X1 U968 ( .A(n1096), .B(n1266), .ZN(n1142) );
AND2_X1 U969 ( .A1(n1022), .A2(G227), .ZN(n1266) );
XOR2_X1 U970 ( .A(G131), .B(n1267), .Z(n1096) );
XOR2_X1 U971 ( .A(G137), .B(G134), .Z(n1267) );
XNOR2_X1 U972 ( .A(G110), .B(G140), .ZN(n1147) );
XNOR2_X1 U973 ( .A(KEYINPUT40), .B(n1268), .ZN(n1264) );
NOR2_X1 U974 ( .A1(KEYINPUT1), .A2(n1269), .ZN(n1268) );
NOR2_X1 U975 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U976 ( .A(KEYINPUT59), .B(n1272), .Z(n1271) );
NOR2_X1 U977 ( .A1(n1113), .A2(n1097), .ZN(n1272) );
AND2_X1 U978 ( .A1(n1113), .A2(n1097), .ZN(n1270) );
XOR2_X1 U979 ( .A(n1273), .B(n1274), .Z(n1097) );
NAND3_X1 U980 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1273) );
NAND2_X1 U981 ( .A1(n1278), .A2(G146), .ZN(n1277) );
NAND2_X1 U982 ( .A1(n1279), .A2(n1280), .ZN(n1276) );
INV_X1 U983 ( .A(KEYINPUT55), .ZN(n1280) );
NAND2_X1 U984 ( .A1(n1281), .A2(n1233), .ZN(n1279) );
XNOR2_X1 U985 ( .A(KEYINPUT22), .B(n1282), .ZN(n1281) );
NAND2_X1 U986 ( .A1(KEYINPUT55), .A2(n1283), .ZN(n1275) );
NAND2_X1 U987 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
OR2_X1 U988 ( .A1(n1282), .A2(KEYINPUT22), .ZN(n1285) );
NAND3_X1 U989 ( .A1(n1282), .A2(n1233), .A3(KEYINPUT22), .ZN(n1284) );
INV_X1 U990 ( .A(n1189), .ZN(n1062) );
NOR2_X1 U991 ( .A1(n1065), .A2(n1064), .ZN(n1189) );
INV_X1 U992 ( .A(n1209), .ZN(n1064) );
NAND2_X1 U993 ( .A1(G214), .A2(n1286), .ZN(n1209) );
XNOR2_X1 U994 ( .A(n1287), .B(n1153), .ZN(n1065) );
NAND2_X1 U995 ( .A1(G210), .A2(n1286), .ZN(n1153) );
NAND2_X1 U996 ( .A1(n1259), .A2(n1155), .ZN(n1286) );
NAND2_X1 U997 ( .A1(n1288), .A2(n1155), .ZN(n1287) );
XOR2_X1 U998 ( .A(n1289), .B(KEYINPUT14), .Z(n1288) );
NAND3_X1 U999 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
NAND3_X1 U1000 ( .A1(n1293), .A2(n1197), .A3(n1294), .ZN(n1292) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U1002 ( .A1(n1297), .A2(n1149), .ZN(n1296) );
NAND3_X1 U1003 ( .A1(n1298), .A2(n1299), .A3(n1295), .ZN(n1291) );
INV_X1 U1004 ( .A(KEYINPUT34), .ZN(n1295) );
NAND3_X1 U1005 ( .A1(n1293), .A2(n1197), .A3(n1297), .ZN(n1299) );
XOR2_X1 U1006 ( .A(KEYINPUT24), .B(KEYINPUT16), .Z(n1297) );
NAND2_X1 U1007 ( .A1(n1300), .A2(n1301), .ZN(n1197) );
INV_X1 U1008 ( .A(n1195), .ZN(n1293) );
NOR2_X1 U1009 ( .A1(n1301), .A2(n1300), .ZN(n1195) );
XOR2_X1 U1010 ( .A(n1257), .B(G125), .Z(n1300) );
XNOR2_X1 U1011 ( .A(n1302), .B(n1278), .ZN(n1257) );
INV_X1 U1012 ( .A(n1282), .ZN(n1278) );
XOR2_X1 U1013 ( .A(n1303), .B(KEYINPUT36), .Z(n1282) );
XNOR2_X1 U1014 ( .A(G146), .B(n1304), .ZN(n1302) );
NOR2_X1 U1015 ( .A1(KEYINPUT4), .A2(n1274), .ZN(n1304) );
XNOR2_X1 U1016 ( .A(G128), .B(KEYINPUT49), .ZN(n1274) );
NAND2_X1 U1017 ( .A1(G224), .A2(n1305), .ZN(n1301) );
XNOR2_X1 U1018 ( .A(KEYINPUT61), .B(n1022), .ZN(n1305) );
INV_X1 U1019 ( .A(n1149), .ZN(n1298) );
NAND2_X1 U1020 ( .A1(KEYINPUT34), .A2(n1149), .ZN(n1290) );
XNOR2_X1 U1021 ( .A(n1306), .B(n1115), .ZN(n1149) );
XOR2_X1 U1022 ( .A(G110), .B(G122), .Z(n1115) );
NAND3_X1 U1023 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
OR2_X1 U1024 ( .A1(n1310), .A2(KEYINPUT17), .ZN(n1309) );
INV_X1 U1025 ( .A(n1114), .ZN(n1310) );
NAND3_X1 U1026 ( .A1(KEYINPUT17), .A2(n1311), .A3(n1113), .ZN(n1308) );
OR2_X1 U1027 ( .A1(n1113), .A2(n1311), .ZN(n1307) );
NOR2_X1 U1028 ( .A1(KEYINPUT2), .A2(n1114), .ZN(n1311) );
XNOR2_X1 U1029 ( .A(n1312), .B(n1313), .ZN(n1114) );
XNOR2_X1 U1030 ( .A(n1254), .B(n1314), .ZN(n1313) );
NOR2_X1 U1031 ( .A1(KEYINPUT9), .A2(n1223), .ZN(n1314) );
INV_X1 U1032 ( .A(G119), .ZN(n1223) );
INV_X1 U1033 ( .A(G113), .ZN(n1254) );
XNOR2_X1 U1034 ( .A(G116), .B(KEYINPUT38), .ZN(n1312) );
XOR2_X1 U1035 ( .A(G101), .B(n1315), .Z(n1113) );
XOR2_X1 U1036 ( .A(G107), .B(G104), .Z(n1315) );
NOR2_X1 U1037 ( .A1(n1030), .A2(n1226), .ZN(n1050) );
INV_X1 U1038 ( .A(n1220), .ZN(n1226) );
XOR2_X1 U1039 ( .A(n1044), .B(n1130), .Z(n1220) );
INV_X1 U1040 ( .A(G475), .ZN(n1130) );
NOR2_X1 U1041 ( .A1(n1128), .A2(G902), .ZN(n1044) );
XOR2_X1 U1042 ( .A(n1316), .B(n1317), .Z(n1128) );
XOR2_X1 U1043 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1044 ( .A(n1320), .B(n1321), .ZN(n1319) );
NOR2_X1 U1045 ( .A1(KEYINPUT58), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1046 ( .A(n1323), .B(n1324), .ZN(n1322) );
AND3_X1 U1047 ( .A1(G214), .A2(n1022), .A3(n1259), .ZN(n1323) );
INV_X1 U1048 ( .A(G237), .ZN(n1259) );
NAND2_X1 U1049 ( .A1(KEYINPUT52), .A2(G122), .ZN(n1320) );
NOR2_X1 U1050 ( .A1(KEYINPUT20), .A2(n1238), .ZN(n1318) );
XNOR2_X1 U1051 ( .A(n1099), .B(G140), .ZN(n1238) );
INV_X1 U1052 ( .A(G125), .ZN(n1099) );
XOR2_X1 U1053 ( .A(n1325), .B(n1326), .Z(n1316) );
XNOR2_X1 U1054 ( .A(n1233), .B(G131), .ZN(n1326) );
INV_X1 U1055 ( .A(G146), .ZN(n1233) );
XNOR2_X1 U1056 ( .A(G104), .B(G113), .ZN(n1325) );
XOR2_X1 U1057 ( .A(G478), .B(n1327), .Z(n1030) );
AND2_X1 U1058 ( .A1(n1155), .A2(n1124), .ZN(n1327) );
XNOR2_X1 U1059 ( .A(n1328), .B(n1329), .ZN(n1124) );
NOR2_X1 U1060 ( .A1(KEYINPUT5), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1061 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1062 ( .A(n1333), .B(n1334), .Z(n1332) );
NOR2_X1 U1063 ( .A1(KEYINPUT56), .A2(n1324), .ZN(n1334) );
INV_X1 U1064 ( .A(n1303), .ZN(n1324) );
XOR2_X1 U1065 ( .A(G143), .B(KEYINPUT12), .Z(n1303) );
XOR2_X1 U1066 ( .A(n1335), .B(G107), .Z(n1333) );
NAND2_X1 U1067 ( .A1(KEYINPUT8), .A2(n1336), .ZN(n1335) );
INV_X1 U1068 ( .A(G116), .ZN(n1336) );
XNOR2_X1 U1069 ( .A(G122), .B(n1337), .ZN(n1331) );
XOR2_X1 U1070 ( .A(G134), .B(G128), .Z(n1337) );
NAND2_X1 U1071 ( .A1(G217), .A2(n1242), .ZN(n1328) );
AND2_X1 U1072 ( .A1(G234), .A2(n1022), .ZN(n1242) );
INV_X1 U1073 ( .A(G953), .ZN(n1022) );
INV_X1 U1074 ( .A(G902), .ZN(n1155) );
endmodule


