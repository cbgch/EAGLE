//Key = 1111111100101000110111010100010010100001000010101100101110110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363;

XOR2_X1 U754 ( .A(n1043), .B(n1044), .Z(G9) );
XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT48), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR3_X1 U757 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND3_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND2_X1 U759 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U760 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND4_X1 U761 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U764 ( .A1(n1059), .A2(n1065), .A3(n1058), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1057), .A2(n1070), .ZN(n1063) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1058), .A2(n1073), .ZN(n1072) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U772 ( .A1(n1059), .A2(n1078), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U775 ( .A(n1083), .ZN(n1053) );
AND3_X1 U776 ( .A1(n1050), .A2(n1051), .A3(n1084), .ZN(n1045) );
NAND4_X1 U777 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1050) );
NOR4_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
XOR2_X1 U779 ( .A(G478), .B(n1093), .Z(n1092) );
XNOR2_X1 U780 ( .A(n1077), .B(KEYINPUT25), .ZN(n1090) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1089) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U783 ( .A1(n1098), .A2(KEYINPUT51), .ZN(n1096) );
XNOR2_X1 U784 ( .A(KEYINPUT57), .B(KEYINPUT19), .ZN(n1094) );
NOR3_X1 U785 ( .A1(n1068), .A2(n1099), .A3(n1100), .ZN(n1087) );
NAND2_X1 U786 ( .A1(n1101), .A2(G475), .ZN(n1086) );
XOR2_X1 U787 ( .A(n1102), .B(KEYINPUT11), .Z(n1101) );
NAND2_X1 U788 ( .A1(G469), .A2(n1103), .ZN(n1085) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1105), .ZN(G72) );
NAND3_X1 U790 ( .A1(n1106), .A2(n1107), .A3(G953), .ZN(n1105) );
XOR2_X1 U791 ( .A(n1108), .B(KEYINPUT16), .Z(n1104) );
NAND2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1051), .ZN(n1110) );
NAND2_X1 U794 ( .A1(n1107), .A2(n1112), .ZN(n1111) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1048), .ZN(n1112) );
OR2_X1 U796 ( .A1(n1107), .A2(n1106), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1114), .A2(G227), .ZN(n1106) );
XOR2_X1 U798 ( .A(n1115), .B(KEYINPUT23), .Z(n1114) );
OR3_X1 U799 ( .A1(n1048), .A2(n1116), .A3(n1113), .ZN(n1107) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U802 ( .A(KEYINPUT55), .B(n1121), .Z(n1117) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1119), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1122), .B(n1123), .Z(n1119) );
XOR2_X1 U805 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U806 ( .A(n1126), .B(KEYINPUT36), .Z(n1122) );
NOR2_X1 U807 ( .A1(n1051), .A2(G900), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(G69) );
NAND2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U810 ( .A1(G953), .A2(n1131), .A3(KEYINPUT12), .ZN(n1130) );
INV_X1 U811 ( .A(n1132), .ZN(n1129) );
NAND3_X1 U812 ( .A1(KEYINPUT12), .A2(n1133), .A3(n1132), .ZN(n1127) );
XOR2_X1 U813 ( .A(n1134), .B(n1135), .Z(n1132) );
AND2_X1 U814 ( .A1(n1049), .A2(n1051), .ZN(n1135) );
NAND3_X1 U815 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1134) );
NAND2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
XNOR2_X1 U817 ( .A(n1141), .B(KEYINPUT58), .ZN(n1139) );
NAND2_X1 U818 ( .A1(n1137), .A2(n1142), .ZN(n1133) );
NAND2_X1 U819 ( .A1(G953), .A2(n1131), .ZN(n1142) );
INV_X1 U820 ( .A(G224), .ZN(n1131) );
INV_X1 U821 ( .A(n1143), .ZN(n1137) );
NOR3_X1 U822 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(G66) );
NOR3_X1 U823 ( .A1(n1147), .A2(n1051), .A3(n1084), .ZN(n1146) );
INV_X1 U824 ( .A(G952), .ZN(n1084) );
AND2_X1 U825 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
INV_X1 U826 ( .A(KEYINPUT41), .ZN(n1147) );
XNOR2_X1 U827 ( .A(n1149), .B(n1150), .ZN(n1144) );
NOR3_X1 U828 ( .A1(n1151), .A2(KEYINPUT40), .A3(n1152), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1148), .A2(n1153), .ZN(G63) );
NOR3_X1 U830 ( .A1(n1093), .A2(n1154), .A3(n1155), .ZN(n1153) );
AND3_X1 U831 ( .A1(n1156), .A2(G478), .A3(n1157), .ZN(n1155) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1156), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1048), .A2(n1049), .ZN(n1159) );
NOR2_X1 U835 ( .A1(n1148), .A2(n1161), .ZN(G60) );
XOR2_X1 U836 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U837 ( .A1(KEYINPUT47), .A2(n1164), .ZN(n1163) );
NAND2_X1 U838 ( .A1(n1157), .A2(G475), .ZN(n1162) );
XOR2_X1 U839 ( .A(G104), .B(n1165), .Z(G6) );
NOR2_X1 U840 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U841 ( .A(KEYINPUT32), .B(n1168), .Z(n1167) );
NOR2_X1 U842 ( .A1(n1148), .A2(n1169), .ZN(G57) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1171) );
AND2_X1 U845 ( .A1(G472), .A2(n1157), .ZN(n1173) );
NOR3_X1 U846 ( .A1(n1174), .A2(n1148), .A3(n1175), .ZN(G54) );
NOR4_X1 U847 ( .A1(n1176), .A2(n1177), .A3(KEYINPUT43), .A4(n1178), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1181), .A2(n1182), .ZN(n1176) );
NOR2_X1 U850 ( .A1(n1051), .A2(G952), .ZN(n1148) );
NOR3_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1174) );
NOR2_X1 U852 ( .A1(n1182), .A2(n1180), .ZN(n1185) );
XNOR2_X1 U853 ( .A(n1181), .B(KEYINPUT14), .ZN(n1180) );
INV_X1 U854 ( .A(n1179), .ZN(n1182) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1179), .ZN(n1184) );
NAND2_X1 U856 ( .A1(n1186), .A2(n1187), .ZN(n1179) );
NAND2_X1 U857 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
AND2_X1 U858 ( .A1(n1157), .A2(G469), .ZN(n1181) );
INV_X1 U859 ( .A(n1151), .ZN(n1157) );
NOR2_X1 U860 ( .A1(KEYINPUT43), .A2(n1178), .ZN(n1183) );
XOR2_X1 U861 ( .A(n1190), .B(KEYINPUT7), .Z(n1178) );
NOR2_X1 U862 ( .A1(n1191), .A2(n1192), .ZN(G51) );
XOR2_X1 U863 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U864 ( .A1(n1195), .A2(n1151), .ZN(n1194) );
NAND2_X1 U865 ( .A1(G902), .A2(n1196), .ZN(n1151) );
OR2_X1 U866 ( .A1(n1049), .A2(n1048), .ZN(n1196) );
NAND4_X1 U867 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1048) );
NOR4_X1 U868 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR4_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1074), .A4(n1066), .ZN(n1204) );
NOR2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
AND3_X1 U871 ( .A1(KEYINPUT60), .A2(n1091), .A3(n1168), .ZN(n1207) );
INV_X1 U872 ( .A(n1209), .ZN(n1202) );
OR2_X1 U873 ( .A1(n1210), .A2(n1079), .ZN(n1199) );
OR3_X1 U874 ( .A1(n1211), .A2(KEYINPUT60), .A3(n1212), .ZN(n1198) );
NAND2_X1 U875 ( .A1(n1213), .A2(n1060), .ZN(n1197) );
NAND2_X1 U876 ( .A1(n1214), .A2(n1215), .ZN(n1060) );
NAND4_X1 U877 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1049) );
AND4_X1 U878 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
NOR2_X1 U879 ( .A1(n1044), .A2(n1224), .ZN(n1218) );
NOR2_X1 U880 ( .A1(n1166), .A2(n1215), .ZN(n1044) );
NAND2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1217) );
XOR2_X1 U882 ( .A(KEYINPUT30), .B(n1227), .Z(n1226) );
OR2_X1 U883 ( .A1(n1214), .A2(n1166), .ZN(n1216) );
NAND2_X1 U884 ( .A1(n1059), .A2(n1228), .ZN(n1166) );
XNOR2_X1 U885 ( .A(n1229), .B(n1230), .ZN(n1193) );
NAND2_X1 U886 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U887 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
NOR2_X1 U888 ( .A1(G952), .A2(n1235), .ZN(n1191) );
XOR2_X1 U889 ( .A(KEYINPUT49), .B(G953), .Z(n1235) );
XOR2_X1 U890 ( .A(n1236), .B(n1237), .Z(G48) );
NAND2_X1 U891 ( .A1(n1238), .A2(n1213), .ZN(n1237) );
XOR2_X1 U892 ( .A(n1214), .B(KEYINPUT39), .Z(n1238) );
INV_X1 U893 ( .A(n1168), .ZN(n1214) );
XOR2_X1 U894 ( .A(n1239), .B(n1240), .Z(G45) );
NOR2_X1 U895 ( .A1(KEYINPUT35), .A2(n1241), .ZN(n1240) );
NOR4_X1 U896 ( .A1(n1205), .A2(n1074), .A3(n1242), .A4(n1243), .ZN(n1239) );
XOR2_X1 U897 ( .A(n1066), .B(KEYINPUT9), .Z(n1242) );
INV_X1 U898 ( .A(n1244), .ZN(n1205) );
XOR2_X1 U899 ( .A(G140), .B(n1203), .Z(G42) );
AND2_X1 U900 ( .A1(n1245), .A2(n1246), .ZN(n1203) );
XOR2_X1 U901 ( .A(n1247), .B(n1209), .Z(G39) );
NAND4_X1 U902 ( .A1(n1248), .A2(n1246), .A3(n1061), .A4(n1077), .ZN(n1209) );
INV_X1 U903 ( .A(n1212), .ZN(n1246) );
XOR2_X1 U904 ( .A(G134), .B(n1201), .Z(G36) );
NOR3_X1 U905 ( .A1(n1215), .A2(n1074), .A3(n1212), .ZN(n1201) );
XOR2_X1 U906 ( .A(G131), .B(n1249), .Z(G33) );
NOR2_X1 U907 ( .A1(n1211), .A2(n1212), .ZN(n1249) );
NAND3_X1 U908 ( .A1(n1250), .A2(n1244), .A3(n1058), .ZN(n1212) );
INV_X1 U909 ( .A(n1091), .ZN(n1058) );
NAND2_X1 U910 ( .A1(n1082), .A2(n1251), .ZN(n1091) );
XNOR2_X1 U911 ( .A(G128), .B(n1252), .ZN(G30) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1253), .ZN(n1252) );
INV_X1 U913 ( .A(n1215), .ZN(n1253) );
AND4_X1 U914 ( .A1(n1077), .A2(n1244), .A3(n1225), .A4(n1254), .ZN(n1213) );
NOR2_X1 U915 ( .A1(n1066), .A2(n1076), .ZN(n1254) );
INV_X1 U916 ( .A(n1250), .ZN(n1066) );
XNOR2_X1 U917 ( .A(G101), .B(n1223), .ZN(G3) );
NAND3_X1 U918 ( .A1(n1228), .A2(n1255), .A3(n1061), .ZN(n1223) );
XOR2_X1 U919 ( .A(n1256), .B(n1257), .Z(G27) );
NAND2_X1 U920 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1257) );
NAND2_X1 U921 ( .A1(n1258), .A2(n1225), .ZN(n1256) );
XOR2_X1 U922 ( .A(n1210), .B(KEYINPUT56), .Z(n1258) );
NAND3_X1 U923 ( .A1(n1057), .A2(n1244), .A3(n1245), .ZN(n1210) );
AND3_X1 U924 ( .A1(n1076), .A2(n1077), .A3(n1168), .ZN(n1245) );
NAND2_X1 U925 ( .A1(n1083), .A2(n1259), .ZN(n1244) );
NAND3_X1 U926 ( .A1(G953), .A2(n1115), .A3(n1260), .ZN(n1259) );
INV_X1 U927 ( .A(G900), .ZN(n1115) );
XOR2_X1 U928 ( .A(n1261), .B(n1222), .Z(G24) );
NAND3_X1 U929 ( .A1(n1262), .A2(n1059), .A3(n1208), .ZN(n1222) );
INV_X1 U930 ( .A(n1243), .ZN(n1208) );
NAND3_X1 U931 ( .A1(n1263), .A2(n1225), .A3(n1264), .ZN(n1243) );
XOR2_X1 U932 ( .A(n1265), .B(KEYINPUT27), .Z(n1264) );
INV_X1 U933 ( .A(n1266), .ZN(n1262) );
XOR2_X1 U934 ( .A(n1267), .B(n1221), .Z(G21) );
NAND4_X1 U935 ( .A1(n1225), .A2(n1077), .A3(n1061), .A4(n1268), .ZN(n1221) );
NOR2_X1 U936 ( .A1(n1266), .A2(n1076), .ZN(n1268) );
XNOR2_X1 U937 ( .A(G116), .B(n1269), .ZN(G18) );
NAND2_X1 U938 ( .A1(n1227), .A2(n1225), .ZN(n1269) );
NOR3_X1 U939 ( .A1(n1215), .A2(n1074), .A3(n1266), .ZN(n1227) );
INV_X1 U940 ( .A(n1255), .ZN(n1074) );
NAND2_X1 U941 ( .A1(n1270), .A2(n1263), .ZN(n1215) );
XOR2_X1 U942 ( .A(G113), .B(n1224), .Z(G15) );
NOR3_X1 U943 ( .A1(n1266), .A2(n1079), .A3(n1211), .ZN(n1224) );
NAND2_X1 U944 ( .A1(n1168), .A2(n1255), .ZN(n1211) );
NAND2_X1 U945 ( .A1(n1271), .A2(n1272), .ZN(n1255) );
OR3_X1 U946 ( .A1(n1077), .A2(n1076), .A3(KEYINPUT45), .ZN(n1272) );
NAND2_X1 U947 ( .A1(KEYINPUT45), .A2(n1059), .ZN(n1271) );
NOR2_X1 U948 ( .A1(n1077), .A2(n1248), .ZN(n1059) );
NOR2_X1 U949 ( .A1(n1263), .A2(n1270), .ZN(n1168) );
INV_X1 U950 ( .A(n1225), .ZN(n1079) );
NAND2_X1 U951 ( .A1(n1057), .A2(n1273), .ZN(n1266) );
AND2_X1 U952 ( .A1(n1069), .A2(n1274), .ZN(n1057) );
XNOR2_X1 U953 ( .A(G110), .B(n1220), .ZN(G12) );
NAND4_X1 U954 ( .A1(n1061), .A2(n1228), .A3(n1076), .A4(n1077), .ZN(n1220) );
XOR2_X1 U955 ( .A(n1275), .B(n1152), .Z(n1077) );
NAND2_X1 U956 ( .A1(G217), .A2(n1276), .ZN(n1152) );
NAND2_X1 U957 ( .A1(n1149), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U958 ( .A(n1278), .B(n1279), .ZN(n1149) );
XOR2_X1 U959 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U960 ( .A(n1282), .B(n1283), .Z(n1281) );
NOR2_X1 U961 ( .A1(KEYINPUT31), .A2(n1284), .ZN(n1283) );
XOR2_X1 U962 ( .A(n1267), .B(G128), .Z(n1284) );
NAND3_X1 U963 ( .A1(G234), .A2(n1285), .A3(G221), .ZN(n1282) );
XOR2_X1 U964 ( .A(KEYINPUT2), .B(G953), .Z(n1285) );
NAND2_X1 U965 ( .A1(KEYINPUT10), .A2(n1247), .ZN(n1280) );
INV_X1 U966 ( .A(G137), .ZN(n1247) );
XNOR2_X1 U967 ( .A(n1188), .B(n1286), .ZN(n1278) );
XNOR2_X1 U968 ( .A(n1287), .B(n1288), .ZN(n1286) );
NOR2_X1 U969 ( .A1(KEYINPUT26), .A2(n1236), .ZN(n1288) );
INV_X1 U970 ( .A(G146), .ZN(n1236) );
NAND2_X1 U971 ( .A1(KEYINPUT52), .A2(n1289), .ZN(n1287) );
XOR2_X1 U972 ( .A(KEYINPUT29), .B(G125), .Z(n1289) );
INV_X1 U973 ( .A(n1248), .ZN(n1076) );
XNOR2_X1 U974 ( .A(n1098), .B(n1097), .ZN(n1248) );
XOR2_X1 U975 ( .A(G472), .B(KEYINPUT1), .Z(n1097) );
AND2_X1 U976 ( .A1(n1290), .A2(n1277), .ZN(n1098) );
XOR2_X1 U977 ( .A(n1170), .B(n1291), .Z(n1290) );
NOR2_X1 U978 ( .A1(KEYINPUT15), .A2(n1172), .ZN(n1291) );
NAND3_X1 U979 ( .A1(n1292), .A2(n1051), .A3(G210), .ZN(n1172) );
XOR2_X1 U980 ( .A(n1293), .B(n1294), .Z(n1170) );
XOR2_X1 U981 ( .A(G101), .B(n1295), .Z(n1294) );
XOR2_X1 U982 ( .A(n1296), .B(n1297), .Z(n1293) );
NOR3_X1 U983 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
NOR2_X1 U984 ( .A1(KEYINPUT46), .A2(n1301), .ZN(n1300) );
NOR3_X1 U985 ( .A1(n1302), .A2(G113), .A3(n1303), .ZN(n1299) );
INV_X1 U986 ( .A(KEYINPUT46), .ZN(n1302) );
AND2_X1 U987 ( .A1(n1303), .A2(G113), .ZN(n1298) );
NAND2_X1 U988 ( .A1(KEYINPUT44), .A2(n1301), .ZN(n1303) );
XOR2_X1 U989 ( .A(G116), .B(G119), .Z(n1301) );
AND3_X1 U990 ( .A1(n1225), .A2(n1273), .A3(n1250), .ZN(n1228) );
NOR2_X1 U991 ( .A1(n1068), .A2(n1069), .ZN(n1250) );
NOR2_X1 U992 ( .A1(n1304), .A2(n1100), .ZN(n1069) );
NOR2_X1 U993 ( .A1(n1103), .A2(G469), .ZN(n1100) );
AND2_X1 U994 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U995 ( .A(n1103), .B(KEYINPUT42), .Z(n1306) );
NAND2_X1 U996 ( .A1(n1307), .A2(n1277), .ZN(n1103) );
XOR2_X1 U997 ( .A(n1308), .B(n1309), .Z(n1307) );
INV_X1 U998 ( .A(n1190), .ZN(n1309) );
XOR2_X1 U999 ( .A(n1310), .B(n1311), .Z(n1190) );
XOR2_X1 U1000 ( .A(n1124), .B(n1296), .Z(n1311) );
XOR2_X1 U1001 ( .A(n1312), .B(n1313), .Z(n1296) );
INV_X1 U1002 ( .A(n1125), .ZN(n1313) );
XNOR2_X1 U1003 ( .A(G128), .B(n1314), .ZN(n1125) );
XOR2_X1 U1004 ( .A(G137), .B(G134), .Z(n1314) );
NAND2_X1 U1005 ( .A1(KEYINPUT34), .A2(n1126), .ZN(n1312) );
INV_X1 U1006 ( .A(G131), .ZN(n1126) );
XNOR2_X1 U1007 ( .A(KEYINPUT53), .B(n1315), .ZN(n1124) );
NOR2_X1 U1008 ( .A1(KEYINPUT38), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1009 ( .A(KEYINPUT50), .B(n1317), .Z(n1316) );
XOR2_X1 U1010 ( .A(n1318), .B(n1319), .Z(n1310) );
NAND2_X1 U1011 ( .A1(KEYINPUT6), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1012 ( .A(KEYINPUT22), .B(G101), .Z(n1320) );
NAND3_X1 U1013 ( .A1(n1321), .A2(n1322), .A3(n1186), .ZN(n1308) );
OR2_X1 U1014 ( .A1(n1189), .A2(n1188), .ZN(n1186) );
NAND3_X1 U1015 ( .A1(KEYINPUT0), .A2(n1188), .A3(n1189), .ZN(n1322) );
XOR2_X1 U1016 ( .A(G110), .B(G140), .Z(n1188) );
OR2_X1 U1017 ( .A1(n1189), .A2(KEYINPUT0), .ZN(n1321) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1051), .ZN(n1189) );
XNOR2_X1 U1019 ( .A(G469), .B(KEYINPUT3), .ZN(n1305) );
INV_X1 U1020 ( .A(n1274), .ZN(n1068) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1276), .ZN(n1274) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1277), .ZN(n1276) );
NAND2_X1 U1023 ( .A1(n1323), .A2(n1083), .ZN(n1273) );
NAND3_X1 U1024 ( .A1(n1324), .A2(n1051), .A3(G952), .ZN(n1083) );
NAND2_X1 U1025 ( .A1(n1143), .A2(n1260), .ZN(n1323) );
AND2_X1 U1026 ( .A1(n1325), .A2(n1324), .ZN(n1260) );
NAND2_X1 U1027 ( .A1(G237), .A2(G234), .ZN(n1324) );
XOR2_X1 U1028 ( .A(n1277), .B(KEYINPUT21), .Z(n1325) );
NOR2_X1 U1029 ( .A1(G898), .A2(n1051), .ZN(n1143) );
NOR2_X1 U1030 ( .A1(n1082), .A2(n1081), .ZN(n1225) );
INV_X1 U1031 ( .A(n1251), .ZN(n1081) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1326), .ZN(n1251) );
XNOR2_X1 U1033 ( .A(n1327), .B(n1195), .ZN(n1082) );
NAND2_X1 U1034 ( .A1(G210), .A2(n1326), .ZN(n1195) );
NAND2_X1 U1035 ( .A1(n1292), .A2(n1277), .ZN(n1326) );
NAND2_X1 U1036 ( .A1(n1328), .A2(n1277), .ZN(n1327) );
INV_X1 U1037 ( .A(G902), .ZN(n1277) );
XOR2_X1 U1038 ( .A(n1230), .B(n1329), .Z(n1328) );
NAND3_X1 U1039 ( .A1(n1330), .A2(n1331), .A3(n1232), .ZN(n1329) );
OR2_X1 U1040 ( .A1(n1234), .A2(n1233), .ZN(n1232) );
NAND3_X1 U1041 ( .A1(KEYINPUT5), .A2(n1234), .A3(n1233), .ZN(n1331) );
NAND2_X1 U1042 ( .A1(G224), .A2(n1051), .ZN(n1234) );
OR2_X1 U1043 ( .A1(n1233), .A2(KEYINPUT5), .ZN(n1330) );
XOR2_X1 U1044 ( .A(n1332), .B(n1295), .Z(n1233) );
NOR2_X1 U1045 ( .A1(KEYINPUT18), .A2(n1333), .ZN(n1295) );
XOR2_X1 U1046 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1047 ( .A(KEYINPUT24), .B(G146), .Z(n1335) );
NOR2_X1 U1048 ( .A1(KEYINPUT33), .A2(n1241), .ZN(n1334) );
INV_X1 U1049 ( .A(G143), .ZN(n1241) );
XNOR2_X1 U1050 ( .A(G125), .B(G128), .ZN(n1332) );
NAND2_X1 U1051 ( .A1(n1138), .A2(n1336), .ZN(n1230) );
NAND2_X1 U1052 ( .A1(n1140), .A2(n1141), .ZN(n1336) );
OR2_X1 U1053 ( .A1(n1141), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U1054 ( .A(n1337), .B(n1338), .ZN(n1140) );
XOR2_X1 U1055 ( .A(G101), .B(n1339), .Z(n1338) );
XOR2_X1 U1056 ( .A(G116), .B(G113), .Z(n1339) );
XOR2_X1 U1057 ( .A(n1340), .B(n1319), .Z(n1337) );
XOR2_X1 U1058 ( .A(G104), .B(G107), .Z(n1319) );
NAND2_X1 U1059 ( .A1(KEYINPUT61), .A2(n1267), .ZN(n1340) );
INV_X1 U1060 ( .A(G119), .ZN(n1267) );
XOR2_X1 U1061 ( .A(G110), .B(n1341), .Z(n1141) );
NOR2_X1 U1062 ( .A1(KEYINPUT37), .A2(n1261), .ZN(n1341) );
INV_X1 U1063 ( .A(G122), .ZN(n1261) );
NOR2_X1 U1064 ( .A1(n1265), .A2(n1263), .ZN(n1061) );
XOR2_X1 U1065 ( .A(n1342), .B(n1093), .Z(n1263) );
NOR2_X1 U1066 ( .A1(n1156), .A2(G902), .ZN(n1093) );
XNOR2_X1 U1067 ( .A(n1343), .B(n1344), .ZN(n1156) );
XOR2_X1 U1068 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1069 ( .A(G143), .B(G128), .Z(n1346) );
NOR2_X1 U1070 ( .A1(KEYINPUT13), .A2(n1347), .ZN(n1345) );
XNOR2_X1 U1071 ( .A(G134), .B(KEYINPUT20), .ZN(n1347) );
XNOR2_X1 U1072 ( .A(n1348), .B(n1349), .ZN(n1343) );
NAND2_X1 U1073 ( .A1(KEYINPUT4), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1074 ( .A(G107), .B(n1351), .Z(n1350) );
XOR2_X1 U1075 ( .A(G122), .B(G116), .Z(n1351) );
NAND4_X1 U1076 ( .A1(KEYINPUT17), .A2(G217), .A3(G234), .A4(n1051), .ZN(n1348) );
NAND2_X1 U1077 ( .A1(KEYINPUT62), .A2(n1160), .ZN(n1342) );
INV_X1 U1078 ( .A(G478), .ZN(n1160) );
INV_X1 U1079 ( .A(n1270), .ZN(n1265) );
NOR2_X1 U1080 ( .A1(n1352), .A2(n1099), .ZN(n1270) );
NOR2_X1 U1081 ( .A1(n1102), .A2(G475), .ZN(n1099) );
INV_X1 U1082 ( .A(n1353), .ZN(n1102) );
XNOR2_X1 U1083 ( .A(KEYINPUT59), .B(n1354), .ZN(n1352) );
NOR2_X1 U1084 ( .A1(n1353), .A2(n1355), .ZN(n1354) );
XNOR2_X1 U1085 ( .A(G475), .B(KEYINPUT8), .ZN(n1355) );
NOR2_X1 U1086 ( .A1(n1164), .A2(G902), .ZN(n1353) );
XOR2_X1 U1087 ( .A(n1356), .B(n1357), .Z(n1164) );
XOR2_X1 U1088 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1089 ( .A(G122), .B(G104), .Z(n1359) );
XOR2_X1 U1090 ( .A(KEYINPUT28), .B(G131), .Z(n1358) );
XOR2_X1 U1091 ( .A(n1360), .B(n1361), .Z(n1356) );
XNOR2_X1 U1092 ( .A(n1317), .B(n1120), .ZN(n1361) );
XNOR2_X1 U1093 ( .A(G140), .B(G125), .ZN(n1120) );
XOR2_X1 U1094 ( .A(G143), .B(G146), .Z(n1317) );
XOR2_X1 U1095 ( .A(n1362), .B(n1363), .Z(n1360) );
AND3_X1 U1096 ( .A1(G214), .A2(n1051), .A3(n1292), .ZN(n1363) );
INV_X1 U1097 ( .A(G237), .ZN(n1292) );
INV_X1 U1098 ( .A(G953), .ZN(n1051) );
NAND2_X1 U1099 ( .A1(KEYINPUT63), .A2(G113), .ZN(n1362) );
endmodule


