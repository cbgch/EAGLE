//Key = 1101100101110001000000001110010101011010110101111000101101101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374;

XOR2_X1 U747 ( .A(n1050), .B(n1051), .Z(G9) );
XOR2_X1 U748 ( .A(KEYINPUT54), .B(G107), .Z(n1051) );
NOR2_X1 U749 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND3_X1 U751 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1054) );
NAND2_X1 U752 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U753 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND4_X1 U754 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
OR2_X1 U755 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U756 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U758 ( .A1(n1065), .A2(n1074), .A3(n1064), .ZN(n1073) );
NAND2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U760 ( .A1(n1066), .A2(n1077), .ZN(n1072) );
NAND2_X1 U761 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U762 ( .A1(n1064), .A2(n1080), .ZN(n1079) );
NAND2_X1 U763 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U764 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1085), .ZN(n1078) );
NAND2_X1 U766 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U767 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
INV_X1 U768 ( .A(n1090), .ZN(n1060) );
AND3_X1 U769 ( .A1(n1057), .A2(n1058), .A3(n1091), .ZN(n1052) );
NAND4_X1 U770 ( .A1(n1070), .A2(n1066), .A3(n1092), .A4(n1093), .ZN(n1057) );
NOR3_X1 U771 ( .A1(n1094), .A2(n1083), .A3(n1088), .ZN(n1093) );
XOR2_X1 U772 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U773 ( .A(KEYINPUT26), .B(n1097), .Z(n1096) );
XOR2_X1 U774 ( .A(n1098), .B(n1099), .Z(n1092) );
XOR2_X1 U775 ( .A(KEYINPUT34), .B(G469), .Z(n1099) );
XOR2_X1 U776 ( .A(n1100), .B(n1101), .Z(G72) );
NOR2_X1 U777 ( .A1(n1102), .A2(n1058), .ZN(n1101) );
AND2_X1 U778 ( .A1(G227), .A2(G900), .ZN(n1102) );
NAND2_X1 U779 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U780 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U781 ( .A(n1107), .B(KEYINPUT37), .Z(n1103) );
OR2_X1 U782 ( .A1(n1106), .A2(n1105), .ZN(n1107) );
AND3_X1 U783 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1105) );
XOR2_X1 U784 ( .A(KEYINPUT60), .B(n1111), .Z(n1110) );
NOR2_X1 U785 ( .A1(G900), .A2(n1058), .ZN(n1111) );
NAND3_X1 U786 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1109) );
XOR2_X1 U787 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1108) );
NAND2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1118) );
XNOR2_X1 U790 ( .A(KEYINPUT1), .B(n1119), .ZN(n1112) );
NAND2_X1 U791 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U792 ( .A(n1122), .B(KEYINPUT3), .Z(n1120) );
XOR2_X1 U793 ( .A(n1116), .B(n1123), .Z(n1117) );
INV_X1 U794 ( .A(n1115), .ZN(n1123) );
XNOR2_X1 U795 ( .A(n1124), .B(n1125), .ZN(n1115) );
NOR2_X1 U796 ( .A1(G134), .A2(KEYINPUT32), .ZN(n1125) );
NAND2_X1 U797 ( .A1(n1126), .A2(n1055), .ZN(n1106) );
XOR2_X1 U798 ( .A(n1058), .B(KEYINPUT17), .Z(n1126) );
XOR2_X1 U799 ( .A(n1127), .B(n1128), .Z(G69) );
NOR2_X1 U800 ( .A1(n1129), .A2(n1058), .ZN(n1128) );
NOR2_X1 U801 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U802 ( .A1(n1132), .A2(n1133), .ZN(n1127) );
NAND2_X1 U803 ( .A1(KEYINPUT59), .A2(n1134), .ZN(n1133) );
XOR2_X1 U804 ( .A(n1135), .B(n1136), .Z(n1132) );
AND2_X1 U805 ( .A1(n1056), .A2(n1058), .ZN(n1136) );
OR2_X1 U806 ( .A1(n1134), .A2(KEYINPUT59), .ZN(n1135) );
NAND2_X1 U807 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND2_X1 U808 ( .A1(G953), .A2(n1131), .ZN(n1138) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1137) );
NOR2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XNOR2_X1 U811 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U812 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U813 ( .A(KEYINPUT15), .B(G217), .Z(n1146) );
NOR2_X1 U814 ( .A1(n1141), .A2(n1147), .ZN(G63) );
XOR2_X1 U815 ( .A(n1148), .B(n1149), .Z(n1147) );
AND2_X1 U816 ( .A1(G478), .A2(n1150), .ZN(n1148) );
NOR2_X1 U817 ( .A1(n1151), .A2(n1152), .ZN(G60) );
XOR2_X1 U818 ( .A(KEYINPUT21), .B(n1141), .Z(n1152) );
XOR2_X1 U819 ( .A(n1153), .B(n1154), .Z(n1151) );
AND2_X1 U820 ( .A1(G475), .A2(n1150), .ZN(n1153) );
XNOR2_X1 U821 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1156), .ZN(G57) );
XOR2_X1 U823 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U824 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U825 ( .A1(G472), .A2(n1150), .ZN(n1159) );
XOR2_X1 U826 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U827 ( .A(G101), .B(n1163), .Z(n1162) );
NOR2_X1 U828 ( .A1(KEYINPUT27), .A2(n1164), .ZN(n1161) );
NOR3_X1 U829 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(G54) );
AND2_X1 U830 ( .A1(KEYINPUT9), .A2(n1141), .ZN(n1167) );
NOR3_X1 U831 ( .A1(KEYINPUT9), .A2(n1058), .A3(n1091), .ZN(n1166) );
INV_X1 U832 ( .A(G952), .ZN(n1091) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1165) );
XNOR2_X1 U834 ( .A(n1170), .B(n1171), .ZN(n1169) );
XNOR2_X1 U835 ( .A(n1172), .B(n1116), .ZN(n1170) );
XOR2_X1 U836 ( .A(n1173), .B(n1174), .Z(n1168) );
XNOR2_X1 U837 ( .A(KEYINPUT16), .B(n1175), .ZN(n1174) );
XOR2_X1 U838 ( .A(n1176), .B(n1177), .Z(n1173) );
AND2_X1 U839 ( .A1(G469), .A2(n1150), .ZN(n1177) );
NAND2_X1 U840 ( .A1(KEYINPUT58), .A2(n1178), .ZN(n1176) );
NOR2_X1 U841 ( .A1(n1141), .A2(n1179), .ZN(G51) );
XOR2_X1 U842 ( .A(n1180), .B(KEYINPUT31), .Z(n1179) );
NAND2_X1 U843 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND3_X1 U844 ( .A1(n1150), .A2(n1097), .A3(n1183), .ZN(n1182) );
XOR2_X1 U845 ( .A(n1184), .B(KEYINPUT28), .Z(n1181) );
NAND2_X1 U846 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U847 ( .A1(n1150), .A2(n1097), .ZN(n1186) );
INV_X1 U848 ( .A(n1145), .ZN(n1150) );
NAND2_X1 U849 ( .A1(G902), .A2(n1187), .ZN(n1145) );
OR2_X1 U850 ( .A1(n1056), .A2(n1055), .ZN(n1187) );
NAND4_X1 U851 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1055) );
AND4_X1 U852 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NAND2_X1 U853 ( .A1(KEYINPUT43), .A2(n1196), .ZN(n1190) );
NAND2_X1 U854 ( .A1(n1064), .A2(n1197), .ZN(n1188) );
NAND2_X1 U855 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U856 ( .A1(n1068), .A2(n1200), .ZN(n1199) );
NAND2_X1 U857 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
OR4_X1 U858 ( .A1(n1203), .A2(n1076), .A3(n1081), .A4(KEYINPUT43), .ZN(n1202) );
NAND2_X1 U859 ( .A1(n1204), .A2(n1070), .ZN(n1198) );
NAND4_X1 U860 ( .A1(n1205), .A2(n1050), .A3(n1206), .A4(n1207), .ZN(n1056) );
AND4_X1 U861 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1155), .ZN(n1207) );
NAND3_X1 U862 ( .A1(n1211), .A2(n1066), .A3(n1068), .ZN(n1155) );
NOR3_X1 U863 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1206) );
NOR4_X1 U864 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
INV_X1 U865 ( .A(KEYINPUT52), .ZN(n1215) );
NOR3_X1 U866 ( .A1(KEYINPUT52), .A2(n1219), .A3(n1086), .ZN(n1213) );
NOR4_X1 U867 ( .A1(n1220), .A2(n1217), .A3(n1221), .A4(n1216), .ZN(n1219) );
NAND3_X1 U868 ( .A1(n1069), .A2(n1066), .A3(n1211), .ZN(n1050) );
INV_X1 U869 ( .A(n1183), .ZN(n1185) );
XOR2_X1 U870 ( .A(n1222), .B(n1223), .Z(n1183) );
NOR2_X1 U871 ( .A1(n1058), .A2(G952), .ZN(n1141) );
XOR2_X1 U872 ( .A(n1224), .B(n1189), .Z(G48) );
NAND3_X1 U873 ( .A1(n1068), .A2(n1225), .A3(n1204), .ZN(n1189) );
XOR2_X1 U874 ( .A(n1226), .B(n1195), .Z(G45) );
NAND4_X1 U875 ( .A1(n1227), .A2(n1225), .A3(n1228), .A4(n1229), .ZN(n1195) );
NAND2_X1 U876 ( .A1(n1230), .A2(n1231), .ZN(G42) );
NAND2_X1 U877 ( .A1(G140), .A2(n1232), .ZN(n1231) );
NAND2_X1 U878 ( .A1(n1196), .A2(n1233), .ZN(n1232) );
OR2_X1 U879 ( .A1(n1234), .A2(KEYINPUT11), .ZN(n1233) );
NAND3_X1 U880 ( .A1(n1235), .A2(n1236), .A3(KEYINPUT11), .ZN(n1230) );
NAND2_X1 U881 ( .A1(n1196), .A2(n1234), .ZN(n1236) );
INV_X1 U882 ( .A(KEYINPUT0), .ZN(n1234) );
NAND2_X1 U883 ( .A1(KEYINPUT0), .A2(n1237), .ZN(n1235) );
NAND2_X1 U884 ( .A1(n1196), .A2(n1122), .ZN(n1237) );
AND4_X1 U885 ( .A1(n1064), .A2(n1068), .A3(n1238), .A4(n1239), .ZN(n1196) );
NOR2_X1 U886 ( .A1(n1240), .A2(n1081), .ZN(n1238) );
XOR2_X1 U887 ( .A(n1241), .B(n1242), .Z(G39) );
NOR2_X1 U888 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U889 ( .A(KEYINPUT40), .B(n1245), .Z(n1244) );
NOR2_X1 U890 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U891 ( .A(KEYINPUT33), .B(n1070), .Z(n1247) );
INV_X1 U892 ( .A(n1204), .ZN(n1246) );
XNOR2_X1 U893 ( .A(G137), .B(KEYINPUT46), .ZN(n1241) );
XNOR2_X1 U894 ( .A(G134), .B(n1194), .ZN(G36) );
NAND3_X1 U895 ( .A1(n1227), .A2(n1069), .A3(n1064), .ZN(n1194) );
XNOR2_X1 U896 ( .A(G131), .B(n1248), .ZN(G33) );
NAND2_X1 U897 ( .A1(n1064), .A2(n1249), .ZN(n1248) );
XOR2_X1 U898 ( .A(KEYINPUT13), .B(n1250), .Z(n1249) );
NOR2_X1 U899 ( .A1(n1251), .A2(n1201), .ZN(n1250) );
INV_X1 U900 ( .A(n1227), .ZN(n1201) );
NOR3_X1 U901 ( .A1(n1081), .A2(n1240), .A3(n1075), .ZN(n1227) );
INV_X1 U902 ( .A(n1252), .ZN(n1075) );
INV_X1 U903 ( .A(n1243), .ZN(n1064) );
NAND2_X1 U904 ( .A1(n1089), .A2(n1253), .ZN(n1243) );
XOR2_X1 U905 ( .A(n1254), .B(n1193), .Z(G30) );
NAND3_X1 U906 ( .A1(n1069), .A2(n1225), .A3(n1204), .ZN(n1193) );
NOR3_X1 U907 ( .A1(n1081), .A2(n1240), .A3(n1216), .ZN(n1204) );
XOR2_X1 U908 ( .A(n1210), .B(n1255), .Z(G3) );
NAND2_X1 U909 ( .A1(KEYINPUT57), .A2(G101), .ZN(n1255) );
NAND3_X1 U910 ( .A1(n1070), .A2(n1211), .A3(n1252), .ZN(n1210) );
XOR2_X1 U911 ( .A(n1121), .B(n1256), .Z(G27) );
NAND2_X1 U912 ( .A1(KEYINPUT24), .A2(n1257), .ZN(n1256) );
INV_X1 U913 ( .A(n1192), .ZN(n1257) );
NAND3_X1 U914 ( .A1(n1068), .A2(n1065), .A3(n1258), .ZN(n1192) );
NOR3_X1 U915 ( .A1(n1076), .A2(n1240), .A3(n1086), .ZN(n1258) );
INV_X1 U916 ( .A(n1203), .ZN(n1240) );
NAND2_X1 U917 ( .A1(n1090), .A2(n1259), .ZN(n1203) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1261), .ZN(n1259) );
INV_X1 U919 ( .A(G900), .ZN(n1261) );
INV_X1 U920 ( .A(n1221), .ZN(n1065) );
XNOR2_X1 U921 ( .A(G122), .B(n1209), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1262), .A2(n1066), .A3(n1228), .A4(n1229), .ZN(n1209) );
NOR2_X1 U923 ( .A1(n1263), .A2(n1264), .ZN(n1066) );
XOR2_X1 U924 ( .A(G119), .B(n1265), .Z(G21) );
NOR4_X1 U925 ( .A1(KEYINPUT51), .A2(n1217), .A3(n1218), .A4(n1266), .ZN(n1265) );
XNOR2_X1 U926 ( .A(KEYINPUT36), .B(n1216), .ZN(n1266) );
NAND2_X1 U927 ( .A1(n1264), .A2(n1263), .ZN(n1216) );
INV_X1 U928 ( .A(n1267), .ZN(n1264) );
INV_X1 U929 ( .A(n1262), .ZN(n1218) );
INV_X1 U930 ( .A(n1070), .ZN(n1217) );
XOR2_X1 U931 ( .A(G116), .B(n1212), .Z(G18) );
AND3_X1 U932 ( .A1(n1262), .A2(n1069), .A3(n1252), .ZN(n1212) );
NOR2_X1 U933 ( .A1(n1229), .A2(n1268), .ZN(n1069) );
XNOR2_X1 U934 ( .A(G113), .B(n1205), .ZN(G15) );
NAND3_X1 U935 ( .A1(n1252), .A2(n1262), .A3(n1068), .ZN(n1205) );
INV_X1 U936 ( .A(n1251), .ZN(n1068) );
NAND2_X1 U937 ( .A1(n1268), .A2(n1229), .ZN(n1251) );
NOR3_X1 U938 ( .A1(n1086), .A2(n1220), .A3(n1221), .ZN(n1262) );
NAND2_X1 U939 ( .A1(n1084), .A2(n1269), .ZN(n1221) );
XNOR2_X1 U940 ( .A(n1270), .B(KEYINPUT23), .ZN(n1084) );
NOR2_X1 U941 ( .A1(n1263), .A2(n1267), .ZN(n1252) );
XOR2_X1 U942 ( .A(n1271), .B(n1272), .Z(G12) );
NAND2_X1 U943 ( .A1(KEYINPUT47), .A2(n1273), .ZN(n1272) );
INV_X1 U944 ( .A(n1208), .ZN(n1273) );
NAND3_X1 U945 ( .A1(n1070), .A2(n1211), .A3(n1239), .ZN(n1208) );
INV_X1 U946 ( .A(n1076), .ZN(n1239) );
NAND2_X1 U947 ( .A1(n1267), .A2(n1263), .ZN(n1076) );
NAND3_X1 U948 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1263) );
OR2_X1 U949 ( .A1(n1277), .A2(n1143), .ZN(n1276) );
NAND3_X1 U950 ( .A1(n1143), .A2(n1277), .A3(n1278), .ZN(n1275) );
NAND2_X1 U951 ( .A1(G217), .A2(n1279), .ZN(n1277) );
XNOR2_X1 U952 ( .A(n1280), .B(n1281), .ZN(n1143) );
XOR2_X1 U953 ( .A(G110), .B(n1282), .Z(n1281) );
XOR2_X1 U954 ( .A(G137), .B(G119), .Z(n1282) );
XNOR2_X1 U955 ( .A(n1283), .B(n1284), .ZN(n1280) );
XOR2_X1 U956 ( .A(n1285), .B(n1286), .Z(n1283) );
NOR2_X1 U957 ( .A1(KEYINPUT14), .A2(G128), .ZN(n1286) );
NAND2_X1 U958 ( .A1(n1287), .A2(G221), .ZN(n1285) );
NAND2_X1 U959 ( .A1(G217), .A2(G902), .ZN(n1274) );
XOR2_X1 U960 ( .A(n1288), .B(G472), .Z(n1267) );
NAND2_X1 U961 ( .A1(n1289), .A2(n1278), .ZN(n1288) );
XOR2_X1 U962 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U963 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U964 ( .A(KEYINPUT12), .B(n1294), .Z(n1293) );
AND2_X1 U965 ( .A1(n1160), .A2(n1164), .ZN(n1294) );
NOR2_X1 U966 ( .A1(n1164), .A2(n1160), .ZN(n1292) );
XNOR2_X1 U967 ( .A(n1295), .B(n1178), .ZN(n1160) );
XNOR2_X1 U968 ( .A(n1296), .B(n1297), .ZN(n1164) );
NOR2_X1 U969 ( .A1(KEYINPUT56), .A2(n1298), .ZN(n1290) );
XOR2_X1 U970 ( .A(n1163), .B(n1299), .Z(n1298) );
NOR2_X1 U971 ( .A1(KEYINPUT50), .A2(n1300), .ZN(n1299) );
XOR2_X1 U972 ( .A(n1301), .B(KEYINPUT38), .Z(n1300) );
AND3_X1 U973 ( .A1(n1302), .A2(n1058), .A3(G210), .ZN(n1163) );
NOR3_X1 U974 ( .A1(n1081), .A2(n1220), .A3(n1086), .ZN(n1211) );
INV_X1 U975 ( .A(n1225), .ZN(n1086) );
NOR2_X1 U976 ( .A1(n1089), .A2(n1088), .ZN(n1225) );
INV_X1 U977 ( .A(n1253), .ZN(n1088) );
NAND2_X1 U978 ( .A1(G214), .A2(n1303), .ZN(n1253) );
XNOR2_X1 U979 ( .A(n1095), .B(n1304), .ZN(n1089) );
NOR2_X1 U980 ( .A1(n1097), .A2(KEYINPUT22), .ZN(n1304) );
AND2_X1 U981 ( .A1(G210), .A2(n1303), .ZN(n1097) );
NAND2_X1 U982 ( .A1(n1302), .A2(n1278), .ZN(n1303) );
NAND2_X1 U983 ( .A1(n1305), .A2(n1278), .ZN(n1095) );
XOR2_X1 U984 ( .A(n1306), .B(n1222), .Z(n1305) );
XOR2_X1 U985 ( .A(n1307), .B(n1308), .Z(n1222) );
XOR2_X1 U986 ( .A(n1309), .B(n1140), .Z(n1308) );
XOR2_X1 U987 ( .A(n1310), .B(n1311), .Z(n1140) );
XOR2_X1 U988 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U989 ( .A(KEYINPUT30), .B(G110), .Z(n1313) );
XOR2_X1 U990 ( .A(KEYINPUT55), .B(KEYINPUT39), .Z(n1312) );
XOR2_X1 U991 ( .A(n1314), .B(n1315), .Z(n1310) );
XNOR2_X1 U992 ( .A(G107), .B(n1316), .ZN(n1314) );
NOR2_X1 U993 ( .A1(KEYINPUT6), .A2(n1301), .ZN(n1316) );
INV_X1 U994 ( .A(G101), .ZN(n1301) );
NAND2_X1 U995 ( .A1(KEYINPUT45), .A2(n1139), .ZN(n1309) );
NAND2_X1 U996 ( .A1(n1317), .A2(n1318), .ZN(n1139) );
NAND2_X1 U997 ( .A1(n1319), .A2(n1296), .ZN(n1318) );
INV_X1 U998 ( .A(n1297), .ZN(n1319) );
NAND2_X1 U999 ( .A1(n1320), .A2(n1297), .ZN(n1317) );
XNOR2_X1 U1000 ( .A(KEYINPUT61), .B(n1296), .ZN(n1320) );
XNOR2_X1 U1001 ( .A(G113), .B(G119), .ZN(n1296) );
XOR2_X1 U1002 ( .A(n1295), .B(G125), .Z(n1307) );
NAND3_X1 U1003 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(n1295) );
NAND2_X1 U1004 ( .A1(G128), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1005 ( .A1(n1325), .A2(n1326), .ZN(n1322) );
INV_X1 U1006 ( .A(KEYINPUT25), .ZN(n1326) );
NAND2_X1 U1007 ( .A1(n1327), .A2(n1254), .ZN(n1325) );
XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n1324), .ZN(n1327) );
NAND2_X1 U1009 ( .A1(KEYINPUT25), .A2(n1328), .ZN(n1321) );
NAND2_X1 U1010 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1011 ( .A1(KEYINPUT49), .A2(n1324), .ZN(n1330) );
OR3_X1 U1012 ( .A1(G128), .A2(KEYINPUT49), .A3(n1324), .ZN(n1329) );
AND2_X1 U1013 ( .A1(n1331), .A2(n1332), .ZN(n1324) );
NAND2_X1 U1014 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
INV_X1 U1015 ( .A(KEYINPUT44), .ZN(n1334) );
NAND3_X1 U1016 ( .A1(G143), .A2(n1224), .A3(KEYINPUT44), .ZN(n1331) );
NAND2_X1 U1017 ( .A1(KEYINPUT35), .A2(n1223), .ZN(n1306) );
NOR2_X1 U1018 ( .A1(n1130), .A2(G953), .ZN(n1223) );
INV_X1 U1019 ( .A(G224), .ZN(n1130) );
AND2_X1 U1020 ( .A1(n1090), .A2(n1335), .ZN(n1220) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1131), .ZN(n1335) );
INV_X1 U1022 ( .A(G898), .ZN(n1131) );
NAND3_X1 U1023 ( .A1(n1260), .A2(n1058), .A3(G952), .ZN(n1090) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1260) );
NAND2_X1 U1025 ( .A1(n1270), .A2(n1269), .ZN(n1081) );
XOR2_X1 U1026 ( .A(n1083), .B(KEYINPUT4), .Z(n1269) );
AND2_X1 U1027 ( .A1(G221), .A2(n1336), .ZN(n1083) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1278), .ZN(n1336) );
XOR2_X1 U1029 ( .A(n1098), .B(n1337), .Z(n1270) );
NOR2_X1 U1030 ( .A1(G469), .A2(KEYINPUT8), .ZN(n1337) );
NAND2_X1 U1031 ( .A1(n1338), .A2(n1278), .ZN(n1098) );
INV_X1 U1032 ( .A(G902), .ZN(n1278) );
XOR2_X1 U1033 ( .A(n1339), .B(n1172), .Z(n1338) );
XNOR2_X1 U1034 ( .A(n1271), .B(G140), .ZN(n1172) );
XNOR2_X1 U1035 ( .A(n1340), .B(n1341), .ZN(n1339) );
NOR2_X1 U1036 ( .A1(KEYINPUT53), .A2(n1342), .ZN(n1341) );
XNOR2_X1 U1037 ( .A(n1116), .B(n1343), .ZN(n1342) );
XNOR2_X1 U1038 ( .A(n1344), .B(n1345), .ZN(n1343) );
NOR2_X1 U1039 ( .A1(KEYINPUT42), .A2(n1171), .ZN(n1345) );
XOR2_X1 U1040 ( .A(n1346), .B(n1347), .Z(n1171) );
XOR2_X1 U1041 ( .A(G101), .B(n1348), .Z(n1347) );
NOR2_X1 U1042 ( .A1(G107), .A2(KEYINPUT5), .ZN(n1348) );
XNOR2_X1 U1043 ( .A(G104), .B(KEYINPUT30), .ZN(n1346) );
NAND2_X1 U1044 ( .A1(KEYINPUT29), .A2(n1178), .ZN(n1344) );
XNOR2_X1 U1045 ( .A(n1349), .B(n1350), .ZN(n1178) );
XOR2_X1 U1046 ( .A(KEYINPUT7), .B(KEYINPUT10), .Z(n1350) );
XNOR2_X1 U1047 ( .A(G134), .B(n1124), .ZN(n1349) );
XOR2_X1 U1048 ( .A(G131), .B(G137), .Z(n1124) );
XNOR2_X1 U1049 ( .A(n1254), .B(n1351), .ZN(n1116) );
NOR2_X1 U1050 ( .A1(KEYINPUT2), .A2(n1333), .ZN(n1351) );
XOR2_X1 U1051 ( .A(n1226), .B(G146), .Z(n1333) );
INV_X1 U1052 ( .A(G128), .ZN(n1254) );
NOR2_X1 U1053 ( .A1(KEYINPUT63), .A2(n1175), .ZN(n1340) );
NAND2_X1 U1054 ( .A1(G227), .A2(n1058), .ZN(n1175) );
NOR2_X1 U1055 ( .A1(n1228), .A2(n1229), .ZN(n1070) );
XNOR2_X1 U1056 ( .A(n1352), .B(n1353), .ZN(n1229) );
XOR2_X1 U1057 ( .A(KEYINPUT20), .B(G475), .Z(n1353) );
OR2_X1 U1058 ( .A1(n1154), .A2(G902), .ZN(n1352) );
XOR2_X1 U1059 ( .A(n1315), .B(n1354), .Z(n1154) );
XOR2_X1 U1060 ( .A(G113), .B(n1355), .Z(n1354) );
NOR2_X1 U1061 ( .A1(KEYINPUT18), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1062 ( .A(n1357), .B(n1284), .Z(n1356) );
NAND2_X1 U1063 ( .A1(n1358), .A2(n1359), .ZN(n1284) );
NAND2_X1 U1064 ( .A1(n1360), .A2(n1224), .ZN(n1359) );
INV_X1 U1065 ( .A(G146), .ZN(n1224) );
NAND2_X1 U1066 ( .A1(n1113), .A2(n1361), .ZN(n1360) );
NAND2_X1 U1067 ( .A1(G140), .A2(n1121), .ZN(n1361) );
NAND2_X1 U1068 ( .A1(G125), .A2(n1122), .ZN(n1113) );
INV_X1 U1069 ( .A(G140), .ZN(n1122) );
NAND2_X1 U1070 ( .A1(G146), .A2(n1362), .ZN(n1358) );
XOR2_X1 U1071 ( .A(n1121), .B(G140), .Z(n1362) );
INV_X1 U1072 ( .A(G125), .ZN(n1121) );
NAND2_X1 U1073 ( .A1(n1363), .A2(KEYINPUT48), .ZN(n1357) );
XOR2_X1 U1074 ( .A(n1364), .B(n1365), .Z(n1363) );
AND3_X1 U1075 ( .A1(G214), .A2(n1058), .A3(n1302), .ZN(n1365) );
INV_X1 U1076 ( .A(G237), .ZN(n1302) );
INV_X1 U1077 ( .A(G953), .ZN(n1058) );
XOR2_X1 U1078 ( .A(G131), .B(n1226), .Z(n1364) );
INV_X1 U1079 ( .A(G143), .ZN(n1226) );
XOR2_X1 U1080 ( .A(G104), .B(G122), .Z(n1315) );
INV_X1 U1081 ( .A(n1268), .ZN(n1228) );
XOR2_X1 U1082 ( .A(n1366), .B(G478), .Z(n1268) );
OR2_X1 U1083 ( .A1(n1149), .A2(G902), .ZN(n1366) );
XNOR2_X1 U1084 ( .A(n1367), .B(n1368), .ZN(n1149) );
XOR2_X1 U1085 ( .A(n1297), .B(n1369), .Z(n1368) );
XOR2_X1 U1086 ( .A(n1370), .B(n1371), .Z(n1369) );
NOR2_X1 U1087 ( .A1(KEYINPUT19), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1088 ( .A(G143), .B(G128), .Z(n1372) );
NAND2_X1 U1089 ( .A1(G217), .A2(n1287), .ZN(n1370) );
NOR2_X1 U1090 ( .A1(n1279), .A2(G953), .ZN(n1287) );
INV_X1 U1091 ( .A(G234), .ZN(n1279) );
XNOR2_X1 U1092 ( .A(G116), .B(KEYINPUT41), .ZN(n1297) );
XOR2_X1 U1093 ( .A(n1373), .B(n1374), .Z(n1367) );
NOR2_X1 U1094 ( .A1(KEYINPUT62), .A2(G107), .ZN(n1374) );
XNOR2_X1 U1095 ( .A(G122), .B(G134), .ZN(n1373) );
INV_X1 U1096 ( .A(G110), .ZN(n1271) );
endmodule


