//Key = 1010111001010001000100111111111011111001001100001011001111000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;

XNOR2_X1 U692 ( .A(n953), .B(n954), .ZN(G9) );
NAND2_X1 U693 ( .A1(KEYINPUT26), .A2(G107), .ZN(n954) );
NAND4_X1 U694 ( .A1(n955), .A2(n956), .A3(n957), .A4(n958), .ZN(G75) );
NAND4_X1 U695 ( .A1(n959), .A2(n960), .A3(n961), .A4(n962), .ZN(n957) );
NOR4_X1 U696 ( .A1(n963), .A2(n964), .A3(n965), .A4(n966), .ZN(n962) );
XNOR2_X1 U697 ( .A(KEYINPUT46), .B(n967), .ZN(n966) );
XOR2_X1 U698 ( .A(n968), .B(n969), .Z(n965) );
NAND2_X1 U699 ( .A1(n970), .A2(n971), .ZN(n969) );
NAND2_X1 U700 ( .A1(n972), .A2(n973), .ZN(n964) );
AND3_X1 U701 ( .A1(n974), .A2(n975), .A3(n976), .ZN(n961) );
NAND3_X1 U702 ( .A1(n977), .A2(n978), .A3(G210), .ZN(n959) );
NAND2_X1 U703 ( .A1(n979), .A2(n980), .ZN(n956) );
NAND2_X1 U704 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND3_X1 U705 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
NAND3_X1 U706 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n984) );
NAND2_X1 U707 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND3_X1 U708 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NAND2_X1 U709 ( .A1(n994), .A2(n995), .ZN(n992) );
INV_X1 U710 ( .A(KEYINPUT9), .ZN(n995) );
NAND3_X1 U711 ( .A1(n996), .A2(n997), .A3(KEYINPUT9), .ZN(n991) );
NAND2_X1 U712 ( .A1(n994), .A2(n998), .ZN(n987) );
NAND2_X1 U713 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U714 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
OR3_X1 U715 ( .A1(n1002), .A2(n1003), .A3(n994), .ZN(n986) );
INV_X1 U716 ( .A(KEYINPUT20), .ZN(n1002) );
NAND3_X1 U717 ( .A1(n989), .A2(n1004), .A3(n994), .ZN(n981) );
NAND2_X1 U718 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U719 ( .A1(n985), .A2(n1007), .ZN(n1006) );
OR2_X1 U720 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U721 ( .A1(n983), .A2(n1010), .ZN(n1005) );
NAND2_X1 U722 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U723 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
XNOR2_X1 U724 ( .A(KEYINPUT14), .B(n975), .ZN(n1014) );
INV_X1 U725 ( .A(n1015), .ZN(n979) );
INV_X1 U726 ( .A(n1016), .ZN(n955) );
XOR2_X1 U727 ( .A(n1017), .B(n1018), .Z(G72) );
XOR2_X1 U728 ( .A(n1019), .B(n1020), .Z(n1018) );
NAND2_X1 U729 ( .A1(G953), .A2(n1021), .ZN(n1020) );
NAND2_X1 U730 ( .A1(G900), .A2(G227), .ZN(n1021) );
NAND2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NAND2_X1 U732 ( .A1(G953), .A2(n1024), .ZN(n1023) );
XOR2_X1 U733 ( .A(n1025), .B(n1026), .Z(n1022) );
XOR2_X1 U734 ( .A(n1027), .B(n1028), .Z(n1026) );
XOR2_X1 U735 ( .A(n1029), .B(G131), .Z(n1028) );
XOR2_X1 U736 ( .A(n1030), .B(n1031), .Z(n1025) );
XNOR2_X1 U737 ( .A(KEYINPUT5), .B(KEYINPUT37), .ZN(n1031) );
NOR2_X1 U738 ( .A1(n1032), .A2(G953), .ZN(n1017) );
XOR2_X1 U739 ( .A(n1033), .B(n1034), .Z(G69) );
NOR3_X1 U740 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U741 ( .A1(G953), .A2(n1038), .ZN(n1037) );
NOR2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
XNOR2_X1 U743 ( .A(KEYINPUT16), .B(n1041), .ZN(n1040) );
NOR2_X1 U744 ( .A1(G224), .A2(n958), .ZN(n1036) );
OR2_X1 U745 ( .A1(n1042), .A2(n1035), .ZN(n1033) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(G66) );
XOR2_X1 U747 ( .A(n1045), .B(n970), .Z(n1044) );
NAND3_X1 U748 ( .A1(n1046), .A2(n1016), .A3(n1047), .ZN(n1045) );
XOR2_X1 U749 ( .A(n971), .B(KEYINPUT50), .Z(n1047) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1048), .ZN(G63) );
XNOR2_X1 U751 ( .A(n1049), .B(n1050), .ZN(n1048) );
NOR3_X1 U752 ( .A1(n1051), .A2(KEYINPUT63), .A3(n1052), .ZN(n1050) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1053), .ZN(G60) );
XOR2_X1 U754 ( .A(n1054), .B(n1055), .Z(n1053) );
AND2_X1 U755 ( .A1(G475), .A2(n1056), .ZN(n1054) );
XNOR2_X1 U756 ( .A(n1057), .B(n1058), .ZN(G6) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
XOR2_X1 U758 ( .A(KEYINPUT8), .B(KEYINPUT13), .Z(n1060) );
NOR2_X1 U759 ( .A1(n1043), .A2(n1061), .ZN(G57) );
XOR2_X1 U760 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U761 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U762 ( .A(n1066), .B(n1067), .Z(n1062) );
XOR2_X1 U763 ( .A(KEYINPUT15), .B(n1068), .Z(n1067) );
AND2_X1 U764 ( .A1(G472), .A2(n1056), .ZN(n1068) );
NAND2_X1 U765 ( .A1(KEYINPUT4), .A2(n1069), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1043), .A2(n1070), .ZN(G54) );
XOR2_X1 U767 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U768 ( .A1(KEYINPUT47), .A2(n1073), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U770 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1074) );
XOR2_X1 U772 ( .A(KEYINPUT28), .B(KEYINPUT25), .Z(n1079) );
NAND2_X1 U773 ( .A1(n1056), .A2(G469), .ZN(n1071) );
INV_X1 U774 ( .A(n1051), .ZN(n1056) );
NOR2_X1 U775 ( .A1(n1043), .A2(n1080), .ZN(G51) );
XOR2_X1 U776 ( .A(n1081), .B(n1082), .Z(n1080) );
XNOR2_X1 U777 ( .A(n1083), .B(n1084), .ZN(n1082) );
XOR2_X1 U778 ( .A(n1085), .B(n1042), .Z(n1084) );
NAND2_X1 U779 ( .A1(KEYINPUT57), .A2(G125), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1081) );
XOR2_X1 U781 ( .A(KEYINPUT58), .B(n1088), .Z(n1087) );
NOR2_X1 U782 ( .A1(n1051), .A2(n1089), .ZN(n1088) );
XOR2_X1 U783 ( .A(KEYINPUT35), .B(G210), .Z(n1089) );
NAND2_X1 U784 ( .A1(G902), .A2(n1016), .ZN(n1051) );
NAND3_X1 U785 ( .A1(n1032), .A2(n1041), .A3(n1090), .ZN(n1016) );
INV_X1 U786 ( .A(n1039), .ZN(n1090) );
NAND4_X1 U787 ( .A1(n1058), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1039) );
NOR4_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n953), .A4(n1096), .ZN(n1093) );
AND3_X1 U789 ( .A1(n983), .A2(n1097), .A3(n1098), .ZN(n953) );
OR2_X1 U790 ( .A1(n1003), .A2(n1099), .ZN(n1092) );
NAND3_X1 U791 ( .A1(n983), .A2(n1097), .A3(n1001), .ZN(n1058) );
AND4_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1032) );
NOR4_X1 U793 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1103) );
NOR3_X1 U794 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1102) );
AND4_X1 U795 ( .A1(KEYINPUT49), .A2(n1111), .A3(n993), .A4(n1098), .ZN(n1110) );
NOR2_X1 U796 ( .A1(KEYINPUT49), .A2(n1112), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1108) );
XOR2_X1 U798 ( .A(KEYINPUT56), .B(n1115), .Z(n1114) );
NOR2_X1 U799 ( .A1(n958), .A2(G952), .ZN(n1043) );
XOR2_X1 U800 ( .A(n1100), .B(n1116), .Z(G48) );
XNOR2_X1 U801 ( .A(G146), .B(KEYINPUT45), .ZN(n1116) );
NAND3_X1 U802 ( .A1(n1001), .A2(n1117), .A3(n1111), .ZN(n1100) );
XOR2_X1 U803 ( .A(n1118), .B(n1101), .Z(G45) );
NAND4_X1 U804 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1101) );
NOR3_X1 U805 ( .A1(n1123), .A2(n1011), .A3(n993), .ZN(n1122) );
XOR2_X1 U806 ( .A(G140), .B(n1107), .Z(G42) );
AND3_X1 U807 ( .A1(n1001), .A2(n1009), .A3(n1124), .ZN(n1107) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(G39) );
NAND2_X1 U809 ( .A1(KEYINPUT24), .A2(n1106), .ZN(n1126) );
AND4_X1 U810 ( .A1(n1127), .A2(n1124), .A3(n989), .A4(n1128), .ZN(n1106) );
XOR2_X1 U811 ( .A(n1105), .B(n1129), .Z(G36) );
NOR2_X1 U812 ( .A1(KEYINPUT10), .A2(n1030), .ZN(n1129) );
AND3_X1 U813 ( .A1(n1008), .A2(n1098), .A3(n1124), .ZN(n1105) );
XOR2_X1 U814 ( .A(G131), .B(n1104), .Z(G33) );
AND3_X1 U815 ( .A1(n1001), .A2(n1008), .A3(n1124), .ZN(n1104) );
AND3_X1 U816 ( .A1(n1117), .A2(n1119), .A3(n985), .ZN(n1124) );
AND2_X1 U817 ( .A1(n1013), .A2(n1130), .ZN(n985) );
XNOR2_X1 U818 ( .A(KEYINPUT42), .B(n975), .ZN(n1130) );
INV_X1 U819 ( .A(n1131), .ZN(n1013) );
XOR2_X1 U820 ( .A(n1132), .B(n1112), .Z(G30) );
NAND3_X1 U821 ( .A1(n1098), .A2(n1117), .A3(n1111), .ZN(n1112) );
AND4_X1 U822 ( .A1(n1127), .A2(n1115), .A3(n1128), .A4(n1119), .ZN(n1111) );
INV_X1 U823 ( .A(n999), .ZN(n1098) );
XOR2_X1 U824 ( .A(n1133), .B(n1091), .Z(G3) );
NAND3_X1 U825 ( .A1(n1097), .A2(n989), .A3(n1008), .ZN(n1091) );
XOR2_X1 U826 ( .A(n1134), .B(n1135), .Z(G27) );
NOR2_X1 U827 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U828 ( .A(G125), .ZN(n1137) );
XNOR2_X1 U829 ( .A(KEYINPUT62), .B(KEYINPUT33), .ZN(n1136) );
NOR2_X1 U830 ( .A1(n1011), .A2(n1113), .ZN(n1134) );
NAND4_X1 U831 ( .A1(n1001), .A2(n994), .A3(n1009), .A4(n1119), .ZN(n1113) );
NAND2_X1 U832 ( .A1(n1015), .A2(n1138), .ZN(n1119) );
NAND4_X1 U833 ( .A1(G902), .A2(G953), .A3(n1139), .A4(n1024), .ZN(n1138) );
INV_X1 U834 ( .A(G900), .ZN(n1024) );
INV_X1 U835 ( .A(n1003), .ZN(n1001) );
XOR2_X1 U836 ( .A(G122), .B(n1095), .Z(G24) );
AND4_X1 U837 ( .A1(n994), .A2(n983), .A3(n1140), .A4(n1141), .ZN(n1095) );
NOR2_X1 U838 ( .A1(n1142), .A2(n972), .ZN(n1140) );
NOR2_X1 U839 ( .A1(n1128), .A2(n1127), .ZN(n983) );
XOR2_X1 U840 ( .A(G119), .B(n1143), .Z(G21) );
NOR2_X1 U841 ( .A1(KEYINPUT41), .A2(n1041), .ZN(n1143) );
NAND4_X1 U842 ( .A1(n1127), .A2(n994), .A3(n1144), .A4(n1141), .ZN(n1041) );
AND2_X1 U843 ( .A1(n1128), .A2(n989), .ZN(n1144) );
INV_X1 U844 ( .A(n1145), .ZN(n1128) );
NAND2_X1 U845 ( .A1(n1146), .A2(n1147), .ZN(G18) );
OR2_X1 U846 ( .A1(n1148), .A2(n1096), .ZN(n1147) );
XOR2_X1 U847 ( .A(n1149), .B(KEYINPUT12), .Z(n1146) );
NAND2_X1 U848 ( .A1(n1096), .A2(n1148), .ZN(n1149) );
INV_X1 U849 ( .A(G116), .ZN(n1148) );
NOR2_X1 U850 ( .A1(n1099), .A2(n999), .ZN(n1096) );
XOR2_X1 U851 ( .A(G113), .B(n1150), .Z(G15) );
NOR2_X1 U852 ( .A1(n1151), .A2(n1099), .ZN(n1150) );
NAND3_X1 U853 ( .A1(n994), .A2(n1141), .A3(n1008), .ZN(n1099) );
INV_X1 U854 ( .A(n1123), .ZN(n1008) );
NAND2_X1 U855 ( .A1(n1127), .A2(n1145), .ZN(n1123) );
NOR2_X1 U856 ( .A1(n1152), .A2(n996), .ZN(n994) );
INV_X1 U857 ( .A(n960), .ZN(n996) );
XOR2_X1 U858 ( .A(n1003), .B(KEYINPUT38), .Z(n1151) );
NAND2_X1 U859 ( .A1(n1153), .A2(n1121), .ZN(n1003) );
INV_X1 U860 ( .A(n972), .ZN(n1121) );
XOR2_X1 U861 ( .A(n1120), .B(KEYINPUT0), .Z(n1153) );
XOR2_X1 U862 ( .A(G110), .B(n1094), .Z(G12) );
AND3_X1 U863 ( .A1(n1097), .A2(n989), .A3(n1009), .ZN(n1094) );
NOR2_X1 U864 ( .A1(n1127), .A2(n1145), .ZN(n1009) );
XOR2_X1 U865 ( .A(n1154), .B(n1046), .Z(n1145) );
INV_X1 U866 ( .A(n968), .ZN(n1046) );
NAND2_X1 U867 ( .A1(G217), .A2(n1155), .ZN(n968) );
XNOR2_X1 U868 ( .A(KEYINPUT17), .B(n1156), .ZN(n1154) );
NOR3_X1 U869 ( .A1(n1157), .A2(KEYINPUT3), .A3(G902), .ZN(n1156) );
INV_X1 U870 ( .A(n970), .ZN(n1157) );
XOR2_X1 U871 ( .A(n1158), .B(n1159), .Z(n970) );
XOR2_X1 U872 ( .A(n1027), .B(n1160), .Z(n1159) );
XOR2_X1 U873 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U874 ( .A1(KEYINPUT40), .A2(n1163), .ZN(n1162) );
NAND2_X1 U875 ( .A1(G221), .A2(n1164), .ZN(n1161) );
XOR2_X1 U876 ( .A(n1125), .B(n1165), .Z(n1027) );
INV_X1 U877 ( .A(G137), .ZN(n1125) );
XNOR2_X1 U878 ( .A(G110), .B(n1166), .ZN(n1158) );
XOR2_X1 U879 ( .A(G146), .B(G128), .Z(n1166) );
XOR2_X1 U880 ( .A(n973), .B(KEYINPUT30), .Z(n1127) );
XOR2_X1 U881 ( .A(n1167), .B(G472), .Z(n973) );
NAND3_X1 U882 ( .A1(n1168), .A2(n1169), .A3(n971), .ZN(n1167) );
NAND2_X1 U883 ( .A1(KEYINPUT22), .A2(n1170), .ZN(n1169) );
XOR2_X1 U884 ( .A(n1171), .B(n1065), .Z(n1170) );
XNOR2_X1 U885 ( .A(n1172), .B(n1077), .ZN(n1065) );
XOR2_X1 U886 ( .A(G101), .B(n1173), .Z(n1077) );
NAND3_X1 U887 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1168) );
INV_X1 U888 ( .A(KEYINPUT22), .ZN(n1176) );
XOR2_X1 U889 ( .A(n1171), .B(n1173), .Z(n1175) );
INV_X1 U890 ( .A(n1177), .ZN(n1173) );
XOR2_X1 U891 ( .A(n1069), .B(n1064), .Z(n1171) );
XOR2_X1 U892 ( .A(n1083), .B(KEYINPUT23), .Z(n1064) );
NAND2_X1 U893 ( .A1(n1178), .A2(n1179), .ZN(n1069) );
NAND2_X1 U894 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U895 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U896 ( .A1(KEYINPUT6), .A2(n1184), .ZN(n1183) );
INV_X1 U897 ( .A(G113), .ZN(n1184) );
INV_X1 U898 ( .A(KEYINPUT52), .ZN(n1182) );
NAND2_X1 U899 ( .A1(G113), .A2(n1185), .ZN(n1178) );
NAND2_X1 U900 ( .A1(KEYINPUT6), .A2(n1186), .ZN(n1185) );
OR2_X1 U901 ( .A1(n1180), .A2(KEYINPUT52), .ZN(n1186) );
XOR2_X1 U902 ( .A(n1187), .B(G116), .Z(n1180) );
NAND2_X1 U903 ( .A1(KEYINPUT32), .A2(n1188), .ZN(n1187) );
XOR2_X1 U904 ( .A(n1133), .B(n1172), .Z(n1174) );
NAND2_X1 U905 ( .A1(G210), .A2(n1189), .ZN(n1172) );
NAND2_X1 U906 ( .A1(n1190), .A2(n1191), .ZN(n989) );
OR2_X1 U907 ( .A1(n999), .A2(KEYINPUT0), .ZN(n1191) );
NAND2_X1 U908 ( .A1(n972), .A2(n1120), .ZN(n999) );
NAND3_X1 U909 ( .A1(n1142), .A2(n972), .A3(KEYINPUT0), .ZN(n1190) );
XOR2_X1 U910 ( .A(n1192), .B(G475), .Z(n972) );
OR2_X1 U911 ( .A1(n1055), .A2(G902), .ZN(n1192) );
XNOR2_X1 U912 ( .A(n1193), .B(n1194), .ZN(n1055) );
XOR2_X1 U913 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U914 ( .A(n1197), .B(G104), .Z(n1196) );
NAND2_X1 U915 ( .A1(KEYINPUT48), .A2(n1198), .ZN(n1197) );
INV_X1 U916 ( .A(G131), .ZN(n1198) );
NAND2_X1 U917 ( .A1(G214), .A2(n1189), .ZN(n1195) );
NOR2_X1 U918 ( .A1(G953), .A2(G237), .ZN(n1189) );
XNOR2_X1 U919 ( .A(n1165), .B(n1199), .ZN(n1193) );
XOR2_X1 U920 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U921 ( .A(G140), .B(G125), .Z(n1165) );
INV_X1 U922 ( .A(n1120), .ZN(n1142) );
NAND2_X1 U923 ( .A1(n967), .A2(n976), .ZN(n1120) );
NAND3_X1 U924 ( .A1(n1052), .A2(n971), .A3(n1049), .ZN(n976) );
INV_X1 U925 ( .A(G478), .ZN(n1052) );
NAND2_X1 U926 ( .A1(G478), .A2(n1202), .ZN(n967) );
NAND2_X1 U927 ( .A1(n1049), .A2(n971), .ZN(n1202) );
XNOR2_X1 U928 ( .A(n1203), .B(n1204), .ZN(n1049) );
XOR2_X1 U929 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U930 ( .A(G128), .B(G122), .Z(n1206) );
XOR2_X1 U931 ( .A(G143), .B(G134), .Z(n1205) );
XOR2_X1 U932 ( .A(n1207), .B(n1208), .Z(n1203) );
XOR2_X1 U933 ( .A(G116), .B(G107), .Z(n1208) );
NAND2_X1 U934 ( .A1(G217), .A2(n1164), .ZN(n1207) );
AND2_X1 U935 ( .A1(G234), .A2(n958), .ZN(n1164) );
AND2_X1 U936 ( .A1(n1141), .A2(n1117), .ZN(n1097) );
INV_X1 U937 ( .A(n993), .ZN(n1117) );
NAND2_X1 U938 ( .A1(n1152), .A2(n960), .ZN(n993) );
NAND2_X1 U939 ( .A1(G221), .A2(n1155), .ZN(n960) );
NAND2_X1 U940 ( .A1(G234), .A2(n971), .ZN(n1155) );
INV_X1 U941 ( .A(n997), .ZN(n1152) );
XNOR2_X1 U942 ( .A(n963), .B(KEYINPUT18), .ZN(n997) );
XNOR2_X1 U943 ( .A(n1209), .B(G469), .ZN(n963) );
NAND2_X1 U944 ( .A1(n1210), .A2(n971), .ZN(n1209) );
XOR2_X1 U945 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U946 ( .A(n1177), .B(n1076), .Z(n1212) );
XOR2_X1 U947 ( .A(n1213), .B(n1214), .Z(n1076) );
XOR2_X1 U948 ( .A(G110), .B(n1215), .Z(n1214) );
AND2_X1 U949 ( .A1(n958), .A2(G227), .ZN(n1215) );
XNOR2_X1 U950 ( .A(G140), .B(KEYINPUT43), .ZN(n1213) );
XOR2_X1 U951 ( .A(n1216), .B(n1217), .Z(n1177) );
XOR2_X1 U952 ( .A(G137), .B(n1218), .Z(n1217) );
NOR2_X1 U953 ( .A1(G131), .A2(KEYINPUT60), .ZN(n1218) );
NAND2_X1 U954 ( .A1(KEYINPUT39), .A2(n1030), .ZN(n1216) );
INV_X1 U955 ( .A(G134), .ZN(n1030) );
XNOR2_X1 U956 ( .A(n1219), .B(KEYINPUT2), .ZN(n1211) );
NAND2_X1 U957 ( .A1(KEYINPUT51), .A2(n1220), .ZN(n1219) );
XOR2_X1 U958 ( .A(n1133), .B(n1078), .Z(n1220) );
XOR2_X1 U959 ( .A(n1221), .B(n1222), .Z(n1078) );
XNOR2_X1 U960 ( .A(KEYINPUT7), .B(n1029), .ZN(n1222) );
NAND2_X1 U961 ( .A1(n1223), .A2(n1224), .ZN(n1029) );
NAND2_X1 U962 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U963 ( .A(KEYINPUT54), .B(G128), .Z(n1226) );
XOR2_X1 U964 ( .A(n1227), .B(KEYINPUT1), .Z(n1223) );
NAND2_X1 U965 ( .A1(n1228), .A2(n1200), .ZN(n1227) );
XOR2_X1 U966 ( .A(n1132), .B(KEYINPUT27), .Z(n1228) );
NAND3_X1 U967 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1221) );
NAND2_X1 U968 ( .A1(n1059), .A2(n1232), .ZN(n1231) );
INV_X1 U969 ( .A(G104), .ZN(n1059) );
OR3_X1 U970 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1230) );
INV_X1 U971 ( .A(KEYINPUT34), .ZN(n1232) );
NAND2_X1 U972 ( .A1(n1234), .A2(n1233), .ZN(n1229) );
NAND2_X1 U973 ( .A1(KEYINPUT19), .A2(G104), .ZN(n1233) );
XOR2_X1 U974 ( .A(G107), .B(KEYINPUT55), .Z(n1234) );
INV_X1 U975 ( .A(G101), .ZN(n1133) );
AND2_X1 U976 ( .A1(n1115), .A2(n1235), .ZN(n1141) );
NAND2_X1 U977 ( .A1(n1015), .A2(n1236), .ZN(n1235) );
NAND3_X1 U978 ( .A1(n1035), .A2(n1139), .A3(G902), .ZN(n1236) );
NOR2_X1 U979 ( .A1(G898), .A2(n958), .ZN(n1035) );
NAND3_X1 U980 ( .A1(n1139), .A2(n958), .A3(G952), .ZN(n1015) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n1139) );
INV_X1 U982 ( .A(n1011), .ZN(n1115) );
NAND2_X1 U983 ( .A1(n1131), .A2(n975), .ZN(n1011) );
NAND2_X1 U984 ( .A1(G214), .A2(n977), .ZN(n975) );
NAND3_X1 U985 ( .A1(n1237), .A2(n1238), .A3(n974), .ZN(n1131) );
NAND2_X1 U986 ( .A1(n1239), .A2(n1240), .ZN(n974) );
NAND2_X1 U987 ( .A1(G210), .A2(n977), .ZN(n1240) );
NAND4_X1 U988 ( .A1(n977), .A2(n978), .A3(G210), .A4(n1241), .ZN(n1238) );
INV_X1 U989 ( .A(KEYINPUT61), .ZN(n1241) );
OR2_X1 U990 ( .A1(G902), .A2(G237), .ZN(n977) );
NAND2_X1 U991 ( .A1(KEYINPUT61), .A2(n1239), .ZN(n1237) );
INV_X1 U992 ( .A(n978), .ZN(n1239) );
NAND2_X1 U993 ( .A1(n1242), .A2(n971), .ZN(n978) );
INV_X1 U994 ( .A(G902), .ZN(n971) );
XOR2_X1 U995 ( .A(KEYINPUT44), .B(n1243), .Z(n1242) );
NOR2_X1 U996 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NOR2_X1 U997 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U998 ( .A(KEYINPUT11), .B(n1042), .Z(n1247) );
INV_X1 U999 ( .A(n1248), .ZN(n1246) );
NOR2_X1 U1000 ( .A1(n1042), .A2(n1248), .ZN(n1244) );
XOR2_X1 U1001 ( .A(n1086), .B(n1249), .Z(n1248) );
XOR2_X1 U1002 ( .A(G125), .B(n1250), .Z(n1249) );
NOR2_X1 U1003 ( .A1(KEYINPUT53), .A2(n1083), .ZN(n1250) );
XNOR2_X1 U1004 ( .A(n1132), .B(n1200), .ZN(n1083) );
INV_X1 U1005 ( .A(n1225), .ZN(n1200) );
XOR2_X1 U1006 ( .A(n1118), .B(G146), .Z(n1225) );
INV_X1 U1007 ( .A(G143), .ZN(n1118) );
INV_X1 U1008 ( .A(G128), .ZN(n1132) );
NAND2_X1 U1009 ( .A1(n1251), .A2(n958), .ZN(n1086) );
INV_X1 U1010 ( .A(G953), .ZN(n958) );
XOR2_X1 U1011 ( .A(KEYINPUT59), .B(G224), .Z(n1251) );
XNOR2_X1 U1012 ( .A(n1252), .B(n1253), .ZN(n1042) );
XOR2_X1 U1013 ( .A(n1163), .B(n1201), .Z(n1253) );
XOR2_X1 U1014 ( .A(G122), .B(G113), .Z(n1201) );
INV_X1 U1015 ( .A(n1188), .ZN(n1163) );
XNOR2_X1 U1016 ( .A(G119), .B(KEYINPUT31), .ZN(n1188) );
XOR2_X1 U1017 ( .A(n1254), .B(n1255), .Z(n1252) );
XNOR2_X1 U1018 ( .A(G110), .B(n1256), .ZN(n1255) );
NAND3_X1 U1019 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NAND2_X1 U1020 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
OR3_X1 U1021 ( .A1(n1261), .A2(n1260), .A3(n1262), .ZN(n1258) );
INV_X1 U1022 ( .A(KEYINPUT36), .ZN(n1261) );
NAND2_X1 U1023 ( .A1(n1262), .A2(n1263), .ZN(n1257) );
NAND2_X1 U1024 ( .A1(n1264), .A2(KEYINPUT36), .ZN(n1263) );
XNOR2_X1 U1025 ( .A(n1260), .B(KEYINPUT21), .ZN(n1264) );
XOR2_X1 U1026 ( .A(G104), .B(G107), .Z(n1260) );
XOR2_X1 U1027 ( .A(KEYINPUT7), .B(G101), .Z(n1262) );
NAND2_X1 U1028 ( .A1(KEYINPUT29), .A2(G116), .ZN(n1254) );
endmodule


