//Key = 0100011110000000010000010110100011110110111110010011000011100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354;

XNOR2_X1 U746 ( .A(G107), .B(n1038), .ZN(G9) );
NAND3_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR3_X1 U748 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
XNOR2_X1 U749 ( .A(n1045), .B(KEYINPUT7), .ZN(n1039) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U751 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
NOR3_X1 U753 ( .A1(n1054), .A2(KEYINPUT13), .A3(n1055), .ZN(n1048) );
INV_X1 U754 ( .A(n1056), .ZN(n1055) );
NOR2_X1 U755 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NOR3_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NOR4_X1 U757 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NOR2_X1 U758 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U759 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U760 ( .A1(KEYINPUT48), .A2(n1044), .ZN(n1068) );
NOR3_X1 U761 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1064) );
XNOR2_X1 U762 ( .A(n1073), .B(KEYINPUT39), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1043), .A2(n1074), .ZN(n1063) );
NOR2_X1 U764 ( .A1(n1075), .A2(n1076), .ZN(n1060) );
AND3_X1 U765 ( .A1(KEYINPUT48), .A2(n1077), .A3(n1078), .ZN(n1076) );
NOR3_X1 U766 ( .A1(n1067), .A2(n1079), .A3(n1074), .ZN(n1057) );
NOR3_X1 U767 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U769 ( .A(KEYINPUT50), .B(n1062), .ZN(n1084) );
INV_X1 U770 ( .A(n1085), .ZN(n1083) );
NOR2_X1 U771 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
INV_X1 U772 ( .A(n1088), .ZN(n1087) );
XNOR2_X1 U773 ( .A(n1075), .B(KEYINPUT2), .ZN(n1086) );
NOR2_X1 U774 ( .A1(n1089), .A2(n1059), .ZN(n1080) );
INV_X1 U775 ( .A(n1040), .ZN(n1059) );
NOR2_X1 U776 ( .A1(n1090), .A2(n1045), .ZN(n1089) );
NOR2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U778 ( .A(n1093), .B(KEYINPUT14), .ZN(n1091) );
AND3_X1 U779 ( .A1(n1052), .A2(n1053), .A3(n1094), .ZN(n1046) );
NAND4_X1 U780 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1052) );
NOR4_X1 U781 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1098) );
XOR2_X1 U782 ( .A(n1103), .B(n1104), .Z(n1099) );
XOR2_X1 U783 ( .A(KEYINPUT43), .B(G472), .Z(n1104) );
NOR2_X1 U784 ( .A1(n1105), .A2(n1106), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1107), .B(n1108), .Z(n1096) );
XOR2_X1 U786 ( .A(n1109), .B(KEYINPUT29), .Z(n1108) );
NAND2_X1 U787 ( .A1(KEYINPUT33), .A2(n1110), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1111), .B(n1112), .Z(n1095) );
NAND2_X1 U789 ( .A1(KEYINPUT57), .A2(n1113), .ZN(n1112) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(G72) );
NAND2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
OR2_X1 U792 ( .A1(n1053), .A2(G227), .ZN(n1117) );
NAND3_X1 U793 ( .A1(G953), .A2(n1118), .A3(n1119), .ZN(n1114) );
INV_X1 U794 ( .A(n1116), .ZN(n1119) );
XNOR2_X1 U795 ( .A(n1120), .B(n1121), .ZN(n1116) );
NOR4_X1 U796 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
NOR2_X1 U797 ( .A1(G140), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U798 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR3_X1 U799 ( .A1(G125), .A2(n1129), .A3(n1130), .ZN(n1123) );
AND3_X1 U800 ( .A1(G125), .A2(G140), .A3(n1129), .ZN(n1122) );
XOR2_X1 U801 ( .A(n1127), .B(n1131), .Z(n1129) );
NAND2_X1 U802 ( .A1(n1132), .A2(n1133), .ZN(n1127) );
NAND2_X1 U803 ( .A1(n1134), .A2(G137), .ZN(n1133) );
NAND2_X1 U804 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
XNOR2_X1 U805 ( .A(n1137), .B(KEYINPUT38), .ZN(n1135) );
NAND2_X1 U806 ( .A1(n1138), .A2(n1053), .ZN(n1120) );
XNOR2_X1 U807 ( .A(KEYINPUT37), .B(n1051), .ZN(n1138) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1118) );
NAND2_X1 U809 ( .A1(n1139), .A2(n1140), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
OR2_X1 U811 ( .A1(n1053), .A2(G224), .ZN(n1142) );
NAND3_X1 U812 ( .A1(G953), .A2(n1143), .A3(n1144), .ZN(n1139) );
INV_X1 U813 ( .A(n1141), .ZN(n1144) );
XNOR2_X1 U814 ( .A(n1145), .B(n1146), .ZN(n1141) );
NOR2_X1 U815 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U816 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U817 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U818 ( .A(n1153), .B(n1154), .Z(n1149) );
NOR2_X1 U819 ( .A1(G898), .A2(n1053), .ZN(n1147) );
NAND3_X1 U820 ( .A1(n1050), .A2(n1053), .A3(KEYINPUT26), .ZN(n1145) );
NAND2_X1 U821 ( .A1(G898), .A2(G224), .ZN(n1143) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XNOR2_X1 U823 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U824 ( .A(KEYINPUT19), .B(n1159), .Z(n1158) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U826 ( .A1(n1155), .A2(n1162), .ZN(G63) );
XNOR2_X1 U827 ( .A(n1163), .B(n1164), .ZN(n1162) );
AND2_X1 U828 ( .A1(G478), .A2(n1165), .ZN(n1164) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1166), .ZN(G60) );
XNOR2_X1 U830 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U831 ( .A1(n1113), .A2(n1161), .ZN(n1167) );
INV_X1 U832 ( .A(G475), .ZN(n1113) );
XOR2_X1 U833 ( .A(G104), .B(n1169), .Z(G6) );
NOR3_X1 U834 ( .A1(n1170), .A2(n1155), .A3(n1171), .ZN(G57) );
NOR3_X1 U835 ( .A1(n1172), .A2(KEYINPUT4), .A3(n1173), .ZN(n1171) );
XOR2_X1 U836 ( .A(n1174), .B(n1175), .Z(n1172) );
NOR2_X1 U837 ( .A1(n1176), .A2(KEYINPUT52), .ZN(n1174) );
NOR2_X1 U838 ( .A1(n1177), .A2(n1178), .ZN(n1170) );
XNOR2_X1 U839 ( .A(n1179), .B(n1175), .ZN(n1178) );
XNOR2_X1 U840 ( .A(n1180), .B(KEYINPUT56), .ZN(n1175) );
NAND2_X1 U841 ( .A1(n1176), .A2(n1181), .ZN(n1179) );
INV_X1 U842 ( .A(KEYINPUT52), .ZN(n1181) );
AND2_X1 U843 ( .A1(n1165), .A2(G472), .ZN(n1176) );
NOR2_X1 U844 ( .A1(KEYINPUT4), .A2(n1173), .ZN(n1177) );
XNOR2_X1 U845 ( .A(n1182), .B(n1183), .ZN(n1173) );
XNOR2_X1 U846 ( .A(n1131), .B(n1184), .ZN(n1183) );
XNOR2_X1 U847 ( .A(KEYINPUT11), .B(n1185), .ZN(n1182) );
NOR2_X1 U848 ( .A1(KEYINPUT24), .A2(n1186), .ZN(n1185) );
NOR2_X1 U849 ( .A1(n1155), .A2(n1187), .ZN(G54) );
XOR2_X1 U850 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U851 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR3_X1 U852 ( .A1(n1161), .A2(KEYINPUT46), .A3(n1110), .ZN(n1191) );
XNOR2_X1 U853 ( .A(n1192), .B(n1193), .ZN(n1188) );
NAND2_X1 U854 ( .A1(KEYINPUT17), .A2(n1194), .ZN(n1193) );
NAND2_X1 U855 ( .A1(KEYINPUT44), .A2(n1195), .ZN(n1192) );
XOR2_X1 U856 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U857 ( .A1(KEYINPUT59), .A2(n1198), .ZN(n1196) );
NOR2_X1 U858 ( .A1(n1155), .A2(n1199), .ZN(G51) );
XOR2_X1 U859 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR3_X1 U860 ( .A1(KEYINPUT21), .A2(n1202), .A3(n1203), .ZN(n1201) );
NOR2_X1 U861 ( .A1(n1204), .A2(n1128), .ZN(n1203) );
XOR2_X1 U862 ( .A(n1205), .B(n1206), .Z(n1204) );
XNOR2_X1 U863 ( .A(KEYINPUT34), .B(KEYINPUT23), .ZN(n1205) );
NOR2_X1 U864 ( .A1(n1207), .A2(n1206), .ZN(n1202) );
XNOR2_X1 U865 ( .A(n1208), .B(n1209), .ZN(n1206) );
NAND2_X1 U866 ( .A1(n1165), .A2(n1210), .ZN(n1200) );
INV_X1 U867 ( .A(n1161), .ZN(n1165) );
NAND2_X1 U868 ( .A1(G902), .A2(n1211), .ZN(n1161) );
OR2_X1 U869 ( .A1(n1051), .A2(n1050), .ZN(n1211) );
NAND4_X1 U870 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1050) );
AND4_X1 U871 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
NOR2_X1 U872 ( .A1(n1169), .A2(n1220), .ZN(n1214) );
AND3_X1 U873 ( .A1(n1221), .A2(n1077), .A3(n1040), .ZN(n1220) );
AND3_X1 U874 ( .A1(n1040), .A2(n1069), .A3(n1221), .ZN(n1169) );
NAND4_X1 U875 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1051) );
NOR4_X1 U876 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
INV_X1 U877 ( .A(n1230), .ZN(n1229) );
NOR2_X1 U878 ( .A1(n1231), .A2(n1232), .ZN(n1224) );
INV_X1 U879 ( .A(n1233), .ZN(n1232) );
NAND3_X1 U880 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1223) );
XNOR2_X1 U881 ( .A(n1045), .B(KEYINPUT8), .ZN(n1236) );
NAND3_X1 U882 ( .A1(n1045), .A2(n1069), .A3(n1237), .ZN(n1222) );
NOR2_X1 U883 ( .A1(n1053), .A2(G952), .ZN(n1155) );
XOR2_X1 U884 ( .A(n1238), .B(n1239), .Z(G48) );
NOR2_X1 U885 ( .A1(G146), .A2(KEYINPUT53), .ZN(n1239) );
NAND3_X1 U886 ( .A1(n1240), .A2(n1069), .A3(n1237), .ZN(n1238) );
XNOR2_X1 U887 ( .A(KEYINPUT0), .B(n1241), .ZN(n1240) );
XNOR2_X1 U888 ( .A(G143), .B(n1242), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1234), .A2(n1045), .A3(n1243), .A4(n1244), .ZN(n1242) );
OR2_X1 U890 ( .A1(n1235), .A2(KEYINPUT3), .ZN(n1244) );
NAND2_X1 U891 ( .A1(KEYINPUT3), .A2(n1245), .ZN(n1243) );
NAND2_X1 U892 ( .A1(n1246), .A2(n1043), .ZN(n1245) );
XOR2_X1 U893 ( .A(n1247), .B(n1248), .Z(G42) );
XNOR2_X1 U894 ( .A(KEYINPUT55), .B(n1130), .ZN(n1248) );
NOR2_X1 U895 ( .A1(KEYINPUT31), .A2(n1233), .ZN(n1247) );
NAND3_X1 U896 ( .A1(n1075), .A2(n1249), .A3(n1250), .ZN(n1233) );
XNOR2_X1 U897 ( .A(n1136), .B(n1231), .ZN(G39) );
AND3_X1 U898 ( .A1(n1073), .A2(n1237), .A3(n1075), .ZN(n1231) );
XOR2_X1 U899 ( .A(G134), .B(n1228), .Z(G36) );
NOR3_X1 U900 ( .A1(n1251), .A2(n1044), .A3(n1062), .ZN(n1228) );
INV_X1 U901 ( .A(n1077), .ZN(n1044) );
XOR2_X1 U902 ( .A(G131), .B(n1227), .Z(G33) );
AND3_X1 U903 ( .A1(n1235), .A2(n1069), .A3(n1075), .ZN(n1227) );
INV_X1 U904 ( .A(n1062), .ZN(n1075) );
NAND2_X1 U905 ( .A1(n1252), .A2(n1092), .ZN(n1062) );
XOR2_X1 U906 ( .A(KEYINPUT14), .B(n1093), .Z(n1252) );
INV_X1 U907 ( .A(n1251), .ZN(n1235) );
NAND2_X1 U908 ( .A1(n1246), .A2(n1249), .ZN(n1251) );
AND2_X1 U909 ( .A1(n1088), .A2(n1253), .ZN(n1246) );
XOR2_X1 U910 ( .A(G128), .B(n1226), .Z(G30) );
AND3_X1 U911 ( .A1(n1077), .A2(n1045), .A3(n1237), .ZN(n1226) );
AND4_X1 U912 ( .A1(n1254), .A2(n1253), .A3(n1249), .A4(n1100), .ZN(n1237) );
XNOR2_X1 U913 ( .A(G101), .B(n1216), .ZN(G3) );
NAND3_X1 U914 ( .A1(n1073), .A2(n1088), .A3(n1221), .ZN(n1216) );
XNOR2_X1 U915 ( .A(n1255), .B(n1256), .ZN(G27) );
NOR2_X1 U916 ( .A1(KEYINPUT22), .A2(n1230), .ZN(n1256) );
NAND3_X1 U917 ( .A1(n1250), .A2(n1045), .A3(n1078), .ZN(n1230) );
AND3_X1 U918 ( .A1(n1085), .A2(n1069), .A3(n1253), .ZN(n1250) );
AND2_X1 U919 ( .A1(n1257), .A2(n1056), .ZN(n1253) );
NAND2_X1 U920 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U921 ( .A1(n1124), .A2(G902), .ZN(n1259) );
NOR2_X1 U922 ( .A1(n1053), .A2(G900), .ZN(n1124) );
NAND2_X1 U923 ( .A1(G952), .A2(n1053), .ZN(n1258) );
XOR2_X1 U924 ( .A(n1212), .B(n1260), .Z(G24) );
XNOR2_X1 U925 ( .A(G122), .B(KEYINPUT63), .ZN(n1260) );
NAND3_X1 U926 ( .A1(n1234), .A2(n1040), .A3(n1261), .ZN(n1212) );
AND2_X1 U927 ( .A1(n1262), .A2(n1102), .ZN(n1234) );
XNOR2_X1 U928 ( .A(G119), .B(n1213), .ZN(G21) );
NAND4_X1 U929 ( .A1(n1261), .A2(n1073), .A3(n1254), .A4(n1100), .ZN(n1213) );
XNOR2_X1 U930 ( .A(G116), .B(n1219), .ZN(G18) );
NAND3_X1 U931 ( .A1(n1088), .A2(n1077), .A3(n1261), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1262), .A2(n1263), .ZN(n1077) );
XNOR2_X1 U933 ( .A(G113), .B(n1218), .ZN(G15) );
NAND3_X1 U934 ( .A1(n1088), .A2(n1069), .A3(n1261), .ZN(n1218) );
NOR3_X1 U935 ( .A1(n1042), .A2(n1241), .A3(n1067), .ZN(n1261) );
INV_X1 U936 ( .A(n1078), .ZN(n1067) );
NOR2_X1 U937 ( .A1(n1072), .A2(n1105), .ZN(n1078) );
NAND2_X1 U938 ( .A1(n1264), .A2(n1265), .ZN(n1069) );
OR2_X1 U939 ( .A1(n1074), .A2(KEYINPUT41), .ZN(n1265) );
INV_X1 U940 ( .A(n1073), .ZN(n1074) );
NAND3_X1 U941 ( .A1(n1262), .A2(n1263), .A3(KEYINPUT41), .ZN(n1264) );
INV_X1 U942 ( .A(n1102), .ZN(n1263) );
NOR2_X1 U943 ( .A1(n1266), .A2(n1100), .ZN(n1088) );
XNOR2_X1 U944 ( .A(G110), .B(n1217), .ZN(G12) );
NAND3_X1 U945 ( .A1(n1073), .A2(n1085), .A3(n1221), .ZN(n1217) );
NOR3_X1 U946 ( .A1(n1043), .A2(n1241), .A3(n1042), .ZN(n1221) );
NAND3_X1 U947 ( .A1(n1267), .A2(n1268), .A3(n1056), .ZN(n1042) );
NAND2_X1 U948 ( .A1(G237), .A2(G234), .ZN(n1056) );
NAND2_X1 U949 ( .A1(n1094), .A2(n1053), .ZN(n1268) );
INV_X1 U950 ( .A(G952), .ZN(n1094) );
NAND2_X1 U951 ( .A1(G953), .A2(n1269), .ZN(n1267) );
OR2_X1 U952 ( .A1(n1270), .A2(G898), .ZN(n1269) );
INV_X1 U953 ( .A(n1045), .ZN(n1241) );
NOR2_X1 U954 ( .A1(n1093), .A2(n1106), .ZN(n1045) );
INV_X1 U955 ( .A(n1092), .ZN(n1106) );
NAND2_X1 U956 ( .A1(G214), .A2(n1271), .ZN(n1092) );
XOR2_X1 U957 ( .A(n1101), .B(n1272), .Z(n1093) );
XOR2_X1 U958 ( .A(KEYINPUT49), .B(KEYINPUT1), .Z(n1272) );
XNOR2_X1 U959 ( .A(n1273), .B(n1210), .ZN(n1101) );
AND2_X1 U960 ( .A1(G210), .A2(n1271), .ZN(n1210) );
NAND2_X1 U961 ( .A1(n1274), .A2(n1270), .ZN(n1271) );
INV_X1 U962 ( .A(G237), .ZN(n1274) );
NAND2_X1 U963 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
XOR2_X1 U964 ( .A(n1277), .B(n1209), .Z(n1276) );
XNOR2_X1 U965 ( .A(n1278), .B(n1279), .ZN(n1209) );
XOR2_X1 U966 ( .A(G122), .B(n1154), .Z(n1279) );
NOR2_X1 U967 ( .A1(KEYINPUT15), .A2(G110), .ZN(n1154) );
NAND2_X1 U968 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
NAND2_X1 U969 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U970 ( .A(n1153), .B(n1284), .Z(n1282) );
OR3_X1 U971 ( .A1(n1153), .A2(n1284), .A3(n1283), .ZN(n1280) );
INV_X1 U972 ( .A(KEYINPUT12), .ZN(n1283) );
XOR2_X1 U973 ( .A(G113), .B(n1152), .Z(n1284) );
XOR2_X1 U974 ( .A(G116), .B(n1285), .Z(n1152) );
NOR2_X1 U975 ( .A1(G119), .A2(KEYINPUT10), .ZN(n1285) );
XOR2_X1 U976 ( .A(n1286), .B(n1287), .Z(n1153) );
XNOR2_X1 U977 ( .A(n1288), .B(n1289), .ZN(n1286) );
NAND2_X1 U978 ( .A1(KEYINPUT51), .A2(n1290), .ZN(n1288) );
NAND2_X1 U979 ( .A1(n1291), .A2(KEYINPUT47), .ZN(n1277) );
XNOR2_X1 U980 ( .A(n1292), .B(n1128), .ZN(n1291) );
INV_X1 U981 ( .A(n1207), .ZN(n1128) );
XNOR2_X1 U982 ( .A(G125), .B(n1131), .ZN(n1207) );
XOR2_X1 U983 ( .A(n1208), .B(KEYINPUT45), .Z(n1292) );
NAND2_X1 U984 ( .A1(G224), .A2(n1053), .ZN(n1208) );
INV_X1 U985 ( .A(n1249), .ZN(n1043) );
NOR2_X1 U986 ( .A1(n1293), .A2(n1105), .ZN(n1249) );
INV_X1 U987 ( .A(n1070), .ZN(n1105) );
NAND2_X1 U988 ( .A1(G221), .A2(n1294), .ZN(n1070) );
INV_X1 U989 ( .A(n1072), .ZN(n1293) );
XNOR2_X1 U990 ( .A(n1109), .B(n1295), .ZN(n1072) );
XNOR2_X1 U991 ( .A(KEYINPUT27), .B(n1110), .ZN(n1295) );
INV_X1 U992 ( .A(G469), .ZN(n1110) );
NAND2_X1 U993 ( .A1(n1296), .A2(n1275), .ZN(n1109) );
XOR2_X1 U994 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U995 ( .A(n1194), .B(n1299), .ZN(n1298) );
XOR2_X1 U996 ( .A(KEYINPUT62), .B(KEYINPUT18), .Z(n1299) );
NAND2_X1 U997 ( .A1(G227), .A2(n1053), .ZN(n1194) );
XOR2_X1 U998 ( .A(n1190), .B(n1300), .Z(n1297) );
XNOR2_X1 U999 ( .A(n1301), .B(n1197), .ZN(n1300) );
XNOR2_X1 U1000 ( .A(n1302), .B(n1287), .ZN(n1197) );
XNOR2_X1 U1001 ( .A(n1303), .B(n1290), .ZN(n1302) );
NAND2_X1 U1002 ( .A1(KEYINPUT5), .A2(n1289), .ZN(n1303) );
NAND2_X1 U1003 ( .A1(KEYINPUT58), .A2(n1131), .ZN(n1301) );
XNOR2_X1 U1004 ( .A(n1186), .B(n1304), .ZN(n1190) );
XNOR2_X1 U1005 ( .A(n1130), .B(G110), .ZN(n1304) );
NAND2_X1 U1006 ( .A1(n1305), .A2(n1306), .ZN(n1085) );
NAND3_X1 U1007 ( .A1(n1266), .A2(n1100), .A3(n1307), .ZN(n1306) );
INV_X1 U1008 ( .A(KEYINPUT9), .ZN(n1307) );
NAND2_X1 U1009 ( .A1(KEYINPUT9), .A2(n1040), .ZN(n1305) );
NOR2_X1 U1010 ( .A1(n1100), .A2(n1254), .ZN(n1040) );
INV_X1 U1011 ( .A(n1266), .ZN(n1254) );
XNOR2_X1 U1012 ( .A(n1308), .B(G472), .ZN(n1266) );
NAND2_X1 U1013 ( .A1(KEYINPUT61), .A2(n1103), .ZN(n1308) );
NAND2_X1 U1014 ( .A1(n1275), .A2(n1309), .ZN(n1103) );
XOR2_X1 U1015 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1016 ( .A(n1180), .B(n1131), .ZN(n1311) );
INV_X1 U1017 ( .A(n1198), .ZN(n1131) );
XOR2_X1 U1018 ( .A(G143), .B(n1312), .Z(n1198) );
XNOR2_X1 U1019 ( .A(n1313), .B(n1289), .ZN(n1180) );
INV_X1 U1020 ( .A(G101), .ZN(n1289) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1022 ( .A(n1315), .B(n1316), .ZN(n1310) );
NAND2_X1 U1023 ( .A1(KEYINPUT42), .A2(n1317), .ZN(n1316) );
INV_X1 U1024 ( .A(n1186), .ZN(n1317) );
XNOR2_X1 U1025 ( .A(G137), .B(n1134), .ZN(n1186) );
INV_X1 U1026 ( .A(n1137), .ZN(n1134) );
XNOR2_X1 U1027 ( .A(n1318), .B(n1319), .ZN(n1137) );
XNOR2_X1 U1028 ( .A(G131), .B(KEYINPUT40), .ZN(n1318) );
NAND2_X1 U1029 ( .A1(KEYINPUT32), .A2(n1184), .ZN(n1315) );
XNOR2_X1 U1030 ( .A(n1320), .B(n1321), .ZN(n1184) );
XNOR2_X1 U1031 ( .A(n1322), .B(G116), .ZN(n1321) );
INV_X1 U1032 ( .A(G119), .ZN(n1322) );
INV_X1 U1033 ( .A(G113), .ZN(n1320) );
XOR2_X1 U1034 ( .A(n1323), .B(n1160), .Z(n1100) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1294), .ZN(n1160) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1270), .ZN(n1294) );
INV_X1 U1037 ( .A(G902), .ZN(n1270) );
NAND2_X1 U1038 ( .A1(n1275), .A2(n1157), .ZN(n1323) );
XOR2_X1 U1039 ( .A(n1324), .B(n1325), .Z(n1157) );
XNOR2_X1 U1040 ( .A(n1312), .B(n1326), .ZN(n1325) );
XOR2_X1 U1041 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1042 ( .A1(KEYINPUT54), .A2(n1136), .ZN(n1328) );
INV_X1 U1043 ( .A(G137), .ZN(n1136) );
NAND2_X1 U1044 ( .A1(n1329), .A2(n1330), .ZN(n1327) );
NAND2_X1 U1045 ( .A1(G125), .A2(n1130), .ZN(n1330) );
INV_X1 U1046 ( .A(G140), .ZN(n1130) );
XOR2_X1 U1047 ( .A(n1331), .B(KEYINPUT20), .Z(n1329) );
NAND2_X1 U1048 ( .A1(n1332), .A2(n1255), .ZN(n1331) );
INV_X1 U1049 ( .A(G125), .ZN(n1255) );
XNOR2_X1 U1050 ( .A(G140), .B(KEYINPUT25), .ZN(n1332) );
XOR2_X1 U1051 ( .A(G128), .B(G146), .Z(n1312) );
XOR2_X1 U1052 ( .A(n1333), .B(n1334), .Z(n1324) );
AND3_X1 U1053 ( .A1(G221), .A2(n1053), .A3(G234), .ZN(n1334) );
XNOR2_X1 U1054 ( .A(G110), .B(G119), .ZN(n1333) );
NOR2_X1 U1055 ( .A1(n1102), .A2(n1262), .ZN(n1073) );
XOR2_X1 U1056 ( .A(n1335), .B(n1111), .Z(n1262) );
NAND2_X1 U1057 ( .A1(n1168), .A2(n1275), .ZN(n1111) );
XOR2_X1 U1058 ( .A(n1336), .B(n1337), .Z(n1168) );
XOR2_X1 U1059 ( .A(n1151), .B(n1338), .Z(n1337) );
XOR2_X1 U1060 ( .A(n1339), .B(n1287), .Z(n1338) );
XOR2_X1 U1061 ( .A(G104), .B(KEYINPUT6), .Z(n1287) );
NAND2_X1 U1062 ( .A1(n1340), .A2(KEYINPUT35), .ZN(n1339) );
XOR2_X1 U1063 ( .A(n1341), .B(n1342), .Z(n1340) );
XNOR2_X1 U1064 ( .A(n1343), .B(G131), .ZN(n1342) );
INV_X1 U1065 ( .A(G143), .ZN(n1343) );
NAND2_X1 U1066 ( .A1(G214), .A2(n1314), .ZN(n1341) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1314) );
XNOR2_X1 U1068 ( .A(G113), .B(G122), .ZN(n1151) );
XOR2_X1 U1069 ( .A(n1344), .B(n1345), .Z(n1336) );
NOR2_X1 U1070 ( .A1(G140), .A2(KEYINPUT30), .ZN(n1345) );
XNOR2_X1 U1071 ( .A(G146), .B(G125), .ZN(n1344) );
NAND2_X1 U1072 ( .A1(KEYINPUT28), .A2(G475), .ZN(n1335) );
XNOR2_X1 U1073 ( .A(n1346), .B(G478), .ZN(n1102) );
NAND2_X1 U1074 ( .A1(n1275), .A2(n1347), .ZN(n1346) );
XNOR2_X1 U1075 ( .A(KEYINPUT60), .B(n1348), .ZN(n1347) );
INV_X1 U1076 ( .A(n1163), .ZN(n1348) );
XNOR2_X1 U1077 ( .A(n1349), .B(n1350), .ZN(n1163) );
XOR2_X1 U1078 ( .A(n1319), .B(n1351), .Z(n1350) );
XNOR2_X1 U1079 ( .A(n1290), .B(n1352), .ZN(n1351) );
AND3_X1 U1080 ( .A1(G217), .A2(n1053), .A3(G234), .ZN(n1352) );
INV_X1 U1081 ( .A(G953), .ZN(n1053) );
INV_X1 U1082 ( .A(G107), .ZN(n1290) );
XOR2_X1 U1083 ( .A(G134), .B(KEYINPUT36), .Z(n1319) );
XOR2_X1 U1084 ( .A(n1353), .B(n1354), .Z(n1349) );
XOR2_X1 U1085 ( .A(G122), .B(G116), .Z(n1354) );
XNOR2_X1 U1086 ( .A(G128), .B(G143), .ZN(n1353) );
XNOR2_X1 U1087 ( .A(G902), .B(KEYINPUT16), .ZN(n1275) );
endmodule


