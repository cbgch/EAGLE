//Key = 0011010101000100001011010110000010100001001001100000001010010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391;

XNOR2_X1 U762 ( .A(G107), .B(n1059), .ZN(G9) );
NAND3_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
AND3_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
XNOR2_X1 U765 ( .A(n1066), .B(KEYINPUT39), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(G75) );
AND4_X1 U767 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(G952), .ZN(n1068) );
AND3_X1 U768 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1069) );
NAND3_X1 U769 ( .A1(n1063), .A2(n1075), .A3(n1076), .ZN(n1074) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND3_X1 U771 ( .A1(n1061), .A2(n1079), .A3(n1080), .ZN(n1078) );
XOR2_X1 U772 ( .A(KEYINPUT48), .B(n1081), .Z(n1079) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1077) );
NAND3_X1 U774 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1066), .A2(n1086), .ZN(n1085) );
XOR2_X1 U776 ( .A(KEYINPUT6), .B(n1087), .Z(n1086) );
NAND3_X1 U777 ( .A1(n1088), .A2(n1080), .A3(n1089), .ZN(n1084) );
NAND3_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1087), .ZN(n1083) );
NAND4_X1 U779 ( .A1(n1081), .A2(n1087), .A3(n1080), .A4(n1092), .ZN(n1072) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1063), .A2(n1095), .ZN(n1094) );
OR2_X1 U782 ( .A1(n1096), .A2(n1065), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1076), .A2(n1097), .ZN(n1093) );
NAND2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U786 ( .A(n1102), .ZN(n1098) );
INV_X1 U787 ( .A(n1103), .ZN(n1081) );
AND3_X1 U788 ( .A1(n1104), .A2(n1073), .A3(n1071), .ZN(n1067) );
NAND4_X1 U789 ( .A1(n1087), .A2(n1080), .A3(n1105), .A4(n1106), .ZN(n1073) );
NOR3_X1 U790 ( .A1(n1101), .A2(n1107), .A3(n1108), .ZN(n1106) );
XOR2_X1 U791 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U792 ( .A1(KEYINPUT25), .A2(n1111), .ZN(n1109) );
INV_X1 U793 ( .A(G472), .ZN(n1111) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1107) );
NAND2_X1 U795 ( .A1(KEYINPUT7), .A2(n1114), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1105) );
XNOR2_X1 U797 ( .A(KEYINPUT52), .B(G952), .ZN(n1104) );
NAND2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(G72) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U800 ( .A(n1121), .B(n1122), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1123), .A2(KEYINPUT19), .ZN(n1122) );
INV_X1 U802 ( .A(n1124), .ZN(n1123) );
NAND2_X1 U803 ( .A1(n1125), .A2(G953), .ZN(n1117) );
XOR2_X1 U804 ( .A(n1121), .B(n1126), .Z(n1125) );
AND2_X1 U805 ( .A1(G227), .A2(G900), .ZN(n1126) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
NAND2_X1 U807 ( .A1(G953), .A2(n1129), .ZN(n1128) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1127) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(n1130) );
NOR2_X1 U811 ( .A1(KEYINPUT4), .A2(G131), .ZN(n1135) );
XOR2_X1 U812 ( .A(n1136), .B(G137), .Z(n1134) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(G69) );
NAND2_X1 U814 ( .A1(G953), .A2(n1139), .ZN(n1138) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1139) );
NAND2_X1 U816 ( .A1(n1140), .A2(KEYINPUT18), .ZN(n1137) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U818 ( .A1(G953), .A2(n1143), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U820 ( .A(KEYINPUT33), .B(n1146), .Z(n1145) );
NAND2_X1 U821 ( .A1(KEYINPUT46), .A2(n1147), .ZN(n1141) );
NAND3_X1 U822 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NAND2_X1 U823 ( .A1(G953), .A2(n1151), .ZN(n1150) );
NAND2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NAND2_X1 U825 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U826 ( .A1(KEYINPUT41), .A2(n1156), .ZN(n1155) );
NAND3_X1 U827 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1148) );
INV_X1 U828 ( .A(KEYINPUT41), .ZN(n1159) );
NAND2_X1 U829 ( .A1(n1160), .A2(n1156), .ZN(n1158) );
INV_X1 U830 ( .A(KEYINPUT30), .ZN(n1156) );
NAND2_X1 U831 ( .A1(n1154), .A2(n1161), .ZN(n1157) );
OR2_X1 U832 ( .A1(n1152), .A2(KEYINPUT30), .ZN(n1161) );
XNOR2_X1 U833 ( .A(n1162), .B(n1163), .ZN(n1152) );
NOR2_X1 U834 ( .A1(n1164), .A2(KEYINPUT12), .ZN(n1163) );
INV_X1 U835 ( .A(n1165), .ZN(n1164) );
NOR2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(G66) );
XNOR2_X1 U837 ( .A(n1168), .B(n1169), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U839 ( .A1(n1166), .A2(n1172), .ZN(G63) );
XOR2_X1 U840 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U841 ( .A1(KEYINPUT21), .A2(n1175), .ZN(n1173) );
NAND2_X1 U842 ( .A1(n1176), .A2(G478), .ZN(n1175) );
NOR2_X1 U843 ( .A1(n1166), .A2(n1177), .ZN(G60) );
NOR3_X1 U844 ( .A1(n1115), .A2(n1178), .A3(n1179), .ZN(n1177) );
AND3_X1 U845 ( .A1(n1180), .A2(G475), .A3(n1176), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1181), .A2(n1180), .ZN(n1178) );
NOR2_X1 U847 ( .A1(n1070), .A2(n1116), .ZN(n1181) );
INV_X1 U848 ( .A(G475), .ZN(n1116) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(G6) );
NOR2_X1 U850 ( .A1(n1166), .A2(n1184), .ZN(G57) );
XOR2_X1 U851 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U853 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U855 ( .A1(n1193), .A2(n1194), .ZN(n1189) );
XNOR2_X1 U856 ( .A(n1191), .B(KEYINPUT1), .ZN(n1193) );
XNOR2_X1 U857 ( .A(n1195), .B(n1196), .ZN(n1191) );
XNOR2_X1 U858 ( .A(n1197), .B(KEYINPUT56), .ZN(n1185) );
NAND2_X1 U859 ( .A1(KEYINPUT26), .A2(n1198), .ZN(n1197) );
NAND2_X1 U860 ( .A1(n1176), .A2(G472), .ZN(n1198) );
NOR2_X1 U861 ( .A1(n1166), .A2(n1199), .ZN(G54) );
XOR2_X1 U862 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U863 ( .A(n1202), .B(n1203), .ZN(n1201) );
NAND2_X1 U864 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
NAND3_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1204) );
NAND2_X1 U867 ( .A1(n1206), .A2(n1207), .ZN(n1210) );
INV_X1 U868 ( .A(n1211), .ZN(n1207) );
XNOR2_X1 U869 ( .A(KEYINPUT23), .B(n1212), .ZN(n1206) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U871 ( .A(KEYINPUT24), .B(G110), .Z(n1214) );
XOR2_X1 U872 ( .A(n1215), .B(KEYINPUT37), .Z(n1213) );
XNOR2_X1 U873 ( .A(n1208), .B(KEYINPUT63), .ZN(n1209) );
XOR2_X1 U874 ( .A(KEYINPUT20), .B(n1216), .Z(n1200) );
AND2_X1 U875 ( .A1(G469), .A2(n1176), .ZN(n1216) );
NOR2_X1 U876 ( .A1(n1166), .A2(n1217), .ZN(G51) );
XOR2_X1 U877 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U878 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR2_X1 U879 ( .A1(n1222), .A2(n1171), .ZN(n1221) );
INV_X1 U880 ( .A(n1176), .ZN(n1171) );
NOR2_X1 U881 ( .A1(n1223), .A2(n1070), .ZN(n1176) );
NOR3_X1 U882 ( .A1(n1144), .A2(n1146), .A3(n1124), .ZN(n1070) );
NAND4_X1 U883 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1124) );
NOR4_X1 U884 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
NOR3_X1 U885 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1226) );
NOR3_X1 U886 ( .A1(n1235), .A2(n1061), .A3(n1236), .ZN(n1234) );
INV_X1 U887 ( .A(KEYINPUT31), .ZN(n1235) );
NOR2_X1 U888 ( .A1(KEYINPUT31), .A2(n1237), .ZN(n1233) );
NOR2_X1 U889 ( .A1(n1238), .A2(n1239), .ZN(n1232) );
INV_X1 U890 ( .A(n1080), .ZN(n1239) );
XNOR2_X1 U891 ( .A(n1240), .B(KEYINPUT55), .ZN(n1238) );
INV_X1 U892 ( .A(n1241), .ZN(n1146) );
NAND4_X1 U893 ( .A1(n1183), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1144) );
AND4_X1 U894 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1244) );
NAND4_X1 U895 ( .A1(n1249), .A2(n1064), .A3(n1066), .A4(n1250), .ZN(n1243) );
AND2_X1 U896 ( .A1(n1065), .A2(n1063), .ZN(n1250) );
XOR2_X1 U897 ( .A(KEYINPUT58), .B(n1061), .Z(n1249) );
NAND3_X1 U898 ( .A1(n1251), .A2(n1063), .A3(n1096), .ZN(n1183) );
NAND3_X1 U899 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1220) );
OR2_X1 U900 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND2_X1 U901 ( .A1(KEYINPUT11), .A2(n1257), .ZN(n1253) );
NAND3_X1 U902 ( .A1(n1258), .A2(n1259), .A3(n1255), .ZN(n1257) );
NAND2_X1 U903 ( .A1(G125), .A2(n1260), .ZN(n1259) );
NAND3_X1 U904 ( .A1(n1192), .A2(n1256), .A3(n1261), .ZN(n1258) );
NAND2_X1 U905 ( .A1(n1262), .A2(n1263), .ZN(n1252) );
INV_X1 U906 ( .A(KEYINPUT11), .ZN(n1263) );
NOR2_X1 U907 ( .A1(n1120), .A2(G952), .ZN(n1166) );
XOR2_X1 U908 ( .A(G146), .B(n1231), .Z(G48) );
AND3_X1 U909 ( .A1(n1096), .A2(n1066), .A3(n1264), .ZN(n1231) );
XOR2_X1 U910 ( .A(n1237), .B(n1265), .Z(G45) );
NOR2_X1 U911 ( .A1(G143), .A2(KEYINPUT60), .ZN(n1265) );
NAND2_X1 U912 ( .A1(n1266), .A2(n1061), .ZN(n1237) );
INV_X1 U913 ( .A(n1236), .ZN(n1266) );
NAND3_X1 U914 ( .A1(n1267), .A2(n1102), .A3(n1268), .ZN(n1236) );
AND3_X1 U915 ( .A1(n1066), .A2(n1269), .A3(n1270), .ZN(n1268) );
XOR2_X1 U916 ( .A(n1215), .B(n1271), .Z(G42) );
NAND2_X1 U917 ( .A1(n1240), .A2(n1080), .ZN(n1271) );
AND2_X1 U918 ( .A1(n1272), .A2(n1061), .ZN(n1240) );
XOR2_X1 U919 ( .A(G137), .B(n1230), .Z(G39) );
AND3_X1 U920 ( .A1(n1076), .A2(n1080), .A3(n1264), .ZN(n1230) );
XOR2_X1 U921 ( .A(n1273), .B(n1229), .Z(G36) );
AND2_X1 U922 ( .A1(n1274), .A2(n1065), .ZN(n1229) );
XOR2_X1 U923 ( .A(n1136), .B(KEYINPUT59), .Z(n1273) );
XOR2_X1 U924 ( .A(G131), .B(n1228), .Z(G33) );
AND2_X1 U925 ( .A1(n1096), .A2(n1274), .ZN(n1228) );
AND4_X1 U926 ( .A1(n1102), .A2(n1080), .A3(n1061), .A4(n1269), .ZN(n1274) );
NOR2_X1 U927 ( .A1(n1275), .A2(n1091), .ZN(n1080) );
NAND3_X1 U928 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(G30) );
NAND2_X1 U929 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U930 ( .A1(KEYINPUT16), .A2(n1281), .ZN(n1277) );
NAND2_X1 U931 ( .A1(n1282), .A2(n1224), .ZN(n1281) );
XOR2_X1 U932 ( .A(KEYINPUT17), .B(G128), .Z(n1282) );
NAND2_X1 U933 ( .A1(n1283), .A2(n1284), .ZN(n1276) );
INV_X1 U934 ( .A(KEYINPUT16), .ZN(n1284) );
NAND2_X1 U935 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U936 ( .A1(KEYINPUT17), .A2(n1280), .ZN(n1286) );
OR3_X1 U937 ( .A1(n1279), .A2(KEYINPUT17), .A3(n1280), .ZN(n1285) );
INV_X1 U938 ( .A(n1224), .ZN(n1279) );
NAND3_X1 U939 ( .A1(n1065), .A2(n1066), .A3(n1264), .ZN(n1224) );
AND4_X1 U940 ( .A1(n1061), .A2(n1101), .A3(n1287), .A4(n1269), .ZN(n1264) );
XNOR2_X1 U941 ( .A(n1242), .B(n1288), .ZN(G3) );
NOR2_X1 U942 ( .A1(KEYINPUT35), .A2(n1289), .ZN(n1288) );
NAND3_X1 U943 ( .A1(n1076), .A2(n1251), .A3(n1102), .ZN(n1242) );
XOR2_X1 U944 ( .A(n1256), .B(n1225), .Z(G27) );
NAND3_X1 U945 ( .A1(n1087), .A2(n1066), .A3(n1272), .ZN(n1225) );
AND4_X1 U946 ( .A1(n1100), .A2(n1096), .A3(n1101), .A4(n1269), .ZN(n1272) );
NAND2_X1 U947 ( .A1(n1103), .A2(n1290), .ZN(n1269) );
NAND4_X1 U948 ( .A1(G902), .A2(G953), .A3(n1291), .A4(n1129), .ZN(n1290) );
INV_X1 U949 ( .A(G900), .ZN(n1129) );
XNOR2_X1 U950 ( .A(G122), .B(n1248), .ZN(G24) );
NAND4_X1 U951 ( .A1(n1267), .A2(n1292), .A3(n1063), .A4(n1270), .ZN(n1248) );
NOR2_X1 U952 ( .A1(n1287), .A2(n1101), .ZN(n1063) );
XOR2_X1 U953 ( .A(n1293), .B(n1247), .Z(G21) );
NAND4_X1 U954 ( .A1(n1292), .A2(n1076), .A3(n1101), .A4(n1287), .ZN(n1247) );
INV_X1 U955 ( .A(n1100), .ZN(n1287) );
XOR2_X1 U956 ( .A(n1294), .B(n1246), .Z(G18) );
NAND3_X1 U957 ( .A1(n1102), .A2(n1065), .A3(n1292), .ZN(n1246) );
NOR2_X1 U958 ( .A1(n1295), .A2(n1267), .ZN(n1065) );
XOR2_X1 U959 ( .A(n1296), .B(n1245), .Z(G15) );
NAND3_X1 U960 ( .A1(n1096), .A2(n1102), .A3(n1292), .ZN(n1245) );
AND3_X1 U961 ( .A1(n1066), .A2(n1064), .A3(n1087), .ZN(n1292) );
NOR2_X1 U962 ( .A1(n1297), .A2(n1089), .ZN(n1087) );
INV_X1 U963 ( .A(n1088), .ZN(n1297) );
NOR2_X1 U964 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
AND2_X1 U965 ( .A1(n1267), .A2(n1298), .ZN(n1096) );
XOR2_X1 U966 ( .A(KEYINPUT2), .B(n1270), .Z(n1298) );
XOR2_X1 U967 ( .A(n1241), .B(n1299), .Z(G12) );
NOR2_X1 U968 ( .A1(G110), .A2(KEYINPUT10), .ZN(n1299) );
NAND4_X1 U969 ( .A1(n1076), .A2(n1251), .A3(n1100), .A4(n1101), .ZN(n1241) );
XOR2_X1 U970 ( .A(n1300), .B(n1170), .Z(n1101) );
NAND2_X1 U971 ( .A1(G217), .A2(n1301), .ZN(n1170) );
NAND2_X1 U972 ( .A1(n1168), .A2(n1223), .ZN(n1300) );
XNOR2_X1 U973 ( .A(n1302), .B(n1303), .ZN(n1168) );
XOR2_X1 U974 ( .A(G119), .B(n1304), .Z(n1303) );
XOR2_X1 U975 ( .A(G137), .B(G128), .Z(n1304) );
XOR2_X1 U976 ( .A(n1305), .B(n1306), .Z(n1302) );
AND2_X1 U977 ( .A1(G221), .A2(n1307), .ZN(n1306) );
XOR2_X1 U978 ( .A(n1308), .B(G110), .Z(n1305) );
NAND2_X1 U979 ( .A1(n1309), .A2(KEYINPUT45), .ZN(n1308) );
XNOR2_X1 U980 ( .A(n1133), .B(n1310), .ZN(n1309) );
NOR2_X1 U981 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1310) );
XOR2_X1 U982 ( .A(n1311), .B(G472), .Z(n1100) );
NAND2_X1 U983 ( .A1(KEYINPUT54), .A2(n1110), .ZN(n1311) );
AND2_X1 U984 ( .A1(n1312), .A2(n1223), .ZN(n1110) );
XOR2_X1 U985 ( .A(n1313), .B(n1314), .Z(n1312) );
XOR2_X1 U986 ( .A(n1187), .B(n1196), .Z(n1314) );
XOR2_X1 U987 ( .A(n1315), .B(G101), .Z(n1187) );
NAND2_X1 U988 ( .A1(G210), .A2(n1316), .ZN(n1315) );
XOR2_X1 U989 ( .A(n1195), .B(n1317), .Z(n1313) );
XOR2_X1 U990 ( .A(KEYINPUT61), .B(n1192), .Z(n1317) );
XOR2_X1 U991 ( .A(n1318), .B(n1319), .Z(n1195) );
NOR2_X1 U992 ( .A1(KEYINPUT0), .A2(n1320), .ZN(n1319) );
XOR2_X1 U993 ( .A(KEYINPUT29), .B(G116), .Z(n1320) );
XOR2_X1 U994 ( .A(n1293), .B(G113), .Z(n1318) );
AND3_X1 U995 ( .A1(n1066), .A2(n1064), .A3(n1061), .ZN(n1251) );
NOR2_X1 U996 ( .A1(n1088), .A2(n1089), .ZN(n1061) );
AND2_X1 U997 ( .A1(G221), .A2(n1301), .ZN(n1089) );
NAND2_X1 U998 ( .A1(G234), .A2(n1223), .ZN(n1301) );
XOR2_X1 U999 ( .A(n1321), .B(G469), .Z(n1088) );
NAND4_X1 U1000 ( .A1(n1322), .A2(n1223), .A3(n1323), .A4(n1324), .ZN(n1321) );
NAND3_X1 U1001 ( .A1(G110), .A2(n1325), .A3(G140), .ZN(n1324) );
NAND2_X1 U1002 ( .A1(n1326), .A2(n1215), .ZN(n1323) );
XOR2_X1 U1003 ( .A(G110), .B(n1325), .Z(n1326) );
NAND2_X1 U1004 ( .A1(n1211), .A2(n1327), .ZN(n1322) );
INV_X1 U1005 ( .A(n1325), .ZN(n1327) );
XNOR2_X1 U1006 ( .A(n1208), .B(n1328), .ZN(n1325) );
NOR2_X1 U1007 ( .A1(KEYINPUT57), .A2(n1203), .ZN(n1328) );
XNOR2_X1 U1008 ( .A(n1329), .B(n1330), .ZN(n1203) );
NOR2_X1 U1009 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NOR2_X1 U1010 ( .A1(n1289), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1011 ( .A(n1334), .B(KEYINPUT42), .Z(n1333) );
NOR2_X1 U1012 ( .A1(G101), .A2(n1335), .ZN(n1331) );
XOR2_X1 U1013 ( .A(n1334), .B(KEYINPUT53), .Z(n1335) );
XOR2_X1 U1014 ( .A(n1336), .B(KEYINPUT50), .Z(n1334) );
XOR2_X1 U1015 ( .A(n1132), .B(n1196), .Z(n1329) );
XNOR2_X1 U1016 ( .A(n1337), .B(n1338), .ZN(n1196) );
NOR2_X1 U1017 ( .A1(KEYINPUT22), .A2(n1136), .ZN(n1338) );
XNOR2_X1 U1018 ( .A(G131), .B(G137), .ZN(n1337) );
XOR2_X1 U1019 ( .A(G128), .B(n1339), .Z(n1132) );
AND2_X1 U1020 ( .A1(G227), .A2(n1340), .ZN(n1208) );
NOR2_X1 U1021 ( .A1(n1215), .A2(G110), .ZN(n1211) );
NAND2_X1 U1022 ( .A1(n1103), .A2(n1341), .ZN(n1064) );
NAND4_X1 U1023 ( .A1(G902), .A2(G953), .A3(n1291), .A4(n1151), .ZN(n1341) );
INV_X1 U1024 ( .A(G898), .ZN(n1151) );
NAND3_X1 U1025 ( .A1(n1342), .A2(n1291), .A3(n1071), .ZN(n1103) );
XNOR2_X1 U1026 ( .A(n1120), .B(KEYINPUT9), .ZN(n1071) );
NAND2_X1 U1027 ( .A1(G237), .A2(G234), .ZN(n1291) );
XOR2_X1 U1028 ( .A(KEYINPUT38), .B(G952), .Z(n1342) );
AND2_X1 U1029 ( .A1(n1343), .A2(n1275), .ZN(n1066) );
INV_X1 U1030 ( .A(n1090), .ZN(n1275) );
XNOR2_X1 U1031 ( .A(n1344), .B(n1222), .ZN(n1090) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1345), .ZN(n1222) );
NAND2_X1 U1033 ( .A1(n1346), .A2(n1223), .ZN(n1344) );
XOR2_X1 U1034 ( .A(n1218), .B(n1347), .Z(n1346) );
NOR2_X1 U1035 ( .A1(n1348), .A2(n1262), .ZN(n1347) );
NAND2_X1 U1036 ( .A1(n1349), .A2(n1350), .ZN(n1262) );
NAND2_X1 U1037 ( .A1(n1351), .A2(n1256), .ZN(n1350) );
XOR2_X1 U1038 ( .A(n1260), .B(n1194), .Z(n1351) );
NAND3_X1 U1039 ( .A1(n1261), .A2(n1192), .A3(G125), .ZN(n1349) );
INV_X1 U1040 ( .A(n1194), .ZN(n1192) );
INV_X1 U1041 ( .A(n1260), .ZN(n1261) );
NOR2_X1 U1042 ( .A1(n1256), .A2(n1255), .ZN(n1348) );
NAND2_X1 U1043 ( .A1(n1194), .A2(n1260), .ZN(n1255) );
NAND2_X1 U1044 ( .A1(G224), .A2(n1340), .ZN(n1260) );
XOR2_X1 U1045 ( .A(n1280), .B(n1352), .Z(n1194) );
NOR2_X1 U1046 ( .A1(KEYINPUT47), .A2(n1339), .ZN(n1352) );
XNOR2_X1 U1047 ( .A(n1353), .B(KEYINPUT43), .ZN(n1339) );
INV_X1 U1048 ( .A(G128), .ZN(n1280) );
XOR2_X1 U1049 ( .A(n1354), .B(n1160), .Z(n1218) );
INV_X1 U1050 ( .A(n1154), .ZN(n1160) );
XNOR2_X1 U1051 ( .A(G110), .B(n1355), .ZN(n1154) );
NOR2_X1 U1052 ( .A1(G122), .A2(KEYINPUT28), .ZN(n1355) );
XOR2_X1 U1053 ( .A(n1162), .B(n1356), .Z(n1354) );
NOR2_X1 U1054 ( .A1(KEYINPUT27), .A2(n1165), .ZN(n1356) );
NAND3_X1 U1055 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1165) );
NAND2_X1 U1056 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
INV_X1 U1057 ( .A(n1336), .ZN(n1360) );
OR3_X1 U1058 ( .A1(n1361), .A2(n1362), .A3(n1289), .ZN(n1358) );
INV_X1 U1059 ( .A(KEYINPUT32), .ZN(n1361) );
NAND2_X1 U1060 ( .A1(n1362), .A2(n1289), .ZN(n1357) );
INV_X1 U1061 ( .A(G101), .ZN(n1289) );
NAND2_X1 U1062 ( .A1(KEYINPUT62), .A2(n1336), .ZN(n1362) );
XOR2_X1 U1063 ( .A(n1182), .B(G107), .Z(n1336) );
INV_X1 U1064 ( .A(G104), .ZN(n1182) );
NAND3_X1 U1065 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1162) );
NAND2_X1 U1066 ( .A1(KEYINPUT51), .A2(G113), .ZN(n1365) );
OR3_X1 U1067 ( .A1(G113), .A2(KEYINPUT51), .A3(n1366), .ZN(n1364) );
NAND2_X1 U1068 ( .A1(n1366), .A2(n1367), .ZN(n1363) );
NAND2_X1 U1069 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
INV_X1 U1070 ( .A(KEYINPUT51), .ZN(n1369) );
XOR2_X1 U1071 ( .A(n1296), .B(KEYINPUT49), .Z(n1368) );
INV_X1 U1072 ( .A(G113), .ZN(n1296) );
XOR2_X1 U1073 ( .A(n1294), .B(n1293), .Z(n1366) );
INV_X1 U1074 ( .A(G119), .ZN(n1293) );
INV_X1 U1075 ( .A(G116), .ZN(n1294) );
XNOR2_X1 U1076 ( .A(n1091), .B(KEYINPUT36), .ZN(n1343) );
AND2_X1 U1077 ( .A1(G214), .A2(n1345), .ZN(n1091) );
NAND2_X1 U1078 ( .A1(n1370), .A2(n1223), .ZN(n1345) );
INV_X1 U1079 ( .A(G902), .ZN(n1223) );
NOR2_X1 U1080 ( .A1(n1270), .A2(n1267), .ZN(n1076) );
XNOR2_X1 U1081 ( .A(n1115), .B(n1371), .ZN(n1267) );
NOR2_X1 U1082 ( .A1(G475), .A2(KEYINPUT44), .ZN(n1371) );
NOR2_X1 U1083 ( .A1(n1180), .A2(G902), .ZN(n1115) );
XOR2_X1 U1084 ( .A(n1372), .B(G113), .Z(n1180) );
XOR2_X1 U1085 ( .A(n1373), .B(n1374), .Z(n1372) );
XOR2_X1 U1086 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1087 ( .A(G131), .B(G122), .Z(n1376) );
XOR2_X1 U1088 ( .A(KEYINPUT5), .B(KEYINPUT3), .Z(n1375) );
XOR2_X1 U1089 ( .A(n1377), .B(n1378), .Z(n1373) );
XOR2_X1 U1090 ( .A(n1353), .B(n1133), .Z(n1378) );
XOR2_X1 U1091 ( .A(n1215), .B(n1256), .Z(n1133) );
INV_X1 U1092 ( .A(G125), .ZN(n1256) );
INV_X1 U1093 ( .A(G140), .ZN(n1215) );
XNOR2_X1 U1094 ( .A(n1379), .B(G146), .ZN(n1353) );
XOR2_X1 U1095 ( .A(n1380), .B(G104), .Z(n1377) );
NAND2_X1 U1096 ( .A1(G214), .A2(n1316), .ZN(n1380) );
AND2_X1 U1097 ( .A1(n1340), .A2(n1370), .ZN(n1316) );
INV_X1 U1098 ( .A(G237), .ZN(n1370) );
INV_X1 U1099 ( .A(n1295), .ZN(n1270) );
XOR2_X1 U1100 ( .A(n1114), .B(n1113), .Z(n1295) );
NOR2_X1 U1101 ( .A1(n1174), .A2(G902), .ZN(n1113) );
XNOR2_X1 U1102 ( .A(n1381), .B(n1382), .ZN(n1174) );
NOR2_X1 U1103 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
XOR2_X1 U1104 ( .A(KEYINPUT40), .B(n1385), .Z(n1384) );
AND2_X1 U1105 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NOR2_X1 U1106 ( .A1(n1387), .A2(n1386), .ZN(n1383) );
XNOR2_X1 U1107 ( .A(n1136), .B(n1388), .ZN(n1386) );
NOR2_X1 U1108 ( .A1(KEYINPUT8), .A2(n1389), .ZN(n1388) );
XOR2_X1 U1109 ( .A(n1390), .B(G128), .Z(n1389) );
NAND2_X1 U1110 ( .A1(KEYINPUT34), .A2(n1379), .ZN(n1390) );
INV_X1 U1111 ( .A(G143), .ZN(n1379) );
INV_X1 U1112 ( .A(G134), .ZN(n1136) );
XOR2_X1 U1113 ( .A(G107), .B(n1391), .Z(n1387) );
XOR2_X1 U1114 ( .A(G122), .B(G116), .Z(n1391) );
NAND3_X1 U1115 ( .A1(n1307), .A2(G217), .A3(KEYINPUT13), .ZN(n1381) );
AND2_X1 U1116 ( .A1(n1340), .A2(G234), .ZN(n1307) );
XOR2_X1 U1117 ( .A(n1120), .B(KEYINPUT15), .Z(n1340) );
INV_X1 U1118 ( .A(G953), .ZN(n1120) );
INV_X1 U1119 ( .A(G478), .ZN(n1114) );
endmodule


