//Key = 1011001011111010010111011011111001101111010101000111010101100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350;

NOR4_X2 U751 ( .A1(n1052), .A2(n1050), .A3(n1054), .A4(n1051), .ZN(n1197) );
XOR2_X1 U752 ( .A(G107), .B(n1029), .Z(G9) );
NOR2_X1 U753 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NAND4_X1 U755 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1032) );
NAND4_X1 U756 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1037) );
NAND3_X1 U757 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U758 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XOR2_X1 U759 ( .A(n1049), .B(n1050), .Z(n1047) );
NAND2_X1 U760 ( .A1(KEYINPUT50), .A2(n1051), .ZN(n1049) );
NAND3_X1 U761 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1044) );
NAND2_X1 U762 ( .A1(n1048), .A2(n1055), .ZN(n1036) );
NAND2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND4_X1 U764 ( .A1(n1040), .A2(n1050), .A3(n1058), .A4(n1059), .ZN(n1057) );
NAND3_X1 U765 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1058) );
NAND2_X1 U766 ( .A1(n1063), .A2(n1042), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
XNOR2_X1 U768 ( .A(n1042), .B(KEYINPUT37), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1041), .A2(n1066), .ZN(n1060) );
XOR2_X1 U770 ( .A(n1067), .B(KEYINPUT32), .Z(n1056) );
NAND4_X1 U771 ( .A1(n1040), .A2(n1041), .A3(n1068), .A4(n1053), .ZN(n1067) );
INV_X1 U772 ( .A(n1069), .ZN(n1040) );
INV_X1 U773 ( .A(n1070), .ZN(n1048) );
AND3_X1 U774 ( .A1(n1038), .A2(n1039), .A3(n1071), .ZN(n1030) );
NAND4_X1 U775 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1038) );
NOR4_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
XNOR2_X1 U777 ( .A(G469), .B(n1080), .ZN(n1079) );
XOR2_X1 U778 ( .A(n1081), .B(KEYINPUT10), .Z(n1076) );
NOR3_X1 U779 ( .A1(n1054), .A2(n1082), .A3(n1051), .ZN(n1074) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(n1073) );
NOR2_X1 U781 ( .A1(n1085), .A2(KEYINPUT59), .ZN(n1084) );
XOR2_X1 U782 ( .A(KEYINPUT29), .B(n1086), .Z(n1072) );
XOR2_X1 U783 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1039), .ZN(n1088) );
AND2_X1 U785 ( .A1(G227), .A2(G900), .ZN(n1089) );
NAND3_X1 U786 ( .A1(KEYINPUT39), .A2(n1090), .A3(n1091), .ZN(n1087) );
XOR2_X1 U787 ( .A(n1092), .B(KEYINPUT44), .Z(n1091) );
NAND3_X1 U788 ( .A1(n1033), .A2(n1039), .A3(n1093), .ZN(n1092) );
INV_X1 U789 ( .A(n1094), .ZN(n1093) );
NAND3_X1 U790 ( .A1(n1095), .A2(n1096), .A3(n1094), .ZN(n1090) );
XNOR2_X1 U791 ( .A(n1097), .B(n1098), .ZN(n1094) );
XOR2_X1 U792 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U793 ( .A(n1101), .B(KEYINPUT51), .Z(n1100) );
NAND2_X1 U794 ( .A1(KEYINPUT28), .A2(G137), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1102), .B(n1103), .Z(n1097) );
XNOR2_X1 U796 ( .A(n1104), .B(n1105), .ZN(n1103) );
NOR2_X1 U797 ( .A1(G131), .A2(KEYINPUT13), .ZN(n1105) );
NAND2_X1 U798 ( .A1(KEYINPUT9), .A2(n1106), .ZN(n1104) );
NAND2_X1 U799 ( .A1(n1033), .A2(n1039), .ZN(n1096) );
NAND2_X1 U800 ( .A1(G953), .A2(n1107), .ZN(n1095) );
XOR2_X1 U801 ( .A(n1108), .B(n1109), .Z(G69) );
XOR2_X1 U802 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U803 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1112) );
NAND3_X1 U805 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1110) );
XOR2_X1 U806 ( .A(n1116), .B(KEYINPUT52), .Z(n1115) );
NAND2_X1 U807 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U808 ( .A1(G953), .A2(n1119), .ZN(n1114) );
OR2_X1 U809 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
XOR2_X1 U810 ( .A(n1120), .B(n1121), .Z(n1117) );
NAND2_X1 U811 ( .A1(KEYINPUT34), .A2(n1122), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1123), .A2(G953), .ZN(n1108) );
NOR2_X1 U813 ( .A1(n1029), .A2(n1034), .ZN(n1123) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XNOR2_X1 U815 ( .A(n1126), .B(n1127), .ZN(n1125) );
XOR2_X1 U816 ( .A(n1128), .B(KEYINPUT14), .Z(n1127) );
NAND2_X1 U817 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U818 ( .A1(n1124), .A2(n1131), .ZN(G63) );
XOR2_X1 U819 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U820 ( .A1(n1129), .A2(G478), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1124), .A2(n1134), .ZN(G60) );
XNOR2_X1 U822 ( .A(n1135), .B(n1136), .ZN(n1134) );
NAND2_X1 U823 ( .A1(n1129), .A2(G475), .ZN(n1135) );
XNOR2_X1 U824 ( .A(n1137), .B(n1138), .ZN(G6) );
NOR2_X1 U825 ( .A1(KEYINPUT35), .A2(n1139), .ZN(n1138) );
NOR4_X1 U826 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(G57) );
AND2_X1 U827 ( .A1(KEYINPUT58), .A2(n1124), .ZN(n1143) );
NOR3_X1 U828 ( .A1(KEYINPUT58), .A2(n1039), .A3(n1071), .ZN(n1142) );
INV_X1 U829 ( .A(G952), .ZN(n1071) );
NOR2_X1 U830 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
XOR2_X1 U831 ( .A(KEYINPUT30), .B(n1146), .Z(n1144) );
NOR2_X1 U832 ( .A1(n1147), .A2(n1148), .ZN(n1140) );
XNOR2_X1 U833 ( .A(n1146), .B(KEYINPUT11), .ZN(n1148) );
XNOR2_X1 U834 ( .A(n1149), .B(n1150), .ZN(n1146) );
XOR2_X1 U835 ( .A(KEYINPUT6), .B(G101), .Z(n1150) );
NAND2_X1 U836 ( .A1(n1151), .A2(KEYINPUT62), .ZN(n1149) );
XOR2_X1 U837 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U838 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U839 ( .A1(n1129), .A2(G472), .ZN(n1155) );
NAND2_X1 U840 ( .A1(KEYINPUT53), .A2(n1156), .ZN(n1154) );
INV_X1 U841 ( .A(n1145), .ZN(n1147) );
NOR2_X1 U842 ( .A1(n1124), .A2(n1157), .ZN(G54) );
XOR2_X1 U843 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U844 ( .A(KEYINPUT15), .B(n1160), .Z(n1159) );
NOR2_X1 U845 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U846 ( .A(KEYINPUT7), .B(n1163), .Z(n1162) );
AND2_X1 U847 ( .A1(n1164), .A2(n1156), .ZN(n1163) );
NOR2_X1 U848 ( .A1(n1156), .A2(n1164), .ZN(n1161) );
XOR2_X1 U849 ( .A(n1165), .B(n1166), .Z(n1158) );
NAND2_X1 U850 ( .A1(n1129), .A2(G469), .ZN(n1165) );
NOR2_X1 U851 ( .A1(n1124), .A2(n1167), .ZN(G51) );
XOR2_X1 U852 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U853 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR3_X1 U854 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1170) );
NOR2_X1 U855 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR3_X1 U856 ( .A1(G125), .A2(KEYINPUT47), .A3(n1177), .ZN(n1173) );
INV_X1 U857 ( .A(n1175), .ZN(n1177) );
NOR2_X1 U858 ( .A1(KEYINPUT22), .A2(n1178), .ZN(n1175) );
AND2_X1 U859 ( .A1(n1178), .A2(KEYINPUT47), .ZN(n1172) );
XOR2_X1 U860 ( .A(n1179), .B(n1180), .Z(n1168) );
NAND2_X1 U861 ( .A1(n1129), .A2(n1083), .ZN(n1179) );
AND2_X1 U862 ( .A1(G902), .A2(n1181), .ZN(n1129) );
OR3_X1 U863 ( .A1(n1035), .A2(n1034), .A3(n1033), .ZN(n1181) );
NAND4_X1 U864 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1033) );
NOR4_X1 U865 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
INV_X1 U866 ( .A(n1190), .ZN(n1186) );
NOR3_X1 U867 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1184) );
NOR2_X1 U868 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
AND4_X1 U869 ( .A1(n1194), .A2(n1196), .A3(n1197), .A4(n1063), .ZN(n1192) );
AND2_X1 U870 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
INV_X1 U871 ( .A(KEYINPUT43), .ZN(n1194) );
NOR2_X1 U872 ( .A1(n1070), .A2(n1200), .ZN(n1191) );
XNOR2_X1 U873 ( .A(KEYINPUT38), .B(n1201), .ZN(n1200) );
NAND4_X1 U874 ( .A1(n1202), .A2(n1203), .A3(n1139), .A4(n1204), .ZN(n1034) );
NOR4_X1 U875 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
INV_X1 U876 ( .A(n1209), .ZN(n1208) );
NAND3_X1 U877 ( .A1(n1197), .A2(n1210), .A3(n1065), .ZN(n1139) );
XOR2_X1 U878 ( .A(n1029), .B(KEYINPUT54), .Z(n1035) );
AND3_X1 U879 ( .A1(n1197), .A2(n1210), .A3(n1063), .ZN(n1029) );
NOR2_X1 U880 ( .A1(n1039), .A2(G952), .ZN(n1124) );
NAND2_X1 U881 ( .A1(n1211), .A2(n1212), .ZN(G48) );
NAND2_X1 U882 ( .A1(n1213), .A2(n1182), .ZN(n1212) );
NAND2_X1 U883 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U884 ( .A1(KEYINPUT25), .A2(KEYINPUT23), .ZN(n1215) );
NAND3_X1 U885 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1211) );
INV_X1 U886 ( .A(KEYINPUT25), .ZN(n1218) );
OR2_X1 U887 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1217) );
NAND2_X1 U888 ( .A1(KEYINPUT23), .A2(n1219), .ZN(n1216) );
OR2_X1 U889 ( .A1(n1182), .A2(G146), .ZN(n1219) );
NAND2_X1 U890 ( .A1(n1220), .A2(n1065), .ZN(n1182) );
XOR2_X1 U891 ( .A(G143), .B(n1189), .Z(G45) );
AND4_X1 U892 ( .A1(n1077), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1189) );
AND2_X1 U893 ( .A1(n1197), .A2(n1068), .ZN(n1223) );
XOR2_X1 U894 ( .A(G140), .B(n1188), .Z(G42) );
AND3_X1 U895 ( .A1(n1065), .A2(n1066), .A3(n1224), .ZN(n1188) );
NAND2_X1 U896 ( .A1(n1225), .A2(n1226), .ZN(G39) );
NAND2_X1 U897 ( .A1(G137), .A2(n1183), .ZN(n1226) );
XOR2_X1 U898 ( .A(KEYINPUT27), .B(n1227), .Z(n1225) );
NOR2_X1 U899 ( .A1(G137), .A2(n1183), .ZN(n1227) );
NAND3_X1 U900 ( .A1(n1199), .A2(n1224), .A3(n1041), .ZN(n1183) );
XOR2_X1 U901 ( .A(G134), .B(n1228), .Z(G36) );
NOR2_X1 U902 ( .A1(n1070), .A2(n1201), .ZN(n1228) );
NAND3_X1 U903 ( .A1(n1068), .A2(n1063), .A3(n1229), .ZN(n1201) );
NOR3_X1 U904 ( .A1(n1198), .A2(n1051), .A3(n1050), .ZN(n1229) );
XOR2_X1 U905 ( .A(G131), .B(n1187), .Z(G33) );
AND3_X1 U906 ( .A1(n1224), .A2(n1065), .A3(n1068), .ZN(n1187) );
NOR4_X1 U907 ( .A1(n1070), .A2(n1198), .A3(n1050), .A4(n1051), .ZN(n1224) );
INV_X1 U908 ( .A(n1221), .ZN(n1198) );
NAND2_X1 U909 ( .A1(n1052), .A2(n1230), .ZN(n1070) );
XOR2_X1 U910 ( .A(n1231), .B(n1195), .Z(G30) );
NAND2_X1 U911 ( .A1(n1220), .A2(n1063), .ZN(n1195) );
AND3_X1 U912 ( .A1(n1197), .A2(n1221), .A3(n1199), .ZN(n1220) );
XNOR2_X1 U913 ( .A(G101), .B(n1202), .ZN(G3) );
NAND4_X1 U914 ( .A1(n1041), .A2(n1068), .A3(n1197), .A4(n1232), .ZN(n1202) );
XOR2_X1 U915 ( .A(n1176), .B(n1190), .Z(G27) );
NAND4_X1 U916 ( .A1(n1065), .A2(n1233), .A3(n1066), .A4(n1221), .ZN(n1190) );
NAND2_X1 U917 ( .A1(n1069), .A2(n1234), .ZN(n1221) );
NAND2_X1 U918 ( .A1(n1235), .A2(n1107), .ZN(n1234) );
XOR2_X1 U919 ( .A(G900), .B(KEYINPUT63), .Z(n1107) );
XOR2_X1 U920 ( .A(n1236), .B(n1203), .Z(G24) );
NAND4_X1 U921 ( .A1(n1233), .A2(n1210), .A3(n1222), .A4(n1077), .ZN(n1203) );
AND2_X1 U922 ( .A1(n1042), .A2(n1232), .ZN(n1210) );
NOR2_X1 U923 ( .A1(n1237), .A2(n1238), .ZN(n1042) );
XOR2_X1 U924 ( .A(n1239), .B(n1209), .Z(G21) );
NAND3_X1 U925 ( .A1(n1041), .A2(n1199), .A3(n1240), .ZN(n1209) );
NOR2_X1 U926 ( .A1(n1241), .A2(n1242), .ZN(n1199) );
XOR2_X1 U927 ( .A(G116), .B(n1207), .Z(G18) );
AND3_X1 U928 ( .A1(n1068), .A2(n1063), .A3(n1240), .ZN(n1207) );
NOR2_X1 U929 ( .A1(n1077), .A2(n1081), .ZN(n1063) );
NAND2_X1 U930 ( .A1(n1243), .A2(n1244), .ZN(G15) );
NAND2_X1 U931 ( .A1(n1206), .A2(n1245), .ZN(n1244) );
XOR2_X1 U932 ( .A(KEYINPUT26), .B(n1246), .Z(n1243) );
NOR2_X1 U933 ( .A1(n1206), .A2(n1245), .ZN(n1246) );
AND3_X1 U934 ( .A1(n1068), .A2(n1065), .A3(n1240), .ZN(n1206) );
AND2_X1 U935 ( .A1(n1233), .A2(n1232), .ZN(n1240) );
INV_X1 U936 ( .A(n1045), .ZN(n1233) );
NAND3_X1 U937 ( .A1(n1247), .A2(n1230), .A3(n1053), .ZN(n1045) );
NOR2_X1 U938 ( .A1(n1248), .A2(n1051), .ZN(n1053) );
INV_X1 U939 ( .A(n1052), .ZN(n1247) );
AND2_X1 U940 ( .A1(n1081), .A2(n1077), .ZN(n1065) );
NOR2_X1 U941 ( .A1(n1238), .A2(n1242), .ZN(n1068) );
XOR2_X1 U942 ( .A(n1249), .B(n1250), .Z(G12) );
NAND2_X1 U943 ( .A1(KEYINPUT33), .A2(n1205), .ZN(n1250) );
AND4_X1 U944 ( .A1(n1041), .A2(n1066), .A3(n1197), .A4(n1232), .ZN(n1205) );
NAND2_X1 U945 ( .A1(n1069), .A2(n1251), .ZN(n1232) );
NAND2_X1 U946 ( .A1(n1235), .A2(n1119), .ZN(n1251) );
XOR2_X1 U947 ( .A(KEYINPUT19), .B(G898), .Z(n1119) );
AND3_X1 U948 ( .A1(G902), .A2(n1252), .A3(G953), .ZN(n1235) );
NAND3_X1 U949 ( .A1(n1252), .A2(n1039), .A3(G952), .ZN(n1069) );
NAND2_X1 U950 ( .A1(G237), .A2(G234), .ZN(n1252) );
INV_X1 U951 ( .A(n1059), .ZN(n1051) );
NAND2_X1 U952 ( .A1(G221), .A2(n1253), .ZN(n1059) );
INV_X1 U953 ( .A(n1230), .ZN(n1054) );
NAND2_X1 U954 ( .A1(G214), .A2(n1254), .ZN(n1230) );
INV_X1 U955 ( .A(n1248), .ZN(n1050) );
NAND2_X1 U956 ( .A1(n1255), .A2(n1256), .ZN(n1248) );
OR2_X1 U957 ( .A1(n1080), .A2(G469), .ZN(n1256) );
XOR2_X1 U958 ( .A(n1257), .B(KEYINPUT48), .Z(n1255) );
NAND2_X1 U959 ( .A1(G469), .A2(n1080), .ZN(n1257) );
NAND2_X1 U960 ( .A1(n1258), .A2(n1259), .ZN(n1080) );
XNOR2_X1 U961 ( .A(n1166), .B(n1260), .ZN(n1258) );
XNOR2_X1 U962 ( .A(n1164), .B(n1156), .ZN(n1260) );
XNOR2_X1 U963 ( .A(n1261), .B(n1178), .ZN(n1164) );
NAND2_X1 U964 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U965 ( .A(n1264), .B(n1265), .ZN(n1166) );
XOR2_X1 U966 ( .A(G140), .B(G110), .Z(n1265) );
NAND2_X1 U967 ( .A1(G227), .A2(n1039), .ZN(n1264) );
XOR2_X1 U968 ( .A(n1266), .B(n1083), .Z(n1052) );
AND2_X1 U969 ( .A1(G210), .A2(n1254), .ZN(n1083) );
NAND2_X1 U970 ( .A1(n1267), .A2(n1259), .ZN(n1254) );
XNOR2_X1 U971 ( .A(n1085), .B(KEYINPUT56), .ZN(n1266) );
AND3_X1 U972 ( .A1(n1268), .A2(n1259), .A3(n1269), .ZN(n1085) );
XOR2_X1 U973 ( .A(KEYINPUT41), .B(n1270), .Z(n1269) );
NOR2_X1 U974 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U975 ( .A1(n1271), .A2(n1272), .ZN(n1268) );
XOR2_X1 U976 ( .A(n1273), .B(n1102), .Z(n1272) );
XOR2_X1 U977 ( .A(n1176), .B(n1180), .Z(n1273) );
AND2_X1 U978 ( .A1(G224), .A2(n1039), .ZN(n1180) );
XOR2_X1 U979 ( .A(n1171), .B(KEYINPUT18), .Z(n1271) );
XNOR2_X1 U980 ( .A(n1274), .B(n1275), .ZN(n1171) );
XOR2_X1 U981 ( .A(n1118), .B(n1121), .Z(n1275) );
NAND2_X1 U982 ( .A1(n1276), .A2(n1277), .ZN(n1118) );
NAND2_X1 U983 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND2_X1 U984 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U985 ( .A1(G110), .A2(n1282), .ZN(n1281) );
INV_X1 U986 ( .A(KEYINPUT4), .ZN(n1280) );
NAND2_X1 U987 ( .A1(n1283), .A2(n1249), .ZN(n1276) );
NAND2_X1 U988 ( .A1(n1282), .A2(n1284), .ZN(n1283) );
OR2_X1 U989 ( .A1(n1278), .A2(KEYINPUT4), .ZN(n1284) );
XOR2_X1 U990 ( .A(n1236), .B(KEYINPUT12), .Z(n1278) );
INV_X1 U991 ( .A(G122), .ZN(n1236) );
INV_X1 U992 ( .A(KEYINPUT5), .ZN(n1282) );
XNOR2_X1 U993 ( .A(n1122), .B(KEYINPUT46), .ZN(n1274) );
AND2_X1 U994 ( .A1(n1285), .A2(n1263), .ZN(n1122) );
NAND2_X1 U995 ( .A1(G101), .A2(n1286), .ZN(n1263) );
XNOR2_X1 U996 ( .A(KEYINPUT0), .B(n1262), .ZN(n1285) );
OR2_X1 U997 ( .A1(n1286), .A2(G101), .ZN(n1262) );
XOR2_X1 U998 ( .A(G107), .B(G104), .Z(n1286) );
NOR2_X1 U999 ( .A1(n1241), .A2(n1237), .ZN(n1066) );
INV_X1 U1000 ( .A(n1242), .ZN(n1237) );
NOR2_X1 U1001 ( .A1(n1287), .A2(n1086), .ZN(n1242) );
NOR2_X1 U1002 ( .A1(n1288), .A2(G472), .ZN(n1086) );
XNOR2_X1 U1003 ( .A(KEYINPUT45), .B(n1082), .ZN(n1287) );
AND2_X1 U1004 ( .A1(G472), .A2(n1288), .ZN(n1082) );
NAND2_X1 U1005 ( .A1(n1289), .A2(n1259), .ZN(n1288) );
XOR2_X1 U1006 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1007 ( .A(n1152), .B(n1156), .Z(n1291) );
XNOR2_X1 U1008 ( .A(n1292), .B(n1293), .ZN(n1156) );
XOR2_X1 U1009 ( .A(KEYINPUT57), .B(G131), .Z(n1293) );
NAND2_X1 U1010 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
NAND2_X1 U1011 ( .A1(G137), .A2(n1101), .ZN(n1295) );
XOR2_X1 U1012 ( .A(n1296), .B(KEYINPUT31), .Z(n1294) );
OR2_X1 U1013 ( .A1(n1101), .A2(G137), .ZN(n1296) );
INV_X1 U1014 ( .A(G134), .ZN(n1101) );
XOR2_X1 U1015 ( .A(n1121), .B(n1178), .Z(n1152) );
INV_X1 U1016 ( .A(n1102), .ZN(n1178) );
XOR2_X1 U1017 ( .A(n1231), .B(n1297), .Z(n1102) );
XOR2_X1 U1018 ( .A(G146), .B(G143), .Z(n1297) );
INV_X1 U1019 ( .A(G128), .ZN(n1231) );
XOR2_X1 U1020 ( .A(n1245), .B(n1298), .Z(n1121) );
XOR2_X1 U1021 ( .A(G119), .B(G116), .Z(n1298) );
XOR2_X1 U1022 ( .A(n1145), .B(G101), .Z(n1290) );
NAND3_X1 U1023 ( .A1(n1267), .A2(n1039), .A3(G210), .ZN(n1145) );
INV_X1 U1024 ( .A(n1238), .ZN(n1241) );
XNOR2_X1 U1025 ( .A(n1078), .B(KEYINPUT20), .ZN(n1238) );
XNOR2_X1 U1026 ( .A(n1299), .B(n1130), .ZN(n1078) );
AND2_X1 U1027 ( .A1(G217), .A2(n1253), .ZN(n1130) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1259), .ZN(n1253) );
NAND2_X1 U1029 ( .A1(n1126), .A2(n1259), .ZN(n1299) );
XNOR2_X1 U1030 ( .A(n1300), .B(n1301), .ZN(n1126) );
XNOR2_X1 U1031 ( .A(n1302), .B(n1303), .ZN(n1301) );
NAND2_X1 U1032 ( .A1(n1304), .A2(KEYINPUT8), .ZN(n1302) );
XOR2_X1 U1033 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1034 ( .A(G128), .B(G110), .Z(n1306) );
NAND2_X1 U1035 ( .A1(KEYINPUT17), .A2(n1239), .ZN(n1305) );
INV_X1 U1036 ( .A(G119), .ZN(n1239) );
XOR2_X1 U1037 ( .A(n1307), .B(G137), .Z(n1300) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1308), .ZN(n1307) );
NOR2_X1 U1039 ( .A1(n1222), .A2(n1077), .ZN(n1041) );
XOR2_X1 U1040 ( .A(G475), .B(n1309), .Z(n1077) );
NOR2_X1 U1041 ( .A1(G902), .A2(n1136), .ZN(n1309) );
NAND2_X1 U1042 ( .A1(n1310), .A2(n1311), .ZN(n1136) );
NAND2_X1 U1043 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1044 ( .A1(KEYINPUT55), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1045 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U1046 ( .A(n1317), .B(n1318), .Z(n1315) );
XOR2_X1 U1047 ( .A(n1319), .B(n1303), .Z(n1312) );
NAND2_X1 U1048 ( .A1(n1320), .A2(n1321), .ZN(n1310) );
NAND2_X1 U1049 ( .A1(n1322), .A2(n1316), .ZN(n1321) );
INV_X1 U1050 ( .A(KEYINPUT1), .ZN(n1316) );
NAND2_X1 U1051 ( .A1(n1323), .A2(KEYINPUT55), .ZN(n1322) );
XNOR2_X1 U1052 ( .A(n1303), .B(n1319), .ZN(n1323) );
NOR2_X1 U1053 ( .A1(KEYINPUT60), .A2(n1324), .ZN(n1319) );
XOR2_X1 U1054 ( .A(n1325), .B(n1326), .Z(n1324) );
NAND4_X1 U1055 ( .A1(KEYINPUT3), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1326) );
NAND3_X1 U1056 ( .A1(KEYINPUT61), .A2(n1330), .A3(n1331), .ZN(n1329) );
OR2_X1 U1057 ( .A1(n1331), .A2(n1330), .ZN(n1328) );
NOR2_X1 U1058 ( .A1(KEYINPUT16), .A2(n1332), .ZN(n1330) );
INV_X1 U1059 ( .A(G143), .ZN(n1331) );
NAND2_X1 U1060 ( .A1(n1332), .A2(n1333), .ZN(n1327) );
INV_X1 U1061 ( .A(KEYINPUT61), .ZN(n1333) );
NAND3_X1 U1062 ( .A1(n1267), .A2(n1039), .A3(G214), .ZN(n1332) );
INV_X1 U1063 ( .A(G237), .ZN(n1267) );
INV_X1 U1064 ( .A(G131), .ZN(n1325) );
XOR2_X1 U1065 ( .A(n1214), .B(n1106), .Z(n1303) );
XOR2_X1 U1066 ( .A(G140), .B(n1176), .Z(n1106) );
INV_X1 U1067 ( .A(G125), .ZN(n1176) );
INV_X1 U1068 ( .A(G146), .ZN(n1214) );
XNOR2_X1 U1069 ( .A(n1318), .B(n1317), .ZN(n1320) );
NAND2_X1 U1070 ( .A1(KEYINPUT36), .A2(n1137), .ZN(n1317) );
INV_X1 U1071 ( .A(G104), .ZN(n1137) );
XOR2_X1 U1072 ( .A(n1334), .B(G122), .Z(n1318) );
NAND2_X1 U1073 ( .A1(KEYINPUT49), .A2(n1245), .ZN(n1334) );
INV_X1 U1074 ( .A(G113), .ZN(n1245) );
INV_X1 U1075 ( .A(n1081), .ZN(n1222) );
XOR2_X1 U1076 ( .A(n1335), .B(G478), .Z(n1081) );
NAND2_X1 U1077 ( .A1(n1133), .A2(n1259), .ZN(n1335) );
INV_X1 U1078 ( .A(G902), .ZN(n1259) );
XOR2_X1 U1079 ( .A(n1336), .B(n1337), .Z(n1133) );
XOR2_X1 U1080 ( .A(n1338), .B(n1339), .Z(n1337) );
NAND2_X1 U1081 ( .A1(KEYINPUT24), .A2(G134), .ZN(n1339) );
NAND3_X1 U1082 ( .A1(G217), .A2(n1308), .A3(KEYINPUT2), .ZN(n1338) );
AND2_X1 U1083 ( .A1(G234), .A2(n1039), .ZN(n1308) );
INV_X1 U1084 ( .A(G953), .ZN(n1039) );
XOR2_X1 U1085 ( .A(n1340), .B(n1341), .Z(n1336) );
NOR2_X1 U1086 ( .A1(G128), .A2(KEYINPUT40), .ZN(n1341) );
XOR2_X1 U1087 ( .A(n1342), .B(G143), .Z(n1340) );
NAND3_X1 U1088 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1342) );
OR2_X1 U1089 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND3_X1 U1090 ( .A1(n1347), .A2(n1346), .A3(G107), .ZN(n1344) );
NAND2_X1 U1091 ( .A1(n1348), .A2(n1349), .ZN(n1343) );
INV_X1 U1092 ( .A(G107), .ZN(n1349) );
NAND2_X1 U1093 ( .A1(n1350), .A2(n1346), .ZN(n1348) );
INV_X1 U1094 ( .A(KEYINPUT42), .ZN(n1346) );
XNOR2_X1 U1095 ( .A(n1347), .B(KEYINPUT21), .ZN(n1350) );
XOR2_X1 U1096 ( .A(G116), .B(G122), .Z(n1347) );
INV_X1 U1097 ( .A(G110), .ZN(n1249) );
endmodule


