//Key = 0101101010110101010010111000010101010000100001101010001111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350;

XNOR2_X1 U762 ( .A(G107), .B(n1040), .ZN(G9) );
NAND4_X1 U763 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
NOR2_X1 U764 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND3_X1 U766 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND4_X1 U767 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NAND2_X1 U768 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND2_X1 U769 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U770 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND3_X1 U771 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
INV_X1 U772 ( .A(KEYINPUT22), .ZN(n1064) );
NAND2_X1 U773 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
OR2_X1 U774 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U775 ( .A1(n1043), .A2(n1070), .ZN(n1057) );
NAND2_X1 U776 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U777 ( .A1(n1059), .A2(n1073), .ZN(n1072) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U779 ( .A1(KEYINPUT22), .A2(n1065), .ZN(n1075) );
NAND2_X1 U780 ( .A1(n1066), .A2(n1076), .ZN(n1071) );
NAND2_X1 U781 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U782 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
INV_X1 U783 ( .A(n1082), .ZN(n1081) );
INV_X1 U784 ( .A(n1083), .ZN(n1054) );
NAND4_X1 U785 ( .A1(n1043), .A2(n1084), .A3(n1066), .A4(n1085), .ZN(n1050) );
NOR2_X1 U786 ( .A1(n1086), .A2(n1083), .ZN(n1085) );
NAND2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
XOR2_X1 U788 ( .A(KEYINPUT58), .B(n1089), .Z(n1087) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1056), .ZN(n1089) );
NOR3_X1 U790 ( .A1(n1048), .A2(G952), .A3(n1091), .ZN(n1045) );
INV_X1 U791 ( .A(n1051), .ZN(n1091) );
NAND4_X1 U792 ( .A1(n1092), .A2(n1080), .A3(n1093), .A4(n1094), .ZN(n1051) );
NOR4_X1 U793 ( .A1(n1090), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1094) );
XOR2_X1 U794 ( .A(G478), .B(n1098), .Z(n1097) );
XNOR2_X1 U795 ( .A(G472), .B(n1099), .ZN(n1096) );
XNOR2_X1 U796 ( .A(n1100), .B(n1101), .ZN(n1095) );
XNOR2_X1 U797 ( .A(n1102), .B(KEYINPUT52), .ZN(n1101) );
AND3_X1 U798 ( .A1(n1103), .A2(n1056), .A3(n1082), .ZN(n1093) );
INV_X1 U799 ( .A(n1104), .ZN(n1048) );
XOR2_X1 U800 ( .A(n1105), .B(n1106), .Z(G72) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
AND2_X1 U802 ( .A1(G227), .A2(G900), .ZN(n1107) );
NAND2_X1 U803 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NAND2_X1 U804 ( .A1(n1111), .A2(n1108), .ZN(n1110) );
XNOR2_X1 U805 ( .A(n1112), .B(n1113), .ZN(n1111) );
NAND3_X1 U806 ( .A1(G900), .A2(n1113), .A3(G953), .ZN(n1109) );
XOR2_X1 U807 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U808 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U809 ( .A(n1118), .B(n1119), .ZN(n1114) );
NAND2_X1 U810 ( .A1(KEYINPUT46), .A2(n1120), .ZN(n1118) );
XOR2_X1 U811 ( .A(n1121), .B(n1122), .Z(G69) );
XOR2_X1 U812 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U814 ( .A1(n1127), .A2(n1125), .ZN(n1123) );
NOR2_X1 U815 ( .A1(G224), .A2(n1108), .ZN(n1127) );
NAND2_X1 U816 ( .A1(n1108), .A2(n1128), .ZN(n1121) );
NAND3_X1 U817 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
XOR2_X1 U818 ( .A(n1132), .B(KEYINPUT43), .Z(n1131) );
NOR2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U821 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U822 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U824 ( .A1(G478), .A2(n1142), .ZN(n1141) );
NAND2_X1 U825 ( .A1(KEYINPUT11), .A2(n1143), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1133), .A2(n1144), .ZN(G60) );
NOR3_X1 U827 ( .A1(n1102), .A2(n1145), .A3(n1146), .ZN(n1144) );
AND3_X1 U828 ( .A1(n1147), .A2(G475), .A3(n1142), .ZN(n1146) );
INV_X1 U829 ( .A(n1138), .ZN(n1142) );
NOR2_X1 U830 ( .A1(n1148), .A2(n1147), .ZN(n1145) );
AND2_X1 U831 ( .A1(n1049), .A2(G475), .ZN(n1148) );
XNOR2_X1 U832 ( .A(G104), .B(n1149), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1133), .A2(n1150), .ZN(G57) );
XOR2_X1 U834 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
OR3_X1 U836 ( .A1(n1138), .A2(n1155), .A3(n1156), .ZN(n1154) );
NAND2_X1 U837 ( .A1(n1157), .A2(n1156), .ZN(n1153) );
XNOR2_X1 U838 ( .A(n1158), .B(n1159), .ZN(n1156) );
NAND2_X1 U839 ( .A1(KEYINPUT40), .A2(n1160), .ZN(n1158) );
XOR2_X1 U840 ( .A(KEYINPUT29), .B(n1161), .Z(n1157) );
NOR2_X1 U841 ( .A1(n1155), .A2(n1138), .ZN(n1161) );
NOR3_X1 U842 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(G54) );
AND2_X1 U843 ( .A1(KEYINPUT31), .A2(n1133), .ZN(n1164) );
NOR3_X1 U844 ( .A1(KEYINPUT31), .A2(G953), .A3(G952), .ZN(n1163) );
NOR2_X1 U845 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
XOR2_X1 U846 ( .A(KEYINPUT16), .B(n1167), .Z(n1166) );
AND2_X1 U847 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U848 ( .A1(n1169), .A2(n1168), .ZN(n1165) );
XNOR2_X1 U849 ( .A(n1170), .B(n1171), .ZN(n1168) );
NAND2_X1 U850 ( .A1(n1172), .A2(KEYINPUT13), .ZN(n1170) );
XOR2_X1 U851 ( .A(n1173), .B(n1116), .Z(n1172) );
NOR2_X1 U852 ( .A1(KEYINPUT32), .A2(n1174), .ZN(n1173) );
NOR2_X1 U853 ( .A1(n1138), .A2(n1175), .ZN(n1169) );
NOR2_X1 U854 ( .A1(n1133), .A2(n1176), .ZN(G51) );
NOR2_X1 U855 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U856 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U857 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U858 ( .A1(n1183), .A2(n1138), .ZN(n1179) );
NAND2_X1 U859 ( .A1(G902), .A2(n1049), .ZN(n1138) );
NAND4_X1 U860 ( .A1(n1184), .A2(n1112), .A3(n1129), .A4(n1132), .ZN(n1049) );
AND4_X1 U861 ( .A1(n1149), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1129) );
AND3_X1 U862 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NAND4_X1 U863 ( .A1(n1059), .A2(n1068), .A3(n1041), .A4(n1042), .ZN(n1186) );
NAND4_X1 U864 ( .A1(n1065), .A2(n1041), .A3(n1043), .A4(n1044), .ZN(n1149) );
AND4_X1 U865 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1112) );
NOR4_X1 U866 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR2_X1 U867 ( .A1(n1088), .A2(n1199), .ZN(n1198) );
NOR3_X1 U868 ( .A1(n1200), .A2(n1201), .A3(n1074), .ZN(n1195) );
XNOR2_X1 U869 ( .A(n1202), .B(KEYINPUT0), .ZN(n1201) );
NOR2_X1 U870 ( .A1(n1203), .A2(n1204), .ZN(n1193) );
XOR2_X1 U871 ( .A(n1130), .B(KEYINPUT5), .Z(n1184) );
NAND4_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1044), .A4(n1207), .ZN(n1130) );
NOR2_X1 U873 ( .A1(n1063), .A2(n1074), .ZN(n1207) );
XNOR2_X1 U874 ( .A(KEYINPUT9), .B(n1088), .ZN(n1205) );
AND2_X1 U875 ( .A1(n1182), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U876 ( .A(n1208), .B(n1209), .ZN(n1181) );
XNOR2_X1 U877 ( .A(n1210), .B(n1126), .ZN(n1209) );
INV_X1 U878 ( .A(n1211), .ZN(n1126) );
XNOR2_X1 U879 ( .A(G125), .B(n1212), .ZN(n1208) );
INV_X1 U880 ( .A(KEYINPUT3), .ZN(n1182) );
NOR2_X1 U881 ( .A1(n1108), .A2(G952), .ZN(n1133) );
XNOR2_X1 U882 ( .A(G146), .B(n1191), .ZN(G48) );
NAND3_X1 U883 ( .A1(n1213), .A2(n1065), .A3(n1202), .ZN(n1191) );
XNOR2_X1 U884 ( .A(G143), .B(n1192), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1213), .A2(n1068), .A3(n1214), .A4(n1215), .ZN(n1192) );
INV_X1 U886 ( .A(n1200), .ZN(n1213) );
NAND3_X1 U887 ( .A1(n1216), .A2(n1217), .A3(n1044), .ZN(n1200) );
XNOR2_X1 U888 ( .A(n1197), .B(n1218), .ZN(G42) );
NOR2_X1 U889 ( .A1(G140), .A2(KEYINPUT44), .ZN(n1218) );
AND3_X1 U890 ( .A1(n1065), .A2(n1219), .A3(n1069), .ZN(n1197) );
XNOR2_X1 U891 ( .A(G137), .B(n1220), .ZN(G39) );
NAND2_X1 U892 ( .A1(KEYINPUT57), .A2(n1196), .ZN(n1220) );
AND3_X1 U893 ( .A1(n1202), .A2(n1219), .A3(n1066), .ZN(n1196) );
XOR2_X1 U894 ( .A(n1221), .B(n1204), .Z(G36) );
AND3_X1 U895 ( .A1(n1068), .A2(n1042), .A3(n1219), .ZN(n1204) );
XNOR2_X1 U896 ( .A(G134), .B(KEYINPUT15), .ZN(n1221) );
XNOR2_X1 U897 ( .A(n1119), .B(n1203), .ZN(G33) );
AND3_X1 U898 ( .A1(n1219), .A2(n1068), .A3(n1065), .ZN(n1203) );
AND4_X1 U899 ( .A1(n1053), .A2(n1044), .A3(n1217), .A4(n1056), .ZN(n1219) );
INV_X1 U900 ( .A(n1090), .ZN(n1053) );
XNOR2_X1 U901 ( .A(G128), .B(n1222), .ZN(G30) );
NAND2_X1 U902 ( .A1(n1223), .A2(n1216), .ZN(n1222) );
XOR2_X1 U903 ( .A(n1224), .B(KEYINPUT8), .Z(n1223) );
NAND4_X1 U904 ( .A1(n1042), .A2(n1044), .A3(n1225), .A4(n1217), .ZN(n1224) );
XOR2_X1 U905 ( .A(KEYINPUT53), .B(n1202), .Z(n1225) );
INV_X1 U906 ( .A(n1074), .ZN(n1042) );
XNOR2_X1 U907 ( .A(n1185), .B(n1226), .ZN(G3) );
NOR2_X1 U908 ( .A1(KEYINPUT37), .A2(n1227), .ZN(n1226) );
NAND3_X1 U909 ( .A1(n1068), .A2(n1044), .A3(n1228), .ZN(n1185) );
XNOR2_X1 U910 ( .A(G125), .B(n1229), .ZN(G27) );
NAND2_X1 U911 ( .A1(n1230), .A2(n1216), .ZN(n1229) );
XOR2_X1 U912 ( .A(n1199), .B(KEYINPUT48), .Z(n1230) );
NAND4_X1 U913 ( .A1(n1059), .A2(n1069), .A3(n1065), .A4(n1217), .ZN(n1199) );
NAND2_X1 U914 ( .A1(n1083), .A2(n1231), .ZN(n1217) );
NAND4_X1 U915 ( .A1(G902), .A2(G953), .A3(n1232), .A4(n1233), .ZN(n1231) );
INV_X1 U916 ( .A(G900), .ZN(n1233) );
XNOR2_X1 U917 ( .A(G122), .B(n1188), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1214), .A2(n1043), .A3(n1041), .A4(n1234), .ZN(n1188) );
NOR2_X1 U919 ( .A1(n1086), .A2(n1235), .ZN(n1234) );
INV_X1 U920 ( .A(n1063), .ZN(n1043) );
NAND2_X1 U921 ( .A1(n1092), .A2(n1236), .ZN(n1063) );
XNOR2_X1 U922 ( .A(n1237), .B(n1190), .ZN(G21) );
NAND3_X1 U923 ( .A1(n1059), .A2(n1202), .A3(n1228), .ZN(n1190) );
NOR2_X1 U924 ( .A1(n1236), .A2(n1092), .ZN(n1202) );
NAND2_X1 U925 ( .A1(KEYINPUT61), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U926 ( .A(G116), .B(n1239), .ZN(G18) );
NAND4_X1 U927 ( .A1(KEYINPUT50), .A2(n1068), .A3(n1240), .A4(n1041), .ZN(n1239) );
NOR2_X1 U928 ( .A1(n1241), .A2(n1074), .ZN(n1240) );
NAND2_X1 U929 ( .A1(n1214), .A2(n1235), .ZN(n1074) );
XNOR2_X1 U930 ( .A(n1059), .B(KEYINPUT28), .ZN(n1241) );
XNOR2_X1 U931 ( .A(n1242), .B(n1132), .ZN(G15) );
NAND4_X1 U932 ( .A1(n1059), .A2(n1065), .A3(n1068), .A4(n1041), .ZN(n1132) );
AND2_X1 U933 ( .A1(n1243), .A2(n1244), .ZN(n1068) );
XOR2_X1 U934 ( .A(n1092), .B(KEYINPUT62), .Z(n1243) );
NOR2_X1 U935 ( .A1(n1235), .A2(n1214), .ZN(n1065) );
INV_X1 U936 ( .A(n1086), .ZN(n1059) );
NAND3_X1 U937 ( .A1(n1080), .A2(n1082), .A3(n1079), .ZN(n1086) );
NAND2_X1 U938 ( .A1(KEYINPUT55), .A2(n1245), .ZN(n1242) );
XNOR2_X1 U939 ( .A(G110), .B(n1189), .ZN(G12) );
NAND3_X1 U940 ( .A1(n1069), .A2(n1044), .A3(n1228), .ZN(n1189) );
AND2_X1 U941 ( .A1(n1066), .A2(n1041), .ZN(n1228) );
AND2_X1 U942 ( .A1(n1216), .A2(n1206), .ZN(n1041) );
NAND2_X1 U943 ( .A1(n1083), .A2(n1246), .ZN(n1206) );
NAND3_X1 U944 ( .A1(n1125), .A2(n1232), .A3(G902), .ZN(n1246) );
NOR2_X1 U945 ( .A1(G898), .A2(n1108), .ZN(n1125) );
NAND3_X1 U946 ( .A1(n1104), .A2(n1232), .A3(G952), .ZN(n1083) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1232) );
XOR2_X1 U948 ( .A(G953), .B(KEYINPUT24), .Z(n1104) );
INV_X1 U949 ( .A(n1088), .ZN(n1216) );
NAND2_X1 U950 ( .A1(n1090), .A2(n1056), .ZN(n1088) );
NAND2_X1 U951 ( .A1(G214), .A2(n1247), .ZN(n1056) );
XOR2_X1 U952 ( .A(n1248), .B(n1183), .Z(n1090) );
NAND2_X1 U953 ( .A1(G210), .A2(n1247), .ZN(n1183) );
NAND2_X1 U954 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
INV_X1 U955 ( .A(G237), .ZN(n1249) );
NAND2_X1 U956 ( .A1(n1251), .A2(n1250), .ZN(n1248) );
XOR2_X1 U957 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U958 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U959 ( .A(KEYINPUT41), .B(G125), .Z(n1255) );
NOR2_X1 U960 ( .A1(KEYINPUT19), .A2(n1211), .ZN(n1254) );
XNOR2_X1 U961 ( .A(n1256), .B(n1257), .ZN(n1211) );
XOR2_X1 U962 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U963 ( .A(n1260), .B(n1261), .ZN(n1259) );
NOR2_X1 U964 ( .A1(KEYINPUT38), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U965 ( .A(n1263), .B(n1238), .ZN(n1262) );
NAND2_X1 U966 ( .A1(KEYINPUT20), .A2(G116), .ZN(n1263) );
NAND2_X1 U967 ( .A1(KEYINPUT6), .A2(n1264), .ZN(n1260) );
XNOR2_X1 U968 ( .A(KEYINPUT17), .B(n1265), .ZN(n1258) );
XOR2_X1 U969 ( .A(n1266), .B(n1267), .Z(n1256) );
XNOR2_X1 U970 ( .A(n1268), .B(n1269), .ZN(n1266) );
NOR2_X1 U971 ( .A1(KEYINPUT30), .A2(n1227), .ZN(n1269) );
INV_X1 U972 ( .A(G101), .ZN(n1227) );
NOR2_X1 U973 ( .A1(G107), .A2(KEYINPUT7), .ZN(n1268) );
XNOR2_X1 U974 ( .A(n1212), .B(n1270), .ZN(n1252) );
NOR2_X1 U975 ( .A1(KEYINPUT63), .A2(n1210), .ZN(n1270) );
AND2_X1 U976 ( .A1(G224), .A2(n1108), .ZN(n1212) );
NOR2_X1 U977 ( .A1(n1215), .A2(n1214), .ZN(n1066) );
XNOR2_X1 U978 ( .A(G478), .B(n1271), .ZN(n1214) );
NOR2_X1 U979 ( .A1(n1098), .A2(KEYINPUT34), .ZN(n1271) );
AND2_X1 U980 ( .A1(n1143), .A2(n1250), .ZN(n1098) );
XOR2_X1 U981 ( .A(n1272), .B(n1273), .Z(n1143) );
XNOR2_X1 U982 ( .A(n1274), .B(n1275), .ZN(n1273) );
NOR2_X1 U983 ( .A1(G122), .A2(KEYINPUT27), .ZN(n1275) );
NAND3_X1 U984 ( .A1(G234), .A2(n1108), .A3(G217), .ZN(n1274) );
XNOR2_X1 U985 ( .A(n1276), .B(n1277), .ZN(n1272) );
XOR2_X1 U986 ( .A(G116), .B(G107), .Z(n1277) );
NAND4_X1 U987 ( .A1(KEYINPUT60), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(n1276) );
OR3_X1 U988 ( .A1(n1281), .A2(G134), .A3(KEYINPUT2), .ZN(n1280) );
NAND2_X1 U989 ( .A1(KEYINPUT2), .A2(n1282), .ZN(n1279) );
NAND2_X1 U990 ( .A1(G134), .A2(n1281), .ZN(n1278) );
NAND2_X1 U991 ( .A1(KEYINPUT54), .A2(n1283), .ZN(n1281) );
INV_X1 U992 ( .A(n1282), .ZN(n1283) );
XOR2_X1 U993 ( .A(G143), .B(n1284), .Z(n1282) );
INV_X1 U994 ( .A(G128), .ZN(n1284) );
INV_X1 U995 ( .A(n1235), .ZN(n1215) );
XOR2_X1 U996 ( .A(n1102), .B(n1285), .Z(n1235) );
NOR2_X1 U997 ( .A1(n1100), .A2(n1286), .ZN(n1285) );
XOR2_X1 U998 ( .A(KEYINPUT59), .B(KEYINPUT25), .Z(n1286) );
XOR2_X1 U999 ( .A(G475), .B(KEYINPUT21), .Z(n1100) );
NOR2_X1 U1000 ( .A1(n1147), .A2(G902), .ZN(n1102) );
XNOR2_X1 U1001 ( .A(n1287), .B(n1288), .ZN(n1147) );
XOR2_X1 U1002 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1003 ( .A(n1264), .B(n1291), .ZN(n1290) );
NOR2_X1 U1004 ( .A1(KEYINPUT26), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1005 ( .A(KEYINPUT36), .B(G140), .Z(n1292) );
INV_X1 U1006 ( .A(G122), .ZN(n1264) );
XNOR2_X1 U1007 ( .A(n1119), .B(G125), .ZN(n1289) );
INV_X1 U1008 ( .A(G131), .ZN(n1119) );
XOR2_X1 U1009 ( .A(n1293), .B(n1267), .Z(n1287) );
XNOR2_X1 U1010 ( .A(G104), .B(n1245), .ZN(n1267) );
INV_X1 U1011 ( .A(G113), .ZN(n1245) );
XOR2_X1 U1012 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U1013 ( .A1(n1296), .A2(G214), .ZN(n1294) );
INV_X1 U1014 ( .A(n1077), .ZN(n1044) );
NAND2_X1 U1015 ( .A1(n1082), .A2(n1297), .ZN(n1077) );
NAND2_X1 U1016 ( .A1(n1079), .A2(n1080), .ZN(n1297) );
NAND3_X1 U1017 ( .A1(n1175), .A2(n1250), .A3(n1298), .ZN(n1080) );
INV_X1 U1018 ( .A(G469), .ZN(n1175) );
XNOR2_X1 U1019 ( .A(n1103), .B(KEYINPUT4), .ZN(n1079) );
NAND2_X1 U1020 ( .A1(G469), .A2(n1299), .ZN(n1103) );
NAND2_X1 U1021 ( .A1(n1298), .A2(n1250), .ZN(n1299) );
XNOR2_X1 U1022 ( .A(n1300), .B(n1171), .ZN(n1298) );
XNOR2_X1 U1023 ( .A(n1301), .B(n1302), .ZN(n1171) );
XNOR2_X1 U1024 ( .A(G140), .B(n1265), .ZN(n1302) );
XOR2_X1 U1025 ( .A(n1303), .B(n1304), .Z(n1301) );
NAND2_X1 U1026 ( .A1(G227), .A2(n1108), .ZN(n1303) );
NAND3_X1 U1027 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1300) );
OR2_X1 U1028 ( .A1(n1174), .A2(n1308), .ZN(n1307) );
NAND2_X1 U1029 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
INV_X1 U1030 ( .A(KEYINPUT45), .ZN(n1310) );
NAND2_X1 U1031 ( .A1(n1311), .A2(n1308), .ZN(n1309) );
XNOR2_X1 U1032 ( .A(n1174), .B(KEYINPUT23), .ZN(n1311) );
NAND2_X1 U1033 ( .A1(KEYINPUT45), .A2(n1312), .ZN(n1305) );
NAND2_X1 U1034 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
OR2_X1 U1035 ( .A1(n1174), .A2(KEYINPUT23), .ZN(n1314) );
NAND3_X1 U1036 ( .A1(n1174), .A2(n1308), .A3(KEYINPUT23), .ZN(n1313) );
XNOR2_X1 U1037 ( .A(n1116), .B(KEYINPUT1), .ZN(n1308) );
XOR2_X1 U1038 ( .A(G128), .B(n1315), .Z(n1116) );
NOR2_X1 U1039 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NOR2_X1 U1040 ( .A1(KEYINPUT39), .A2(n1295), .ZN(n1317) );
AND2_X1 U1041 ( .A1(KEYINPUT47), .A2(n1295), .ZN(n1316) );
XOR2_X1 U1042 ( .A(G101), .B(n1318), .Z(n1174) );
XOR2_X1 U1043 ( .A(G107), .B(G104), .Z(n1318) );
NAND2_X1 U1044 ( .A1(G221), .A2(n1319), .ZN(n1082) );
NOR2_X1 U1045 ( .A1(n1244), .A2(n1092), .ZN(n1069) );
XNOR2_X1 U1046 ( .A(n1320), .B(n1137), .ZN(n1092) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1319), .ZN(n1137) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1250), .ZN(n1319) );
OR2_X1 U1049 ( .A1(n1136), .A2(G902), .ZN(n1320) );
XNOR2_X1 U1050 ( .A(n1321), .B(n1322), .ZN(n1136) );
NOR2_X1 U1051 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1052 ( .A(n1325), .B(KEYINPUT33), .Z(n1324) );
NAND2_X1 U1053 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND3_X1 U1054 ( .A1(G234), .A2(n1108), .A3(G221), .ZN(n1327) );
AND4_X1 U1055 ( .A1(n1108), .A2(G234), .A3(G137), .A4(G221), .ZN(n1323) );
NAND2_X1 U1056 ( .A1(n1328), .A2(n1329), .ZN(n1321) );
NAND2_X1 U1057 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1058 ( .A(n1332), .B(n1117), .ZN(n1331) );
XOR2_X1 U1059 ( .A(n1333), .B(n1334), .Z(n1330) );
XOR2_X1 U1060 ( .A(n1335), .B(KEYINPUT18), .Z(n1328) );
NAND2_X1 U1061 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1062 ( .A(n1333), .B(n1334), .ZN(n1337) );
XOR2_X1 U1063 ( .A(G128), .B(n1338), .Z(n1334) );
NOR2_X1 U1064 ( .A1(G119), .A2(KEYINPUT14), .ZN(n1338) );
NAND2_X1 U1065 ( .A1(KEYINPUT10), .A2(n1265), .ZN(n1333) );
INV_X1 U1066 ( .A(G110), .ZN(n1265) );
XNOR2_X1 U1067 ( .A(G146), .B(n1117), .ZN(n1336) );
XOR2_X1 U1068 ( .A(G125), .B(G140), .Z(n1117) );
INV_X1 U1069 ( .A(n1236), .ZN(n1244) );
XOR2_X1 U1070 ( .A(n1339), .B(n1099), .Z(n1236) );
NAND2_X1 U1071 ( .A1(n1340), .A2(n1250), .ZN(n1099) );
INV_X1 U1072 ( .A(G902), .ZN(n1250) );
XOR2_X1 U1073 ( .A(n1341), .B(n1152), .Z(n1340) );
XNOR2_X1 U1074 ( .A(n1342), .B(G101), .ZN(n1152) );
NAND2_X1 U1075 ( .A1(n1296), .A2(G210), .ZN(n1342) );
AND2_X1 U1076 ( .A1(n1343), .A2(n1108), .ZN(n1296) );
INV_X1 U1077 ( .A(G953), .ZN(n1108) );
XNOR2_X1 U1078 ( .A(G237), .B(KEYINPUT12), .ZN(n1343) );
XOR2_X1 U1079 ( .A(n1160), .B(n1344), .Z(n1341) );
NOR2_X1 U1080 ( .A1(KEYINPUT49), .A2(n1345), .ZN(n1344) );
XNOR2_X1 U1081 ( .A(n1159), .B(KEYINPUT35), .ZN(n1345) );
XOR2_X1 U1082 ( .A(n1210), .B(n1304), .Z(n1159) );
XNOR2_X1 U1083 ( .A(n1346), .B(n1120), .ZN(n1304) );
XNOR2_X1 U1084 ( .A(G134), .B(n1326), .ZN(n1120) );
INV_X1 U1085 ( .A(G137), .ZN(n1326) );
XNOR2_X1 U1086 ( .A(G131), .B(KEYINPUT42), .ZN(n1346) );
XOR2_X1 U1087 ( .A(G128), .B(n1295), .Z(n1210) );
XNOR2_X1 U1088 ( .A(G143), .B(n1332), .ZN(n1295) );
INV_X1 U1089 ( .A(G146), .ZN(n1332) );
NAND2_X1 U1090 ( .A1(n1347), .A2(n1348), .ZN(n1160) );
NAND2_X1 U1091 ( .A1(G113), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1092 ( .A(n1350), .B(KEYINPUT51), .Z(n1347) );
OR2_X1 U1093 ( .A1(n1349), .A2(G113), .ZN(n1350) );
XNOR2_X1 U1094 ( .A(G116), .B(n1238), .ZN(n1349) );
INV_X1 U1095 ( .A(G119), .ZN(n1238) );
NAND2_X1 U1096 ( .A1(KEYINPUT56), .A2(n1155), .ZN(n1339) );
INV_X1 U1097 ( .A(G472), .ZN(n1155) );
endmodule


