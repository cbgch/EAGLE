//Key = 1101001101100111001101011010111000111011011110000101101001000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402;

XOR2_X1 U763 ( .A(G107), .B(n1063), .Z(G9) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(G75) );
NOR4_X1 U766 ( .A1(G953), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1067) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR3_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1078) );
NOR3_X1 U774 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1084) );
AND2_X1 U775 ( .A1(n1089), .A2(KEYINPUT4), .ZN(n1088) );
NOR3_X1 U776 ( .A1(KEYINPUT4), .A2(n1090), .A3(n1091), .ZN(n1087) );
NOR3_X1 U777 ( .A1(n1081), .A2(n1092), .A3(n1085), .ZN(n1073) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U779 ( .A1(n1095), .A2(n1077), .ZN(n1094) );
INV_X1 U780 ( .A(n1096), .ZN(n1077) );
NOR3_X1 U781 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1095) );
AND2_X1 U782 ( .A1(n1100), .A2(KEYINPUT33), .ZN(n1099) );
NOR3_X1 U783 ( .A1(KEYINPUT33), .A2(n1101), .A3(n1102), .ZN(n1098) );
NOR2_X1 U784 ( .A1(n1103), .A2(n1075), .ZN(n1093) );
NOR2_X1 U785 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR3_X1 U786 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1066) );
AND4_X1 U787 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1068) );
NOR4_X1 U788 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1109) );
AND2_X1 U789 ( .A1(n1114), .A2(G217), .ZN(n1113) );
XNOR2_X1 U790 ( .A(n1115), .B(n1116), .ZN(n1111) );
NOR2_X1 U791 ( .A1(G475), .A2(KEYINPUT20), .ZN(n1116) );
NAND3_X1 U792 ( .A1(n1091), .A2(n1117), .A3(n1118), .ZN(n1110) );
NOR3_X1 U793 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1108) );
AND2_X1 U794 ( .A1(n1122), .A2(KEYINPUT8), .ZN(n1121) );
NOR3_X1 U795 ( .A1(KEYINPUT8), .A2(n1123), .A3(n1122), .ZN(n1120) );
XNOR2_X1 U796 ( .A(KEYINPUT21), .B(n1124), .ZN(n1107) );
NOR2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(n1106) );
XNOR2_X1 U798 ( .A(n1127), .B(KEYINPUT29), .ZN(n1126) );
XOR2_X1 U799 ( .A(n1128), .B(KEYINPUT9), .Z(n1125) );
OR2_X1 U800 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U801 ( .A1(n1131), .A2(n1132), .ZN(G72) );
NAND2_X1 U802 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
INV_X1 U803 ( .A(n1135), .ZN(n1134) );
XOR2_X1 U804 ( .A(KEYINPUT37), .B(n1136), .Z(n1133) );
NAND2_X1 U805 ( .A1(n1137), .A2(n1135), .ZN(n1131) );
NAND2_X1 U806 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND2_X1 U807 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U808 ( .A(n1142), .B(n1143), .Z(n1140) );
NAND2_X1 U809 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
XOR2_X1 U810 ( .A(KEYINPUT53), .B(n1146), .Z(n1145) );
NAND3_X1 U811 ( .A1(n1143), .A2(G900), .A3(G953), .ZN(n1138) );
NOR2_X1 U812 ( .A1(KEYINPUT50), .A2(n1147), .ZN(n1143) );
XOR2_X1 U813 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U814 ( .A(n1150), .B(n1151), .ZN(n1149) );
XNOR2_X1 U815 ( .A(n1152), .B(n1153), .ZN(n1148) );
XOR2_X1 U816 ( .A(KEYINPUT10), .B(n1136), .Z(n1137) );
AND2_X1 U817 ( .A1(G953), .A2(n1154), .ZN(n1136) );
NAND2_X1 U818 ( .A1(G900), .A2(G227), .ZN(n1154) );
XOR2_X1 U819 ( .A(n1155), .B(n1156), .Z(G69) );
XOR2_X1 U820 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U821 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U822 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U823 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
XOR2_X1 U824 ( .A(KEYINPUT2), .B(n1165), .Z(n1164) );
NOR2_X1 U825 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U826 ( .A(n1168), .ZN(n1163) );
NOR2_X1 U827 ( .A1(KEYINPUT5), .A2(n1169), .ZN(n1157) );
NOR2_X1 U828 ( .A1(n1170), .A2(n1141), .ZN(n1169) );
AND2_X1 U829 ( .A1(G224), .A2(G898), .ZN(n1170) );
NAND3_X1 U830 ( .A1(n1171), .A2(n1141), .A3(KEYINPUT0), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1172), .A2(n1173), .ZN(G66) );
XOR2_X1 U832 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U833 ( .A(KEYINPUT34), .B(n1176), .Z(n1175) );
NOR2_X1 U834 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U835 ( .A1(n1172), .A2(n1179), .ZN(G63) );
XNOR2_X1 U836 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U837 ( .A1(n1182), .A2(n1178), .ZN(n1181) );
NOR2_X1 U838 ( .A1(n1172), .A2(n1183), .ZN(G60) );
NOR3_X1 U839 ( .A1(n1115), .A2(n1184), .A3(n1185), .ZN(n1183) );
NOR3_X1 U840 ( .A1(n1186), .A2(n1187), .A3(n1178), .ZN(n1185) );
NOR2_X1 U841 ( .A1(n1188), .A2(n1189), .ZN(n1184) );
AND2_X1 U842 ( .A1(n1070), .A2(G475), .ZN(n1189) );
XOR2_X1 U843 ( .A(n1190), .B(n1191), .Z(G6) );
XNOR2_X1 U844 ( .A(G104), .B(KEYINPUT46), .ZN(n1191) );
NAND3_X1 U845 ( .A1(n1192), .A2(n1193), .A3(n1105), .ZN(n1190) );
NOR2_X1 U846 ( .A1(n1172), .A2(n1194), .ZN(G57) );
XOR2_X1 U847 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U848 ( .A(n1197), .B(n1198), .ZN(n1196) );
XOR2_X1 U849 ( .A(n1199), .B(n1200), .Z(n1195) );
XOR2_X1 U850 ( .A(n1201), .B(n1202), .Z(n1200) );
NOR2_X1 U851 ( .A1(n1203), .A2(n1178), .ZN(n1202) );
NAND3_X1 U852 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1199) );
NAND2_X1 U853 ( .A1(G101), .A2(n1207), .ZN(n1206) );
OR3_X1 U854 ( .A1(n1207), .A2(G101), .A3(n1208), .ZN(n1205) );
INV_X1 U855 ( .A(KEYINPUT51), .ZN(n1207) );
NAND2_X1 U856 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
NAND2_X1 U857 ( .A1(n1210), .A2(KEYINPUT51), .ZN(n1209) );
XNOR2_X1 U858 ( .A(G101), .B(KEYINPUT22), .ZN(n1210) );
NOR2_X1 U859 ( .A1(n1172), .A2(n1211), .ZN(G54) );
XOR2_X1 U860 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U861 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U862 ( .A1(n1122), .A2(n1178), .ZN(n1215) );
XOR2_X1 U863 ( .A(n1216), .B(n1217), .Z(n1212) );
XOR2_X1 U864 ( .A(KEYINPUT24), .B(n1218), .Z(n1217) );
NOR2_X1 U865 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U866 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NOR2_X1 U867 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
AND2_X1 U868 ( .A1(G140), .A2(KEYINPUT41), .ZN(n1223) );
NOR2_X1 U869 ( .A1(G140), .A2(n1225), .ZN(n1219) );
NOR2_X1 U870 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U871 ( .A(KEYINPUT41), .ZN(n1227) );
NOR2_X1 U872 ( .A1(G110), .A2(n1224), .ZN(n1226) );
INV_X1 U873 ( .A(KEYINPUT28), .ZN(n1224) );
NAND2_X1 U874 ( .A1(KEYINPUT18), .A2(n1197), .ZN(n1216) );
NOR2_X1 U875 ( .A1(n1172), .A2(n1228), .ZN(G51) );
XOR2_X1 U876 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U877 ( .A(n1231), .B(n1232), .ZN(n1230) );
NOR2_X1 U878 ( .A1(n1129), .A2(n1178), .ZN(n1232) );
NAND2_X1 U879 ( .A1(G902), .A2(n1070), .ZN(n1178) );
NAND3_X1 U880 ( .A1(n1144), .A2(n1233), .A3(n1234), .ZN(n1070) );
INV_X1 U881 ( .A(n1171), .ZN(n1234) );
NAND4_X1 U882 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1171) );
AND4_X1 U883 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1238) );
AND2_X1 U884 ( .A1(n1243), .A2(n1244), .ZN(n1237) );
NAND3_X1 U885 ( .A1(n1245), .A2(n1105), .A3(n1246), .ZN(n1236) );
NOR3_X1 U886 ( .A1(n1085), .A2(n1247), .A3(n1248), .ZN(n1246) );
XNOR2_X1 U887 ( .A(n1249), .B(KEYINPUT19), .ZN(n1247) );
INV_X1 U888 ( .A(n1193), .ZN(n1085) );
XNOR2_X1 U889 ( .A(n1250), .B(KEYINPUT26), .ZN(n1245) );
NAND2_X1 U890 ( .A1(n1251), .A2(n1250), .ZN(n1235) );
XOR2_X1 U891 ( .A(n1065), .B(KEYINPUT38), .Z(n1251) );
NAND4_X1 U892 ( .A1(n1104), .A2(n1193), .A3(n1097), .A4(n1252), .ZN(n1065) );
XOR2_X1 U893 ( .A(KEYINPUT55), .B(n1146), .Z(n1233) );
AND4_X1 U894 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1146) );
AND3_X1 U895 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1144) );
NOR4_X1 U896 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1259) );
NOR2_X1 U897 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
INV_X1 U898 ( .A(KEYINPUT39), .ZN(n1264) );
NOR3_X1 U899 ( .A1(KEYINPUT39), .A2(n1266), .A3(n1081), .ZN(n1262) );
INV_X1 U900 ( .A(n1089), .ZN(n1081) );
AND2_X1 U901 ( .A1(KEYINPUT30), .A2(n1267), .ZN(n1261) );
NOR3_X1 U902 ( .A1(KEYINPUT30), .A2(n1086), .A3(n1268), .ZN(n1260) );
NAND2_X1 U903 ( .A1(n1269), .A2(n1270), .ZN(n1229) );
XOR2_X1 U904 ( .A(n1271), .B(KEYINPUT48), .Z(n1269) );
NOR2_X1 U905 ( .A1(n1141), .A2(G952), .ZN(n1172) );
XNOR2_X1 U906 ( .A(G146), .B(n1257), .ZN(G48) );
NAND3_X1 U907 ( .A1(n1105), .A2(n1086), .A3(n1272), .ZN(n1257) );
XOR2_X1 U908 ( .A(G143), .B(n1267), .Z(G45) );
NOR2_X1 U909 ( .A1(n1268), .A2(n1273), .ZN(n1267) );
NAND4_X1 U910 ( .A1(n1274), .A2(n1083), .A3(n1127), .A4(n1275), .ZN(n1268) );
XOR2_X1 U911 ( .A(n1265), .B(n1276), .Z(G42) );
NAND2_X1 U912 ( .A1(KEYINPUT13), .A2(G140), .ZN(n1276) );
NAND2_X1 U913 ( .A1(n1266), .A2(n1089), .ZN(n1265) );
AND3_X1 U914 ( .A1(n1105), .A2(n1082), .A3(n1274), .ZN(n1266) );
XNOR2_X1 U915 ( .A(G137), .B(n1258), .ZN(G39) );
NAND3_X1 U916 ( .A1(n1272), .A2(n1096), .A3(n1089), .ZN(n1258) );
XNOR2_X1 U917 ( .A(G134), .B(n1253), .ZN(G36) );
NAND2_X1 U918 ( .A1(n1277), .A2(n1104), .ZN(n1253) );
XNOR2_X1 U919 ( .A(G131), .B(n1254), .ZN(G33) );
NAND2_X1 U920 ( .A1(n1277), .A2(n1105), .ZN(n1254) );
INV_X1 U921 ( .A(n1278), .ZN(n1105) );
AND3_X1 U922 ( .A1(n1274), .A2(n1083), .A3(n1089), .ZN(n1277) );
NOR2_X1 U923 ( .A1(n1090), .A2(n1279), .ZN(n1089) );
INV_X1 U924 ( .A(n1091), .ZN(n1279) );
XNOR2_X1 U925 ( .A(G128), .B(n1255), .ZN(G30) );
NAND3_X1 U926 ( .A1(n1086), .A2(n1104), .A3(n1272), .ZN(n1255) );
AND3_X1 U927 ( .A1(n1119), .A2(n1280), .A3(n1274), .ZN(n1272) );
AND2_X1 U928 ( .A1(n1097), .A2(n1281), .ZN(n1274) );
INV_X1 U929 ( .A(n1248), .ZN(n1097) );
XOR2_X1 U930 ( .A(n1282), .B(G101), .Z(G3) );
NAND2_X1 U931 ( .A1(KEYINPUT63), .A2(n1244), .ZN(n1282) );
NAND3_X1 U932 ( .A1(n1096), .A2(n1192), .A3(n1083), .ZN(n1244) );
NAND2_X1 U933 ( .A1(n1283), .A2(n1284), .ZN(G27) );
OR2_X1 U934 ( .A1(n1256), .A2(G125), .ZN(n1284) );
XOR2_X1 U935 ( .A(n1285), .B(KEYINPUT58), .Z(n1283) );
NAND2_X1 U936 ( .A1(G125), .A2(n1256), .ZN(n1285) );
NAND4_X1 U937 ( .A1(n1086), .A2(n1281), .A3(n1082), .A4(n1286), .ZN(n1256) );
NOR2_X1 U938 ( .A1(n1278), .A2(n1075), .ZN(n1286) );
NAND2_X1 U939 ( .A1(n1287), .A2(n1288), .ZN(n1281) );
OR4_X1 U940 ( .A1(n1289), .A2(n1141), .A3(n1072), .A4(G900), .ZN(n1287) );
INV_X1 U941 ( .A(n1290), .ZN(n1072) );
XNOR2_X1 U942 ( .A(G122), .B(n1243), .ZN(G24) );
NAND4_X1 U943 ( .A1(n1291), .A2(n1193), .A3(n1127), .A4(n1275), .ZN(n1243) );
NOR2_X1 U944 ( .A1(n1280), .A2(n1119), .ZN(n1193) );
XNOR2_X1 U945 ( .A(G119), .B(n1242), .ZN(G21) );
NAND4_X1 U946 ( .A1(n1291), .A2(n1096), .A3(n1119), .A4(n1280), .ZN(n1242) );
XNOR2_X1 U947 ( .A(G116), .B(n1292), .ZN(G18) );
NAND2_X1 U948 ( .A1(KEYINPUT3), .A2(n1293), .ZN(n1292) );
INV_X1 U949 ( .A(n1241), .ZN(n1293) );
NAND3_X1 U950 ( .A1(n1083), .A2(n1104), .A3(n1291), .ZN(n1241) );
NOR3_X1 U951 ( .A1(n1273), .A2(n1249), .A3(n1075), .ZN(n1291) );
INV_X1 U952 ( .A(n1100), .ZN(n1075) );
NOR2_X1 U953 ( .A1(n1275), .A2(n1294), .ZN(n1104) );
INV_X1 U954 ( .A(n1127), .ZN(n1294) );
XNOR2_X1 U955 ( .A(G113), .B(n1240), .ZN(G15) );
NAND3_X1 U956 ( .A1(n1083), .A2(n1100), .A3(n1295), .ZN(n1240) );
NOR3_X1 U957 ( .A1(n1278), .A2(n1249), .A3(n1064), .ZN(n1295) );
NAND2_X1 U958 ( .A1(n1296), .A2(n1275), .ZN(n1278) );
XNOR2_X1 U959 ( .A(KEYINPUT40), .B(n1297), .ZN(n1296) );
NOR2_X1 U960 ( .A1(n1101), .A2(n1112), .ZN(n1100) );
INV_X1 U961 ( .A(n1102), .ZN(n1112) );
AND2_X1 U962 ( .A1(n1298), .A2(n1119), .ZN(n1083) );
XNOR2_X1 U963 ( .A(G110), .B(n1239), .ZN(G12) );
NAND3_X1 U964 ( .A1(n1096), .A2(n1192), .A3(n1082), .ZN(n1239) );
NOR2_X1 U965 ( .A1(n1119), .A2(n1298), .ZN(n1082) );
INV_X1 U966 ( .A(n1280), .ZN(n1298) );
NAND2_X1 U967 ( .A1(n1124), .A2(n1299), .ZN(n1280) );
NAND2_X1 U968 ( .A1(G217), .A2(n1114), .ZN(n1299) );
NAND2_X1 U969 ( .A1(n1289), .A2(n1300), .ZN(n1114) );
OR2_X1 U970 ( .A1(n1174), .A2(G234), .ZN(n1300) );
NAND3_X1 U971 ( .A1(n1301), .A2(n1289), .A3(n1174), .ZN(n1124) );
XNOR2_X1 U972 ( .A(n1302), .B(n1303), .ZN(n1174) );
XOR2_X1 U973 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U974 ( .A(n1306), .B(n1307), .Z(n1305) );
AND3_X1 U975 ( .A1(G221), .A2(n1308), .A3(G234), .ZN(n1307) );
NAND2_X1 U976 ( .A1(KEYINPUT52), .A2(n1309), .ZN(n1306) );
NAND2_X1 U977 ( .A1(KEYINPUT14), .A2(G128), .ZN(n1304) );
XNOR2_X1 U978 ( .A(G110), .B(n1310), .ZN(n1302) );
XOR2_X1 U979 ( .A(G137), .B(G119), .Z(n1310) );
OR2_X1 U980 ( .A1(n1177), .A2(G234), .ZN(n1301) );
INV_X1 U981 ( .A(G217), .ZN(n1177) );
XOR2_X1 U982 ( .A(n1311), .B(n1203), .Z(n1119) );
INV_X1 U983 ( .A(G472), .ZN(n1203) );
NAND2_X1 U984 ( .A1(n1312), .A2(n1289), .ZN(n1311) );
XOR2_X1 U985 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U986 ( .A(n1208), .B(G101), .ZN(n1314) );
AND3_X1 U987 ( .A1(n1308), .A2(n1315), .A3(G210), .ZN(n1208) );
NAND2_X1 U988 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND2_X1 U989 ( .A1(n1318), .A2(n1198), .ZN(n1317) );
XOR2_X1 U990 ( .A(KEYINPUT49), .B(n1319), .Z(n1316) );
NOR2_X1 U991 ( .A1(n1318), .A2(n1198), .ZN(n1319) );
XOR2_X1 U992 ( .A(n1320), .B(n1321), .Z(n1198) );
NOR2_X1 U993 ( .A1(G113), .A2(KEYINPUT12), .ZN(n1321) );
XNOR2_X1 U994 ( .A(n1322), .B(n1197), .ZN(n1318) );
XNOR2_X1 U995 ( .A(KEYINPUT17), .B(n1323), .ZN(n1322) );
NOR2_X1 U996 ( .A1(KEYINPUT31), .A2(n1201), .ZN(n1323) );
NOR3_X1 U997 ( .A1(n1064), .A2(n1249), .A3(n1248), .ZN(n1192) );
NAND2_X1 U998 ( .A1(n1102), .A2(n1101), .ZN(n1248) );
NAND2_X1 U999 ( .A1(n1324), .A2(n1117), .ZN(n1101) );
NAND2_X1 U1000 ( .A1(n1123), .A2(n1122), .ZN(n1117) );
INV_X1 U1001 ( .A(G469), .ZN(n1122) );
INV_X1 U1002 ( .A(n1325), .ZN(n1123) );
NAND2_X1 U1003 ( .A1(G469), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1004 ( .A1(n1326), .A2(n1289), .ZN(n1325) );
XOR2_X1 U1005 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1006 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1007 ( .A(KEYINPUT35), .B(KEYINPUT1), .Z(n1330) );
NOR2_X1 U1008 ( .A1(KEYINPUT60), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1009 ( .A(n1222), .B(n1332), .ZN(n1331) );
XOR2_X1 U1010 ( .A(KEYINPUT62), .B(G140), .Z(n1332) );
INV_X1 U1011 ( .A(G110), .ZN(n1222) );
XNOR2_X1 U1012 ( .A(n1214), .B(n1197), .ZN(n1327) );
XOR2_X1 U1013 ( .A(n1333), .B(n1150), .Z(n1197) );
XOR2_X1 U1014 ( .A(G134), .B(G137), .Z(n1150) );
NAND2_X1 U1015 ( .A1(KEYINPUT43), .A2(n1153), .ZN(n1333) );
XOR2_X1 U1016 ( .A(n1334), .B(n1335), .Z(n1214) );
XNOR2_X1 U1017 ( .A(n1336), .B(n1166), .ZN(n1335) );
AND2_X1 U1018 ( .A1(n1308), .A2(G227), .ZN(n1336) );
XOR2_X1 U1019 ( .A(n1152), .B(KEYINPUT11), .Z(n1334) );
NAND2_X1 U1020 ( .A1(n1337), .A2(n1338), .ZN(n1152) );
NAND2_X1 U1021 ( .A1(G128), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1022 ( .A(KEYINPUT57), .B(n1340), .Z(n1337) );
NOR2_X1 U1023 ( .A1(G128), .A2(n1339), .ZN(n1340) );
NAND2_X1 U1024 ( .A1(G221), .A2(n1341), .ZN(n1102) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1289), .ZN(n1341) );
INV_X1 U1026 ( .A(n1252), .ZN(n1249) );
NAND2_X1 U1027 ( .A1(n1288), .A2(n1342), .ZN(n1252) );
NAND3_X1 U1028 ( .A1(n1159), .A2(n1290), .A3(G902), .ZN(n1342) );
NOR2_X1 U1029 ( .A1(n1141), .A2(G898), .ZN(n1159) );
INV_X1 U1030 ( .A(G953), .ZN(n1141) );
NAND3_X1 U1031 ( .A1(G952), .A2(n1290), .A3(n1343), .ZN(n1288) );
XNOR2_X1 U1032 ( .A(G953), .B(KEYINPUT16), .ZN(n1343) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1290) );
INV_X1 U1034 ( .A(n1250), .ZN(n1064) );
XOR2_X1 U1035 ( .A(n1086), .B(KEYINPUT59), .Z(n1250) );
INV_X1 U1036 ( .A(n1273), .ZN(n1086) );
NAND2_X1 U1037 ( .A1(n1091), .A2(n1090), .ZN(n1273) );
NAND3_X1 U1038 ( .A1(n1344), .A2(n1345), .A3(n1118), .ZN(n1090) );
NAND2_X1 U1039 ( .A1(n1130), .A2(n1129), .ZN(n1118) );
NAND2_X1 U1040 ( .A1(KEYINPUT27), .A2(n1129), .ZN(n1345) );
OR3_X1 U1041 ( .A1(n1130), .A2(KEYINPUT27), .A3(n1129), .ZN(n1344) );
NAND2_X1 U1042 ( .A1(G210), .A2(n1346), .ZN(n1129) );
AND2_X1 U1043 ( .A1(n1347), .A2(n1289), .ZN(n1130) );
XOR2_X1 U1044 ( .A(n1231), .B(n1348), .Z(n1347) );
NAND2_X1 U1045 ( .A1(n1270), .A2(n1271), .ZN(n1348) );
NAND2_X1 U1046 ( .A1(n1349), .A2(n1350), .ZN(n1271) );
NAND2_X1 U1047 ( .A1(G224), .A2(n1308), .ZN(n1350) );
XOR2_X1 U1048 ( .A(n1201), .B(G125), .Z(n1349) );
NAND3_X1 U1049 ( .A1(n1351), .A2(n1308), .A3(G224), .ZN(n1270) );
XNOR2_X1 U1050 ( .A(G125), .B(n1201), .ZN(n1351) );
NAND3_X1 U1051 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1201) );
NAND2_X1 U1052 ( .A1(KEYINPUT47), .A2(n1355), .ZN(n1354) );
INV_X1 U1053 ( .A(n1339), .ZN(n1355) );
OR3_X1 U1054 ( .A1(n1356), .A2(KEYINPUT47), .A3(G128), .ZN(n1353) );
NAND2_X1 U1055 ( .A1(G128), .A2(n1356), .ZN(n1352) );
NAND2_X1 U1056 ( .A1(KEYINPUT7), .A2(n1339), .ZN(n1356) );
XOR2_X1 U1057 ( .A(G146), .B(G143), .Z(n1339) );
NAND2_X1 U1058 ( .A1(n1357), .A2(n1358), .ZN(n1231) );
NAND2_X1 U1059 ( .A1(n1162), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1060 ( .A(KEYINPUT23), .B(n1360), .Z(n1357) );
NOR2_X1 U1061 ( .A1(n1162), .A2(n1359), .ZN(n1360) );
NAND2_X1 U1062 ( .A1(n1361), .A2(n1362), .ZN(n1359) );
NAND2_X1 U1063 ( .A1(KEYINPUT61), .A2(n1363), .ZN(n1362) );
NAND2_X1 U1064 ( .A1(n1168), .A2(n1364), .ZN(n1363) );
OR2_X1 U1065 ( .A1(n1167), .A2(n1166), .ZN(n1364) );
NAND2_X1 U1066 ( .A1(n1166), .A2(n1167), .ZN(n1168) );
NAND2_X1 U1067 ( .A1(n1365), .A2(n1366), .ZN(n1361) );
INV_X1 U1068 ( .A(KEYINPUT61), .ZN(n1366) );
XOR2_X1 U1069 ( .A(n1167), .B(n1166), .Z(n1365) );
XOR2_X1 U1070 ( .A(n1367), .B(n1368), .Z(n1166) );
XOR2_X1 U1071 ( .A(KEYINPUT32), .B(G107), .Z(n1368) );
XNOR2_X1 U1072 ( .A(G104), .B(G101), .ZN(n1367) );
NAND2_X1 U1073 ( .A1(n1369), .A2(n1370), .ZN(n1167) );
NAND2_X1 U1074 ( .A1(G113), .A2(n1320), .ZN(n1370) );
XOR2_X1 U1075 ( .A(KEYINPUT6), .B(n1371), .Z(n1369) );
NOR2_X1 U1076 ( .A1(G113), .A2(n1320), .ZN(n1371) );
XOR2_X1 U1077 ( .A(G116), .B(G119), .Z(n1320) );
XNOR2_X1 U1078 ( .A(G122), .B(G110), .ZN(n1162) );
NAND2_X1 U1079 ( .A1(G214), .A2(n1346), .ZN(n1091) );
NAND2_X1 U1080 ( .A1(n1315), .A2(n1289), .ZN(n1346) );
NOR2_X1 U1081 ( .A1(n1275), .A2(n1297), .ZN(n1096) );
XNOR2_X1 U1082 ( .A(n1127), .B(KEYINPUT36), .ZN(n1297) );
XOR2_X1 U1083 ( .A(n1372), .B(n1182), .Z(n1127) );
INV_X1 U1084 ( .A(G478), .ZN(n1182) );
NAND2_X1 U1085 ( .A1(n1180), .A2(n1289), .ZN(n1372) );
INV_X1 U1086 ( .A(G902), .ZN(n1289) );
XNOR2_X1 U1087 ( .A(n1373), .B(n1374), .ZN(n1180) );
XOR2_X1 U1088 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1089 ( .A(G128), .B(G122), .Z(n1376) );
XOR2_X1 U1090 ( .A(G143), .B(G134), .Z(n1375) );
XOR2_X1 U1091 ( .A(n1377), .B(n1378), .Z(n1373) );
XOR2_X1 U1092 ( .A(G116), .B(G107), .Z(n1378) );
NAND3_X1 U1093 ( .A1(G217), .A2(n1308), .A3(G234), .ZN(n1377) );
NAND3_X1 U1094 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1275) );
OR2_X1 U1095 ( .A1(n1382), .A2(KEYINPUT42), .ZN(n1381) );
NAND3_X1 U1096 ( .A1(KEYINPUT42), .A2(n1382), .A3(G475), .ZN(n1380) );
INV_X1 U1097 ( .A(n1115), .ZN(n1382) );
NAND2_X1 U1098 ( .A1(n1383), .A2(n1187), .ZN(n1379) );
INV_X1 U1099 ( .A(G475), .ZN(n1187) );
NAND2_X1 U1100 ( .A1(n1384), .A2(KEYINPUT42), .ZN(n1383) );
XNOR2_X1 U1101 ( .A(n1115), .B(KEYINPUT45), .ZN(n1384) );
NOR2_X1 U1102 ( .A1(n1188), .A2(G902), .ZN(n1115) );
INV_X1 U1103 ( .A(n1186), .ZN(n1188) );
NAND2_X1 U1104 ( .A1(n1385), .A2(n1386), .ZN(n1186) );
NAND2_X1 U1105 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1389), .Z(n1385) );
NOR2_X1 U1107 ( .A1(n1387), .A2(n1388), .ZN(n1389) );
NAND2_X1 U1108 ( .A1(n1390), .A2(n1391), .ZN(n1388) );
NAND2_X1 U1109 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
XOR2_X1 U1110 ( .A(n1394), .B(n1395), .Z(n1393) );
XNOR2_X1 U1111 ( .A(n1309), .B(KEYINPUT56), .ZN(n1392) );
XOR2_X1 U1112 ( .A(n1396), .B(KEYINPUT25), .Z(n1390) );
NAND2_X1 U1113 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
XNOR2_X1 U1114 ( .A(KEYINPUT56), .B(n1399), .ZN(n1398) );
INV_X1 U1115 ( .A(n1309), .ZN(n1399) );
XOR2_X1 U1116 ( .A(G146), .B(n1151), .Z(n1309) );
XOR2_X1 U1117 ( .A(G125), .B(G140), .Z(n1151) );
XNOR2_X1 U1118 ( .A(n1395), .B(n1394), .ZN(n1397) );
NAND2_X1 U1119 ( .A1(KEYINPUT44), .A2(n1153), .ZN(n1394) );
INV_X1 U1120 ( .A(G131), .ZN(n1153) );
XOR2_X1 U1121 ( .A(n1400), .B(G143), .Z(n1395) );
NAND3_X1 U1122 ( .A1(n1308), .A2(n1315), .A3(G214), .ZN(n1400) );
INV_X1 U1123 ( .A(G237), .ZN(n1315) );
XOR2_X1 U1124 ( .A(G953), .B(KEYINPUT15), .Z(n1308) );
XNOR2_X1 U1125 ( .A(n1401), .B(n1402), .ZN(n1387) );
XOR2_X1 U1126 ( .A(G122), .B(G113), .Z(n1402) );
INV_X1 U1127 ( .A(G104), .ZN(n1401) );
endmodule


