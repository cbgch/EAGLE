//Key = 1101011111100110010000111001101111100101101001100010011010101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370;

XOR2_X1 U749 ( .A(G107), .B(n1029), .Z(G9) );
NOR2_X1 U750 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U751 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR4_X1 U752 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1034) );
NOR2_X1 U753 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NOR2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1036) );
AND2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1042) );
NOR3_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NOR2_X1 U758 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U759 ( .A(KEYINPUT31), .B(n1053), .ZN(n1052) );
NOR3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1049) );
NOR2_X1 U761 ( .A1(n1053), .A2(n1057), .ZN(n1048) );
NAND4_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1032) );
NAND4_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1044), .A4(n1054), .ZN(n1059) );
INV_X1 U764 ( .A(KEYINPUT27), .ZN(n1054) );
NAND4_X1 U765 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1041), .ZN(n1044) );
NAND2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
NAND2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1058) );
XOR2_X1 U771 ( .A(KEYINPUT51), .B(n1040), .Z(n1076) );
AND2_X1 U772 ( .A1(n1062), .A2(n1067), .ZN(n1040) );
NOR3_X1 U773 ( .A1(n1047), .A2(n1055), .A3(n1039), .ZN(n1062) );
NOR3_X1 U774 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U775 ( .A(n1060), .ZN(n1077) );
NAND4_X1 U776 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1060) );
NOR3_X1 U777 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
INV_X1 U778 ( .A(n1085), .ZN(n1084) );
NOR3_X1 U779 ( .A1(n1071), .A2(n1086), .A3(n1087), .ZN(n1080) );
NOR3_X1 U780 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1079) );
AND2_X1 U781 ( .A1(n1091), .A2(G478), .ZN(n1090) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1089) );
XOR2_X1 U783 ( .A(n1094), .B(KEYINPUT26), .Z(n1093) );
NOR2_X1 U784 ( .A1(G472), .A2(n1095), .ZN(n1088) );
NOR3_X1 U785 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1078) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(n1098) );
XNOR2_X1 U787 ( .A(KEYINPUT6), .B(n1101), .ZN(n1100) );
NAND2_X1 U788 ( .A1(KEYINPUT22), .A2(G475), .ZN(n1099) );
XOR2_X1 U789 ( .A(n1102), .B(KEYINPUT54), .Z(n1097) );
NAND2_X1 U790 ( .A1(G472), .A2(n1095), .ZN(n1102) );
XNOR2_X1 U791 ( .A(n1103), .B(n1104), .ZN(n1096) );
NOR2_X1 U792 ( .A1(KEYINPUT59), .A2(n1105), .ZN(n1104) );
INV_X1 U793 ( .A(n1106), .ZN(n1105) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(G72) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1061), .ZN(n1108) );
AND2_X1 U796 ( .A1(G227), .A2(G900), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NAND2_X1 U798 ( .A1(n1112), .A2(n1061), .ZN(n1111) );
XNOR2_X1 U799 ( .A(n1035), .B(n1113), .ZN(n1112) );
OR3_X1 U800 ( .A1(n1114), .A2(n1113), .A3(n1061), .ZN(n1110) );
XNOR2_X1 U801 ( .A(n1115), .B(n1116), .ZN(n1113) );
XNOR2_X1 U802 ( .A(KEYINPUT16), .B(n1117), .ZN(n1116) );
XOR2_X1 U803 ( .A(n1118), .B(n1119), .Z(n1115) );
NOR2_X1 U804 ( .A1(KEYINPUT52), .A2(n1120), .ZN(n1119) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U806 ( .A1(KEYINPUT12), .A2(G131), .ZN(n1122) );
XNOR2_X1 U807 ( .A(G134), .B(G137), .ZN(n1121) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(G69) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U810 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U811 ( .A(n1129), .B(n1130), .Z(n1127) );
NAND2_X1 U812 ( .A1(KEYINPUT45), .A2(n1131), .ZN(n1129) );
NAND2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1123) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U815 ( .A1(G953), .A2(n1136), .ZN(n1135) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1136) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U819 ( .A1(G953), .A2(n1141), .ZN(n1140) );
INV_X1 U820 ( .A(n1125), .ZN(n1139) );
INV_X1 U821 ( .A(n1134), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1142), .A2(n1143), .ZN(n1134) );
NAND2_X1 U823 ( .A1(KEYINPUT13), .A2(n1144), .ZN(n1143) );
OR2_X1 U824 ( .A1(KEYINPUT17), .A2(n1144), .ZN(n1142) );
AND2_X1 U825 ( .A1(n1061), .A2(n1033), .ZN(n1144) );
NOR2_X1 U826 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U828 ( .A1(n1103), .A2(n1149), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1150), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1151), .B(n1152), .ZN(n1150) );
AND2_X1 U831 ( .A1(G478), .A2(n1153), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1145), .A2(n1154), .ZN(G60) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
AND2_X1 U834 ( .A1(G475), .A2(n1153), .ZN(n1156) );
NAND2_X1 U835 ( .A1(KEYINPUT40), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U836 ( .A(G104), .B(n1158), .ZN(G6) );
NAND3_X1 U837 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
NOR3_X1 U838 ( .A1(n1053), .A2(n1162), .A3(n1069), .ZN(n1161) );
XNOR2_X1 U839 ( .A(n1075), .B(KEYINPUT34), .ZN(n1159) );
NOR2_X1 U840 ( .A1(n1145), .A2(n1163), .ZN(G57) );
XOR2_X1 U841 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U842 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U843 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND3_X1 U844 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
NAND2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U846 ( .A1(KEYINPUT48), .A2(n1175), .ZN(n1171) );
NAND2_X1 U847 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XNOR2_X1 U848 ( .A(KEYINPUT37), .B(n1178), .ZN(n1176) );
NAND2_X1 U849 ( .A1(n1179), .A2(n1180), .ZN(n1170) );
INV_X1 U850 ( .A(KEYINPUT48), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NAND3_X1 U852 ( .A1(KEYINPUT37), .A2(n1177), .A3(n1178), .ZN(n1182) );
OR2_X1 U853 ( .A1(n1178), .A2(KEYINPUT37), .ZN(n1181) );
INV_X1 U854 ( .A(n1174), .ZN(n1178) );
NOR2_X1 U855 ( .A1(G101), .A2(KEYINPUT44), .ZN(n1166) );
XOR2_X1 U856 ( .A(n1183), .B(n1184), .Z(n1164) );
AND2_X1 U857 ( .A1(G472), .A2(n1153), .ZN(n1184) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(G54) );
XOR2_X1 U859 ( .A(n1118), .B(n1187), .Z(n1186) );
XOR2_X1 U860 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U861 ( .A1(KEYINPUT56), .A2(n1190), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1153), .A2(G469), .ZN(n1190) );
INV_X1 U863 ( .A(n1149), .ZN(n1153) );
XNOR2_X1 U864 ( .A(G140), .B(n1191), .ZN(n1118) );
NOR2_X1 U865 ( .A1(n1192), .A2(n1193), .ZN(n1185) );
XOR2_X1 U866 ( .A(KEYINPUT8), .B(n1194), .Z(n1193) );
XNOR2_X1 U867 ( .A(KEYINPUT25), .B(G953), .ZN(n1192) );
NOR2_X1 U868 ( .A1(n1145), .A2(n1195), .ZN(G51) );
XOR2_X1 U869 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U870 ( .A1(n1094), .A2(n1149), .ZN(n1197) );
NAND2_X1 U871 ( .A1(G902), .A2(n1198), .ZN(n1149) );
OR2_X1 U872 ( .A1(n1033), .A2(n1035), .ZN(n1198) );
NAND4_X1 U873 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1035) );
NOR4_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR2_X1 U875 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U876 ( .A(n1209), .B(KEYINPUT20), .Z(n1207) );
NOR3_X1 U877 ( .A1(n1210), .A2(n1055), .A3(n1211), .ZN(n1205) );
NOR4_X1 U878 ( .A1(n1212), .A2(n1213), .A3(n1056), .A4(n1214), .ZN(n1204) );
NOR2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1201) );
NAND4_X1 U880 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1033) );
NOR4_X1 U881 ( .A1(n1029), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1220) );
NOR4_X1 U882 ( .A1(n1057), .A2(n1053), .A3(n1213), .A4(n1162), .ZN(n1029) );
NAND2_X1 U883 ( .A1(n1067), .A2(n1224), .ZN(n1219) );
NAND2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND3_X1 U885 ( .A1(n1227), .A2(n1228), .A3(n1160), .ZN(n1226) );
NAND2_X1 U886 ( .A1(n1229), .A2(n1230), .ZN(n1225) );
NAND2_X1 U887 ( .A1(KEYINPUT39), .A2(n1231), .ZN(n1196) );
AND2_X1 U888 ( .A1(n1232), .A2(n1194), .ZN(n1145) );
XOR2_X1 U889 ( .A(G952), .B(KEYINPUT62), .Z(n1194) );
XNOR2_X1 U890 ( .A(KEYINPUT25), .B(n1061), .ZN(n1232) );
XOR2_X1 U891 ( .A(G146), .B(n1233), .Z(G48) );
NOR2_X1 U892 ( .A1(n1208), .A2(n1209), .ZN(n1233) );
NAND4_X1 U893 ( .A1(n1234), .A2(n1160), .A3(n1235), .A4(n1236), .ZN(n1209) );
XOR2_X1 U894 ( .A(n1237), .B(n1238), .Z(G45) );
NAND2_X1 U895 ( .A1(KEYINPUT23), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U896 ( .A(KEYINPUT36), .B(n1240), .ZN(n1239) );
NAND4_X1 U897 ( .A1(n1241), .A2(n1229), .A3(n1227), .A4(n1236), .ZN(n1237) );
INV_X1 U898 ( .A(n1214), .ZN(n1229) );
XNOR2_X1 U899 ( .A(n1063), .B(KEYINPUT9), .ZN(n1241) );
XNOR2_X1 U900 ( .A(n1242), .B(n1216), .ZN(G42) );
NOR3_X1 U901 ( .A1(n1051), .A2(n1243), .A3(n1210), .ZN(n1216) );
INV_X1 U902 ( .A(n1074), .ZN(n1243) );
XOR2_X1 U903 ( .A(n1244), .B(n1245), .Z(G39) );
XNOR2_X1 U904 ( .A(KEYINPUT35), .B(n1246), .ZN(n1245) );
NOR3_X1 U905 ( .A1(n1247), .A2(n1211), .A3(n1210), .ZN(n1244) );
XNOR2_X1 U906 ( .A(KEYINPUT50), .B(n1055), .ZN(n1247) );
XNOR2_X1 U907 ( .A(n1248), .B(n1249), .ZN(G36) );
NAND2_X1 U908 ( .A1(KEYINPUT7), .A2(n1250), .ZN(n1248) );
INV_X1 U909 ( .A(n1203), .ZN(n1250) );
NOR3_X1 U910 ( .A1(n1056), .A2(n1057), .A3(n1210), .ZN(n1203) );
XOR2_X1 U911 ( .A(n1251), .B(n1215), .Z(G33) );
NOR3_X1 U912 ( .A1(n1056), .A2(n1051), .A3(n1210), .ZN(n1215) );
NAND4_X1 U913 ( .A1(n1064), .A2(n1235), .A3(n1236), .A4(n1041), .ZN(n1210) );
NAND2_X1 U914 ( .A1(KEYINPUT3), .A2(n1252), .ZN(n1251) );
INV_X1 U915 ( .A(G131), .ZN(n1252) );
XNOR2_X1 U916 ( .A(n1199), .B(n1253), .ZN(G30) );
NOR2_X1 U917 ( .A1(KEYINPUT15), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U918 ( .A(G128), .B(KEYINPUT18), .ZN(n1254) );
OR4_X1 U919 ( .A1(n1211), .A2(n1057), .A3(n1213), .A4(n1212), .ZN(n1199) );
XNOR2_X1 U920 ( .A(G101), .B(n1217), .ZN(G3) );
NAND2_X1 U921 ( .A1(n1063), .A2(n1255), .ZN(n1217) );
INV_X1 U922 ( .A(n1056), .ZN(n1063) );
XNOR2_X1 U923 ( .A(G125), .B(n1200), .ZN(G27) );
NAND4_X1 U924 ( .A1(n1160), .A2(n1073), .A3(n1256), .A4(n1074), .ZN(n1200) );
NOR2_X1 U925 ( .A1(n1212), .A2(n1208), .ZN(n1256) );
INV_X1 U926 ( .A(n1236), .ZN(n1212) );
NAND2_X1 U927 ( .A1(n1039), .A2(n1257), .ZN(n1236) );
NAND4_X1 U928 ( .A1(G902), .A2(G953), .A3(n1258), .A4(n1114), .ZN(n1257) );
INV_X1 U929 ( .A(G900), .ZN(n1114) );
INV_X1 U930 ( .A(n1047), .ZN(n1073) );
INV_X1 U931 ( .A(n1051), .ZN(n1160) );
XOR2_X1 U932 ( .A(G122), .B(n1259), .Z(G24) );
NOR4_X1 U933 ( .A1(KEYINPUT41), .A2(n1053), .A3(n1260), .A4(n1214), .ZN(n1259) );
NAND2_X1 U934 ( .A1(n1261), .A2(n1262), .ZN(n1214) );
INV_X1 U935 ( .A(n1067), .ZN(n1053) );
NOR2_X1 U936 ( .A1(n1263), .A2(n1264), .ZN(n1067) );
XNOR2_X1 U937 ( .A(G119), .B(n1218), .ZN(G21) );
NAND3_X1 U938 ( .A1(n1230), .A2(n1045), .A3(n1234), .ZN(n1218) );
INV_X1 U939 ( .A(n1211), .ZN(n1234) );
NAND2_X1 U940 ( .A1(n1264), .A2(n1263), .ZN(n1211) );
INV_X1 U941 ( .A(n1265), .ZN(n1264) );
XNOR2_X1 U942 ( .A(n1266), .B(n1223), .ZN(G18) );
NOR3_X1 U943 ( .A1(n1260), .A2(n1057), .A3(n1056), .ZN(n1223) );
OR2_X1 U944 ( .A1(n1261), .A2(n1267), .ZN(n1057) );
XNOR2_X1 U945 ( .A(n1268), .B(n1222), .ZN(G15) );
NOR3_X1 U946 ( .A1(n1051), .A2(n1260), .A3(n1056), .ZN(n1222) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1263), .ZN(n1056) );
INV_X1 U948 ( .A(n1230), .ZN(n1260) );
NOR3_X1 U949 ( .A1(n1208), .A2(n1162), .A3(n1047), .ZN(n1230) );
NAND2_X1 U950 ( .A1(n1072), .A2(n1269), .ZN(n1047) );
NAND2_X1 U951 ( .A1(n1267), .A2(n1261), .ZN(n1051) );
INV_X1 U952 ( .A(n1262), .ZN(n1267) );
NAND2_X1 U953 ( .A1(n1270), .A2(n1271), .ZN(G12) );
NAND2_X1 U954 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U955 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
NAND2_X1 U956 ( .A1(KEYINPUT5), .A2(n1276), .ZN(n1275) );
INV_X1 U957 ( .A(KEYINPUT60), .ZN(n1276) );
NAND3_X1 U958 ( .A1(n1277), .A2(n1278), .A3(KEYINPUT60), .ZN(n1270) );
OR2_X1 U959 ( .A1(G110), .A2(KEYINPUT5), .ZN(n1278) );
NAND2_X1 U960 ( .A1(KEYINPUT5), .A2(n1279), .ZN(n1277) );
NAND2_X1 U961 ( .A1(n1221), .A2(n1274), .ZN(n1279) );
INV_X1 U962 ( .A(n1273), .ZN(n1221) );
NAND2_X1 U963 ( .A1(n1074), .A2(n1255), .ZN(n1273) );
NOR3_X1 U964 ( .A1(n1213), .A2(n1162), .A3(n1055), .ZN(n1255) );
INV_X1 U965 ( .A(n1045), .ZN(n1055) );
NOR2_X1 U966 ( .A1(n1262), .A2(n1261), .ZN(n1045) );
XNOR2_X1 U967 ( .A(n1101), .B(G475), .ZN(n1261) );
NAND2_X1 U968 ( .A1(n1157), .A2(n1280), .ZN(n1101) );
XNOR2_X1 U969 ( .A(n1281), .B(n1282), .ZN(n1157) );
XOR2_X1 U970 ( .A(n1283), .B(n1284), .Z(n1282) );
AND3_X1 U971 ( .A1(G214), .A2(n1061), .A3(n1285), .ZN(n1284) );
NOR2_X1 U972 ( .A1(KEYINPUT21), .A2(G131), .ZN(n1283) );
XOR2_X1 U973 ( .A(n1286), .B(n1287), .Z(n1281) );
AND2_X1 U974 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U975 ( .A(n1290), .B(n1291), .Z(n1286) );
XNOR2_X1 U976 ( .A(n1268), .B(n1292), .ZN(n1291) );
XNOR2_X1 U977 ( .A(KEYINPUT10), .B(n1240), .ZN(n1292) );
XOR2_X1 U978 ( .A(n1293), .B(n1294), .Z(n1290) );
XNOR2_X1 U979 ( .A(G104), .B(n1295), .ZN(n1293) );
NAND2_X1 U980 ( .A1(n1296), .A2(n1297), .ZN(n1262) );
NAND2_X1 U981 ( .A1(G478), .A2(n1091), .ZN(n1297) );
XOR2_X1 U982 ( .A(KEYINPUT14), .B(n1083), .Z(n1296) );
NOR2_X1 U983 ( .A1(n1091), .A2(G478), .ZN(n1083) );
NAND2_X1 U984 ( .A1(n1151), .A2(n1280), .ZN(n1091) );
XNOR2_X1 U985 ( .A(n1298), .B(n1299), .ZN(n1151) );
XNOR2_X1 U986 ( .A(n1300), .B(n1301), .ZN(n1299) );
XNOR2_X1 U987 ( .A(n1240), .B(G134), .ZN(n1301) );
XOR2_X1 U988 ( .A(n1302), .B(n1303), .Z(n1298) );
AND2_X1 U989 ( .A1(n1304), .A2(G217), .ZN(n1303) );
NAND2_X1 U990 ( .A1(n1305), .A2(n1306), .ZN(n1302) );
OR2_X1 U991 ( .A1(n1307), .A2(G107), .ZN(n1306) );
XOR2_X1 U992 ( .A(n1308), .B(KEYINPUT38), .Z(n1305) );
NAND2_X1 U993 ( .A1(G107), .A2(n1307), .ZN(n1308) );
XOR2_X1 U994 ( .A(G116), .B(n1294), .Z(n1307) );
INV_X1 U995 ( .A(n1228), .ZN(n1162) );
NAND2_X1 U996 ( .A1(n1039), .A2(n1309), .ZN(n1228) );
NAND3_X1 U997 ( .A1(n1125), .A2(n1258), .A3(G902), .ZN(n1309) );
NOR2_X1 U998 ( .A1(n1061), .A2(G898), .ZN(n1125) );
NAND3_X1 U999 ( .A1(n1258), .A2(n1061), .A3(G952), .ZN(n1039) );
NAND2_X1 U1000 ( .A1(G237), .A2(n1310), .ZN(n1258) );
INV_X1 U1001 ( .A(n1227), .ZN(n1213) );
NOR2_X1 U1002 ( .A1(n1208), .A2(n1069), .ZN(n1227) );
INV_X1 U1003 ( .A(n1235), .ZN(n1069) );
NOR2_X1 U1004 ( .A1(n1071), .A2(n1072), .ZN(n1235) );
NOR2_X1 U1005 ( .A1(n1311), .A2(n1086), .ZN(n1072) );
NOR2_X1 U1006 ( .A1(n1312), .A2(G469), .ZN(n1086) );
XNOR2_X1 U1007 ( .A(KEYINPUT28), .B(n1082), .ZN(n1311) );
AND2_X1 U1008 ( .A1(G469), .A2(n1312), .ZN(n1082) );
NAND2_X1 U1009 ( .A1(n1313), .A2(n1280), .ZN(n1312) );
XOR2_X1 U1010 ( .A(n1189), .B(n1314), .Z(n1313) );
XNOR2_X1 U1011 ( .A(G140), .B(n1315), .ZN(n1314) );
NOR2_X1 U1012 ( .A1(KEYINPUT4), .A2(n1191), .ZN(n1315) );
XNOR2_X1 U1013 ( .A(n1316), .B(n1317), .ZN(n1191) );
XNOR2_X1 U1014 ( .A(n1240), .B(n1318), .ZN(n1317) );
NOR2_X1 U1015 ( .A1(KEYINPUT49), .A2(n1300), .ZN(n1318) );
XOR2_X1 U1016 ( .A(n1319), .B(n1320), .Z(n1189) );
XOR2_X1 U1017 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1018 ( .A(G110), .B(n1323), .ZN(n1322) );
NOR2_X1 U1019 ( .A1(G104), .A2(KEYINPUT63), .ZN(n1323) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1061), .ZN(n1321) );
XNOR2_X1 U1021 ( .A(n1177), .B(n1324), .ZN(n1319) );
INV_X1 U1022 ( .A(n1269), .ZN(n1071) );
NAND2_X1 U1023 ( .A1(G221), .A2(n1325), .ZN(n1269) );
INV_X1 U1024 ( .A(n1075), .ZN(n1208) );
NOR2_X1 U1025 ( .A1(n1087), .A2(n1064), .ZN(n1075) );
INV_X1 U1026 ( .A(n1038), .ZN(n1064) );
NAND2_X1 U1027 ( .A1(n1326), .A2(n1085), .ZN(n1038) );
NAND2_X1 U1028 ( .A1(n1092), .A2(n1094), .ZN(n1085) );
OR2_X1 U1029 ( .A1(n1094), .A2(n1092), .ZN(n1326) );
AND2_X1 U1030 ( .A1(n1327), .A2(n1280), .ZN(n1092) );
XOR2_X1 U1031 ( .A(n1231), .B(KEYINPUT29), .Z(n1327) );
XOR2_X1 U1032 ( .A(n1328), .B(n1329), .Z(n1231) );
XOR2_X1 U1033 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1034 ( .A(n1117), .B(n1332), .ZN(n1331) );
NOR2_X1 U1035 ( .A1(KEYINPUT19), .A2(n1333), .ZN(n1332) );
XNOR2_X1 U1036 ( .A(n1130), .B(n1334), .ZN(n1333) );
XNOR2_X1 U1037 ( .A(n1131), .B(KEYINPUT53), .ZN(n1334) );
XNOR2_X1 U1038 ( .A(n1335), .B(n1336), .ZN(n1131) );
XNOR2_X1 U1039 ( .A(G119), .B(n1268), .ZN(n1336) );
NAND2_X1 U1040 ( .A1(KEYINPUT33), .A2(n1266), .ZN(n1335) );
XOR2_X1 U1041 ( .A(G104), .B(n1324), .Z(n1130) );
XOR2_X1 U1042 ( .A(G101), .B(G107), .Z(n1324) );
NOR2_X1 U1043 ( .A1(G953), .A2(n1141), .ZN(n1330) );
INV_X1 U1044 ( .A(G224), .ZN(n1141) );
XNOR2_X1 U1045 ( .A(n1174), .B(n1128), .ZN(n1328) );
XNOR2_X1 U1046 ( .A(n1274), .B(n1294), .ZN(n1128) );
XOR2_X1 U1047 ( .A(G122), .B(KEYINPUT43), .Z(n1294) );
INV_X1 U1048 ( .A(G110), .ZN(n1274) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1337), .ZN(n1094) );
INV_X1 U1050 ( .A(n1041), .ZN(n1087) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1337), .ZN(n1041) );
NAND2_X1 U1052 ( .A1(n1285), .A2(n1280), .ZN(n1337) );
NOR2_X1 U1053 ( .A1(n1265), .A2(n1263), .ZN(n1074) );
XOR2_X1 U1054 ( .A(n1338), .B(n1095), .Z(n1263) );
NAND2_X1 U1055 ( .A1(n1339), .A2(n1280), .ZN(n1095) );
XOR2_X1 U1056 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1057 ( .A(n1174), .B(n1183), .ZN(n1341) );
XOR2_X1 U1058 ( .A(n1342), .B(n1343), .Z(n1183) );
XNOR2_X1 U1059 ( .A(G119), .B(n1266), .ZN(n1343) );
INV_X1 U1060 ( .A(G116), .ZN(n1266) );
NAND2_X1 U1061 ( .A1(KEYINPUT1), .A2(n1268), .ZN(n1342) );
INV_X1 U1062 ( .A(G113), .ZN(n1268) );
XOR2_X1 U1063 ( .A(n1344), .B(n1316), .Z(n1174) );
XNOR2_X1 U1064 ( .A(n1345), .B(n1346), .ZN(n1344) );
NAND2_X1 U1065 ( .A1(KEYINPUT32), .A2(n1240), .ZN(n1346) );
INV_X1 U1066 ( .A(G143), .ZN(n1240) );
NAND2_X1 U1067 ( .A1(KEYINPUT0), .A2(G128), .ZN(n1345) );
XNOR2_X1 U1068 ( .A(n1173), .B(n1347), .ZN(n1340) );
XOR2_X1 U1069 ( .A(G101), .B(n1348), .Z(n1347) );
NOR2_X1 U1070 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1348) );
NAND3_X1 U1071 ( .A1(n1285), .A2(n1061), .A3(G210), .ZN(n1168) );
INV_X1 U1072 ( .A(G237), .ZN(n1285) );
INV_X1 U1073 ( .A(n1177), .ZN(n1173) );
XNOR2_X1 U1074 ( .A(n1349), .B(n1350), .ZN(n1177) );
XNOR2_X1 U1075 ( .A(n1246), .B(G131), .ZN(n1350) );
NAND2_X1 U1076 ( .A1(KEYINPUT42), .A2(n1249), .ZN(n1349) );
INV_X1 U1077 ( .A(G134), .ZN(n1249) );
NAND2_X1 U1078 ( .A1(KEYINPUT61), .A2(G472), .ZN(n1338) );
XNOR2_X1 U1079 ( .A(n1103), .B(n1351), .ZN(n1265) );
NOR2_X1 U1080 ( .A1(n1106), .A2(KEYINPUT2), .ZN(n1351) );
NOR2_X1 U1081 ( .A1(n1352), .A2(G902), .ZN(n1106) );
INV_X1 U1082 ( .A(n1147), .ZN(n1352) );
XNOR2_X1 U1083 ( .A(n1353), .B(n1354), .ZN(n1147) );
XOR2_X1 U1084 ( .A(n1355), .B(n1356), .Z(n1354) );
NAND2_X1 U1085 ( .A1(KEYINPUT58), .A2(n1246), .ZN(n1356) );
INV_X1 U1086 ( .A(G137), .ZN(n1246) );
NAND2_X1 U1087 ( .A1(n1357), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1088 ( .A1(KEYINPUT55), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1089 ( .A(n1360), .B(n1361), .Z(n1357) );
NOR2_X1 U1090 ( .A1(KEYINPUT55), .A2(n1359), .ZN(n1361) );
XNOR2_X1 U1091 ( .A(G110), .B(n1362), .ZN(n1359) );
XNOR2_X1 U1092 ( .A(n1300), .B(G119), .ZN(n1362) );
INV_X1 U1093 ( .A(G128), .ZN(n1300) );
NAND2_X1 U1094 ( .A1(n1363), .A2(n1364), .ZN(n1360) );
NAND3_X1 U1095 ( .A1(n1365), .A2(n1288), .A3(n1366), .ZN(n1364) );
XNOR2_X1 U1096 ( .A(KEYINPUT24), .B(n1295), .ZN(n1365) );
NAND2_X1 U1097 ( .A1(n1367), .A2(n1368), .ZN(n1363) );
NAND2_X1 U1098 ( .A1(n1366), .A2(n1288), .ZN(n1368) );
NAND2_X1 U1099 ( .A1(n1369), .A2(n1117), .ZN(n1288) );
INV_X1 U1100 ( .A(G125), .ZN(n1117) );
XNOR2_X1 U1101 ( .A(KEYINPUT46), .B(G140), .ZN(n1369) );
XOR2_X1 U1102 ( .A(n1289), .B(KEYINPUT57), .Z(n1366) );
NAND2_X1 U1103 ( .A1(G125), .A2(n1370), .ZN(n1289) );
XNOR2_X1 U1104 ( .A(KEYINPUT46), .B(n1242), .ZN(n1370) );
INV_X1 U1105 ( .A(G140), .ZN(n1242) );
XNOR2_X1 U1106 ( .A(KEYINPUT24), .B(n1316), .ZN(n1367) );
INV_X1 U1107 ( .A(n1295), .ZN(n1316) );
XOR2_X1 U1108 ( .A(G146), .B(KEYINPUT30), .Z(n1295) );
NAND2_X1 U1109 ( .A1(G221), .A2(n1304), .ZN(n1353) );
AND2_X1 U1110 ( .A1(G234), .A2(n1061), .ZN(n1304) );
INV_X1 U1111 ( .A(G953), .ZN(n1061) );
NAND2_X1 U1112 ( .A1(G217), .A2(n1325), .ZN(n1103) );
NAND2_X1 U1113 ( .A1(n1310), .A2(n1280), .ZN(n1325) );
INV_X1 U1114 ( .A(G902), .ZN(n1280) );
XOR2_X1 U1115 ( .A(G234), .B(KEYINPUT47), .Z(n1310) );
endmodule


