//Key = 0110011101010010001111101110110100000110101001100011110100101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313;

XNOR2_X1 U731 ( .A(G107), .B(n1003), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1004), .A2(n1005), .ZN(G75) );
XOR2_X1 U733 ( .A(n1006), .B(KEYINPUT26), .Z(n1005) );
OR2_X1 U734 ( .A1(n1007), .A2(G952), .ZN(n1006) );
NOR4_X1 U735 ( .A1(n1008), .A2(n1007), .A3(n1009), .A4(n1010), .ZN(n1004) );
INV_X1 U736 ( .A(G952), .ZN(n1009) );
NAND2_X1 U737 ( .A1(n1011), .A2(n1012), .ZN(n1007) );
NAND4_X1 U738 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR4_X1 U739 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
XNOR2_X1 U740 ( .A(n1021), .B(n1022), .ZN(n1018) );
XNOR2_X1 U741 ( .A(n1023), .B(n1024), .ZN(n1017) );
NAND2_X1 U742 ( .A1(n1025), .A2(KEYINPUT7), .ZN(n1023) );
XNOR2_X1 U743 ( .A(G469), .B(KEYINPUT13), .ZN(n1025) );
NOR3_X1 U744 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1015) );
AND2_X1 U745 ( .A1(n1029), .A2(G478), .ZN(n1026) );
XOR2_X1 U746 ( .A(n1030), .B(n1031), .Z(n1014) );
NOR2_X1 U747 ( .A1(n1032), .A2(KEYINPUT56), .ZN(n1031) );
XOR2_X1 U748 ( .A(KEYINPUT53), .B(n1033), .Z(n1013) );
NOR2_X1 U749 ( .A1(G478), .A2(n1029), .ZN(n1033) );
NAND3_X1 U750 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1008) );
NAND2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND3_X1 U752 ( .A1(n1039), .A2(n1040), .A3(n1027), .ZN(n1035) );
XOR2_X1 U753 ( .A(KEYINPUT0), .B(n1037), .Z(n1040) );
AND2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1037) );
NAND2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(n1034) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U757 ( .A1(KEYINPUT16), .A2(n1047), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1041), .A2(n1048), .ZN(n1047) );
AND3_X1 U759 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1041) );
NAND2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U762 ( .A1(n1049), .A2(n1055), .A3(n1042), .ZN(n1054) );
OR2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U764 ( .A1(n1050), .A2(n1058), .ZN(n1053) );
NAND2_X1 U765 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U766 ( .A1(n1049), .A2(n1061), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U768 ( .A1(n1048), .A2(n1064), .ZN(n1063) );
INV_X1 U769 ( .A(KEYINPUT16), .ZN(n1064) );
OR2_X1 U770 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U771 ( .A1(n1042), .A2(n1067), .ZN(n1059) );
NAND2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
INV_X1 U774 ( .A(n1072), .ZN(n1051) );
XOR2_X1 U775 ( .A(n1073), .B(n1074), .Z(G72) );
NOR2_X1 U776 ( .A1(n1075), .A2(n1011), .ZN(n1074) );
NOR2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U778 ( .A1(KEYINPUT47), .A2(n1078), .ZN(n1073) );
XOR2_X1 U779 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U780 ( .A1(n1081), .A2(G953), .ZN(n1080) );
NOR2_X1 U781 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U782 ( .A(KEYINPUT17), .B(n1084), .ZN(n1083) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(n1079) );
NAND2_X1 U784 ( .A1(G953), .A2(n1077), .ZN(n1086) );
XOR2_X1 U785 ( .A(n1087), .B(n1088), .Z(n1085) );
XOR2_X1 U786 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U787 ( .A1(G125), .A2(KEYINPUT15), .ZN(n1090) );
NAND2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND3_X1 U789 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NAND2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U791 ( .A1(KEYINPUT51), .A2(n1098), .ZN(n1096) );
XOR2_X1 U792 ( .A(KEYINPUT55), .B(n1099), .Z(n1098) );
NAND2_X1 U793 ( .A1(KEYINPUT44), .A2(n1100), .ZN(n1094) );
NAND2_X1 U794 ( .A1(G131), .A2(n1101), .ZN(n1100) );
NAND2_X1 U795 ( .A1(n1102), .A2(n1103), .ZN(n1093) );
NAND2_X1 U796 ( .A1(n1104), .A2(n1105), .ZN(n1091) );
NAND2_X1 U797 ( .A1(KEYINPUT51), .A2(n1106), .ZN(n1105) );
NAND3_X1 U798 ( .A1(n1107), .A2(n1108), .A3(n1097), .ZN(n1106) );
INV_X1 U799 ( .A(KEYINPUT61), .ZN(n1097) );
NAND2_X1 U800 ( .A1(n1109), .A2(n1103), .ZN(n1108) );
INV_X1 U801 ( .A(KEYINPUT44), .ZN(n1103) );
NAND3_X1 U802 ( .A1(G131), .A2(n1101), .A3(KEYINPUT44), .ZN(n1107) );
XNOR2_X1 U803 ( .A(n1099), .B(KEYINPUT55), .ZN(n1104) );
XNOR2_X1 U804 ( .A(G140), .B(KEYINPUT58), .ZN(n1087) );
XOR2_X1 U805 ( .A(n1110), .B(n1111), .Z(G69) );
XOR2_X1 U806 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U807 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1114) );
NAND3_X1 U809 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1112) );
XOR2_X1 U810 ( .A(KEYINPUT2), .B(n1118), .Z(n1117) );
NOR2_X1 U811 ( .A1(G898), .A2(n1011), .ZN(n1118) );
NAND2_X1 U812 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
NAND2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NAND2_X1 U814 ( .A1(KEYINPUT6), .A2(n1123), .ZN(n1122) );
OR2_X1 U815 ( .A1(n1124), .A2(KEYINPUT6), .ZN(n1121) );
OR2_X1 U816 ( .A1(n1120), .A2(n1123), .ZN(n1115) );
OR2_X1 U817 ( .A1(KEYINPUT32), .A2(n1124), .ZN(n1123) );
XNOR2_X1 U818 ( .A(G110), .B(n1125), .ZN(n1124) );
NOR2_X1 U819 ( .A1(n1126), .A2(G953), .ZN(n1110) );
NOR2_X1 U820 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U821 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U822 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U823 ( .A1(n1127), .A2(n1133), .ZN(G63) );
NOR2_X1 U824 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U825 ( .A(n1136), .B(KEYINPUT5), .Z(n1135) );
NAND2_X1 U826 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U827 ( .A1(n1139), .A2(G478), .ZN(n1138) );
XOR2_X1 U828 ( .A(KEYINPUT42), .B(n1140), .Z(n1137) );
AND3_X1 U829 ( .A1(n1139), .A2(n1140), .A3(G478), .ZN(n1134) );
XOR2_X1 U830 ( .A(n1141), .B(KEYINPUT14), .Z(n1140) );
NOR2_X1 U831 ( .A1(n1127), .A2(n1142), .ZN(G60) );
XOR2_X1 U832 ( .A(n1143), .B(KEYINPUT4), .Z(n1142) );
NAND2_X1 U833 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U834 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U835 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NAND2_X1 U836 ( .A1(KEYINPUT9), .A2(n1150), .ZN(n1149) );
INV_X1 U837 ( .A(KEYINPUT10), .ZN(n1148) );
NAND2_X1 U838 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
NAND2_X1 U839 ( .A1(KEYINPUT9), .A2(n1153), .ZN(n1152) );
OR2_X1 U840 ( .A1(n1147), .A2(KEYINPUT10), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1139), .A2(G475), .ZN(n1147) );
INV_X1 U842 ( .A(n1150), .ZN(n1151) );
XNOR2_X1 U843 ( .A(G104), .B(n1154), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1127), .A2(n1155), .ZN(G57) );
XOR2_X1 U845 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U846 ( .A(n1158), .B(n1099), .Z(n1157) );
XOR2_X1 U847 ( .A(n1159), .B(n1160), .Z(n1156) );
AND2_X1 U848 ( .A1(G472), .A2(n1139), .ZN(n1160) );
NOR2_X1 U849 ( .A1(n1127), .A2(n1161), .ZN(G54) );
XOR2_X1 U850 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U851 ( .A(n1109), .B(n1164), .ZN(n1163) );
NOR3_X1 U852 ( .A1(n1132), .A2(KEYINPUT59), .A3(n1165), .ZN(n1164) );
INV_X1 U853 ( .A(G469), .ZN(n1165) );
NOR2_X1 U854 ( .A1(n1127), .A2(n1166), .ZN(G51) );
XOR2_X1 U855 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n1169), .ZN(n1168) );
NAND2_X1 U857 ( .A1(n1139), .A2(n1032), .ZN(n1167) );
INV_X1 U858 ( .A(n1132), .ZN(n1139) );
NAND2_X1 U859 ( .A1(G902), .A2(n1010), .ZN(n1132) );
NAND3_X1 U860 ( .A1(n1170), .A2(n1084), .A3(n1126), .ZN(n1010) );
AND2_X1 U861 ( .A1(n1171), .A2(n1172), .ZN(n1126) );
AND4_X1 U862 ( .A1(n1003), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1172) );
NAND3_X1 U863 ( .A1(n1057), .A2(n1049), .A3(n1176), .ZN(n1003) );
AND4_X1 U864 ( .A1(n1177), .A2(n1178), .A3(n1154), .A4(n1179), .ZN(n1171) );
OR4_X1 U865 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
XOR2_X1 U866 ( .A(n1184), .B(KEYINPUT19), .Z(n1180) );
NAND3_X1 U867 ( .A1(n1176), .A2(n1049), .A3(n1056), .ZN(n1154) );
INV_X1 U868 ( .A(n1181), .ZN(n1049) );
INV_X1 U869 ( .A(n1082), .ZN(n1170) );
NAND4_X1 U870 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1082) );
NOR4_X1 U871 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
INV_X1 U872 ( .A(n1193), .ZN(n1192) );
NOR2_X1 U873 ( .A1(n1011), .A2(G952), .ZN(n1127) );
XNOR2_X1 U874 ( .A(G146), .B(n1187), .ZN(G48) );
NAND3_X1 U875 ( .A1(n1056), .A2(n1038), .A3(n1194), .ZN(n1187) );
XNOR2_X1 U876 ( .A(G143), .B(n1185), .ZN(G45) );
NAND3_X1 U877 ( .A1(n1195), .A2(n1038), .A3(n1196), .ZN(n1185) );
XNOR2_X1 U878 ( .A(G140), .B(n1186), .ZN(G42) );
NAND3_X1 U879 ( .A1(n1043), .A2(n1048), .A3(n1197), .ZN(n1186) );
XOR2_X1 U880 ( .A(n1198), .B(n1199), .Z(G39) );
NOR2_X1 U881 ( .A1(KEYINPUT23), .A2(n1193), .ZN(n1199) );
NAND3_X1 U882 ( .A1(n1043), .A2(n1050), .A3(n1194), .ZN(n1193) );
XNOR2_X1 U883 ( .A(G137), .B(KEYINPUT38), .ZN(n1198) );
XOR2_X1 U884 ( .A(G134), .B(n1200), .Z(G36) );
NOR2_X1 U885 ( .A1(KEYINPUT8), .A2(n1084), .ZN(n1200) );
NAND3_X1 U886 ( .A1(n1196), .A2(n1057), .A3(n1043), .ZN(n1084) );
XOR2_X1 U887 ( .A(G131), .B(n1191), .Z(G33) );
AND3_X1 U888 ( .A1(n1196), .A2(n1056), .A3(n1043), .ZN(n1191) );
NOR2_X1 U889 ( .A1(n1201), .A2(n1027), .ZN(n1043) );
AND3_X1 U890 ( .A1(n1048), .A2(n1202), .A3(n1203), .ZN(n1196) );
XOR2_X1 U891 ( .A(G128), .B(n1190), .Z(G30) );
AND3_X1 U892 ( .A1(n1057), .A2(n1038), .A3(n1194), .ZN(n1190) );
AND4_X1 U893 ( .A1(n1048), .A2(n1020), .A3(n1204), .A4(n1202), .ZN(n1194) );
XOR2_X1 U894 ( .A(n1178), .B(n1205), .Z(G3) );
XNOR2_X1 U895 ( .A(G101), .B(KEYINPUT35), .ZN(n1205) );
NAND3_X1 U896 ( .A1(n1176), .A2(n1050), .A3(n1203), .ZN(n1178) );
XOR2_X1 U897 ( .A(G125), .B(n1189), .Z(G27) );
AND2_X1 U898 ( .A1(n1197), .A2(n1206), .ZN(n1189) );
AND4_X1 U899 ( .A1(n1070), .A2(n1056), .A3(n1071), .A4(n1202), .ZN(n1197) );
NAND2_X1 U900 ( .A1(n1072), .A2(n1207), .ZN(n1202) );
NAND4_X1 U901 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1077), .ZN(n1207) );
INV_X1 U902 ( .A(G900), .ZN(n1077) );
XOR2_X1 U903 ( .A(n1209), .B(n1210), .Z(G24) );
NOR2_X1 U904 ( .A1(KEYINPUT34), .A2(n1125), .ZN(n1210) );
NOR3_X1 U905 ( .A1(n1211), .A2(n1212), .A3(n1181), .ZN(n1209) );
NAND2_X1 U906 ( .A1(n1071), .A2(n1213), .ZN(n1181) );
XNOR2_X1 U907 ( .A(n1195), .B(KEYINPUT54), .ZN(n1212) );
INV_X1 U908 ( .A(n1183), .ZN(n1195) );
NAND2_X1 U909 ( .A1(n1214), .A2(n1215), .ZN(n1183) );
XNOR2_X1 U910 ( .A(n1216), .B(n1217), .ZN(G21) );
NOR2_X1 U911 ( .A1(n1218), .A2(n1177), .ZN(n1217) );
NAND4_X1 U912 ( .A1(n1219), .A2(n1050), .A3(n1020), .A4(n1204), .ZN(n1177) );
XNOR2_X1 U913 ( .A(KEYINPUT60), .B(KEYINPUT39), .ZN(n1218) );
XNOR2_X1 U914 ( .A(G116), .B(n1175), .ZN(G18) );
NAND3_X1 U915 ( .A1(n1219), .A2(n1057), .A3(n1203), .ZN(n1175) );
AND2_X1 U916 ( .A1(n1220), .A2(n1215), .ZN(n1057) );
XNOR2_X1 U917 ( .A(KEYINPUT49), .B(n1214), .ZN(n1220) );
NAND2_X1 U918 ( .A1(n1221), .A2(n1222), .ZN(G15) );
OR2_X1 U919 ( .A1(n1174), .A2(G113), .ZN(n1222) );
XOR2_X1 U920 ( .A(n1223), .B(KEYINPUT3), .Z(n1221) );
NAND2_X1 U921 ( .A1(G113), .A2(n1174), .ZN(n1223) );
NAND3_X1 U922 ( .A1(n1219), .A2(n1056), .A3(n1203), .ZN(n1174) );
INV_X1 U923 ( .A(n1068), .ZN(n1203) );
NAND2_X1 U924 ( .A1(n1020), .A2(n1213), .ZN(n1068) );
XNOR2_X1 U925 ( .A(n1224), .B(KEYINPUT11), .ZN(n1213) );
INV_X1 U926 ( .A(n1204), .ZN(n1224) );
INV_X1 U927 ( .A(n1211), .ZN(n1219) );
NAND2_X1 U928 ( .A1(n1206), .A2(n1184), .ZN(n1211) );
INV_X1 U929 ( .A(n1182), .ZN(n1206) );
NAND2_X1 U930 ( .A1(n1042), .A2(n1038), .ZN(n1182) );
NOR2_X1 U931 ( .A1(n1065), .A2(n1028), .ZN(n1042) );
INV_X1 U932 ( .A(n1066), .ZN(n1028) );
XNOR2_X1 U933 ( .A(G110), .B(n1173), .ZN(G12) );
NAND4_X1 U934 ( .A1(n1070), .A2(n1176), .A3(n1071), .A4(n1050), .ZN(n1173) );
NAND2_X1 U935 ( .A1(n1225), .A2(n1226), .ZN(n1050) );
OR3_X1 U936 ( .A1(n1214), .A2(n1215), .A3(KEYINPUT49), .ZN(n1226) );
INV_X1 U937 ( .A(n1227), .ZN(n1214) );
NAND2_X1 U938 ( .A1(KEYINPUT49), .A2(n1056), .ZN(n1225) );
NOR2_X1 U939 ( .A1(n1215), .A2(n1227), .ZN(n1056) );
XNOR2_X1 U940 ( .A(n1228), .B(n1229), .ZN(n1227) );
XNOR2_X1 U941 ( .A(KEYINPUT48), .B(n1230), .ZN(n1229) );
INV_X1 U942 ( .A(n1021), .ZN(n1230) );
NOR2_X1 U943 ( .A1(n1150), .A2(G902), .ZN(n1021) );
XNOR2_X1 U944 ( .A(n1231), .B(n1232), .ZN(n1150) );
XNOR2_X1 U945 ( .A(n1125), .B(G104), .ZN(n1232) );
NAND2_X1 U946 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
NAND2_X1 U947 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U948 ( .A(n1237), .B(KEYINPUT31), .Z(n1236) );
XNOR2_X1 U949 ( .A(G146), .B(n1238), .ZN(n1235) );
NAND2_X1 U950 ( .A1(n1237), .A2(n1239), .ZN(n1233) );
XOR2_X1 U951 ( .A(G146), .B(n1238), .Z(n1239) );
XOR2_X1 U952 ( .A(n1240), .B(n1241), .Z(n1237) );
XOR2_X1 U953 ( .A(n1242), .B(n1243), .Z(n1241) );
NAND2_X1 U954 ( .A1(KEYINPUT46), .A2(G131), .ZN(n1243) );
NAND2_X1 U955 ( .A1(n1244), .A2(G214), .ZN(n1242) );
XNOR2_X1 U956 ( .A(G143), .B(n1245), .ZN(n1240) );
NOR2_X1 U957 ( .A1(KEYINPUT41), .A2(n1246), .ZN(n1245) );
INV_X1 U958 ( .A(G113), .ZN(n1246) );
NAND2_X1 U959 ( .A1(KEYINPUT21), .A2(n1022), .ZN(n1228) );
XOR2_X1 U960 ( .A(G475), .B(KEYINPUT28), .Z(n1022) );
XOR2_X1 U961 ( .A(n1247), .B(n1029), .Z(n1215) );
NAND2_X1 U962 ( .A1(n1141), .A2(n1248), .ZN(n1029) );
XNOR2_X1 U963 ( .A(n1249), .B(n1250), .ZN(n1141) );
XNOR2_X1 U964 ( .A(n1251), .B(n1252), .ZN(n1250) );
NAND2_X1 U965 ( .A1(KEYINPUT25), .A2(n1253), .ZN(n1251) );
XOR2_X1 U966 ( .A(G107), .B(n1254), .Z(n1253) );
XNOR2_X1 U967 ( .A(n1125), .B(G116), .ZN(n1254) );
XOR2_X1 U968 ( .A(n1255), .B(G134), .Z(n1249) );
NAND2_X1 U969 ( .A1(G217), .A2(n1256), .ZN(n1255) );
NAND2_X1 U970 ( .A1(KEYINPUT24), .A2(G478), .ZN(n1247) );
INV_X1 U971 ( .A(n1020), .ZN(n1071) );
XNOR2_X1 U972 ( .A(n1257), .B(G472), .ZN(n1020) );
NAND2_X1 U973 ( .A1(n1258), .A2(n1248), .ZN(n1257) );
XOR2_X1 U974 ( .A(n1158), .B(n1259), .Z(n1258) );
XOR2_X1 U975 ( .A(n1260), .B(n1159), .Z(n1259) );
XNOR2_X1 U976 ( .A(n1261), .B(n1262), .ZN(n1159) );
NAND2_X1 U977 ( .A1(n1244), .A2(G210), .ZN(n1261) );
NOR2_X1 U978 ( .A1(G953), .A2(G237), .ZN(n1244) );
NAND2_X1 U979 ( .A1(KEYINPUT18), .A2(n1099), .ZN(n1260) );
XNOR2_X1 U980 ( .A(n1102), .B(n1263), .ZN(n1158) );
AND3_X1 U981 ( .A1(n1038), .A2(n1184), .A3(n1048), .ZN(n1176) );
AND2_X1 U982 ( .A1(n1264), .A2(n1065), .ZN(n1048) );
XNOR2_X1 U983 ( .A(n1024), .B(G469), .ZN(n1065) );
NAND2_X1 U984 ( .A1(n1265), .A2(n1248), .ZN(n1024) );
XOR2_X1 U985 ( .A(n1162), .B(n1266), .Z(n1265) );
XNOR2_X1 U986 ( .A(KEYINPUT1), .B(n1267), .ZN(n1266) );
NOR2_X1 U987 ( .A1(KEYINPUT43), .A2(n1102), .ZN(n1267) );
INV_X1 U988 ( .A(n1109), .ZN(n1102) );
XOR2_X1 U989 ( .A(G131), .B(n1101), .Z(n1109) );
XNOR2_X1 U990 ( .A(G134), .B(n1268), .ZN(n1101) );
XNOR2_X1 U991 ( .A(n1269), .B(n1270), .ZN(n1162) );
INV_X1 U992 ( .A(G140), .ZN(n1270) );
XOR2_X1 U993 ( .A(n1271), .B(n1272), .Z(n1269) );
XOR2_X1 U994 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U995 ( .A(KEYINPUT27), .B(G104), .Z(n1274) );
XOR2_X1 U996 ( .A(KEYINPUT55), .B(KEYINPUT37), .Z(n1273) );
XOR2_X1 U997 ( .A(n1275), .B(n1276), .Z(n1271) );
XNOR2_X1 U998 ( .A(n1262), .B(n1277), .ZN(n1276) );
NOR2_X1 U999 ( .A1(G953), .A2(n1076), .ZN(n1277) );
INV_X1 U1000 ( .A(G227), .ZN(n1076) );
INV_X1 U1001 ( .A(G101), .ZN(n1262) );
XOR2_X1 U1002 ( .A(n1278), .B(n1279), .Z(n1275) );
NOR2_X1 U1003 ( .A1(G107), .A2(KEYINPUT12), .ZN(n1279) );
XNOR2_X1 U1004 ( .A(KEYINPUT52), .B(n1066), .ZN(n1264) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1280), .ZN(n1066) );
NAND2_X1 U1006 ( .A1(n1072), .A2(n1281), .ZN(n1184) );
NAND4_X1 U1007 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1282), .ZN(n1281) );
INV_X1 U1008 ( .A(G898), .ZN(n1282) );
NAND3_X1 U1009 ( .A1(n1208), .A2(n1011), .A3(G952), .ZN(n1072) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1208) );
NOR2_X1 U1011 ( .A1(n1039), .A2(n1027), .ZN(n1038) );
AND2_X1 U1012 ( .A1(G214), .A2(n1283), .ZN(n1027) );
INV_X1 U1013 ( .A(n1201), .ZN(n1039) );
XNOR2_X1 U1014 ( .A(n1284), .B(n1032), .ZN(n1201) );
AND2_X1 U1015 ( .A1(G210), .A2(n1283), .ZN(n1032) );
OR2_X1 U1016 ( .A1(G902), .A2(G237), .ZN(n1283) );
NAND2_X1 U1017 ( .A1(KEYINPUT45), .A2(n1030), .ZN(n1284) );
AND2_X1 U1018 ( .A1(n1285), .A2(n1248), .ZN(n1030) );
XOR2_X1 U1019 ( .A(KEYINPUT40), .B(n1169), .Z(n1285) );
XNOR2_X1 U1020 ( .A(n1286), .B(n1287), .ZN(n1169) );
XOR2_X1 U1021 ( .A(n1288), .B(n1278), .Z(n1287) );
XNOR2_X1 U1022 ( .A(G110), .B(n1099), .ZN(n1278) );
XOR2_X1 U1023 ( .A(G146), .B(n1252), .Z(n1099) );
XNOR2_X1 U1024 ( .A(G128), .B(n1289), .ZN(n1252) );
INV_X1 U1025 ( .A(G143), .ZN(n1289) );
NAND2_X1 U1026 ( .A1(KEYINPUT22), .A2(n1120), .ZN(n1288) );
XOR2_X1 U1027 ( .A(n1290), .B(n1291), .Z(n1120) );
XOR2_X1 U1028 ( .A(G107), .B(G104), .Z(n1291) );
XNOR2_X1 U1029 ( .A(G101), .B(n1263), .ZN(n1290) );
XNOR2_X1 U1030 ( .A(n1292), .B(n1293), .ZN(n1263) );
XNOR2_X1 U1031 ( .A(KEYINPUT30), .B(n1216), .ZN(n1293) );
INV_X1 U1032 ( .A(G119), .ZN(n1216) );
XNOR2_X1 U1033 ( .A(G116), .B(G113), .ZN(n1292) );
XOR2_X1 U1034 ( .A(n1294), .B(n1295), .Z(n1286) );
XNOR2_X1 U1035 ( .A(G125), .B(n1125), .ZN(n1295) );
INV_X1 U1036 ( .A(G122), .ZN(n1125) );
NAND2_X1 U1037 ( .A1(G224), .A2(n1011), .ZN(n1294) );
XNOR2_X1 U1038 ( .A(n1204), .B(KEYINPUT29), .ZN(n1070) );
XOR2_X1 U1039 ( .A(n1019), .B(KEYINPUT36), .Z(n1204) );
XNOR2_X1 U1040 ( .A(n1131), .B(n1296), .ZN(n1019) );
NOR2_X1 U1041 ( .A1(G902), .A2(n1129), .ZN(n1296) );
XOR2_X1 U1042 ( .A(n1297), .B(n1298), .Z(n1129) );
XOR2_X1 U1043 ( .A(n1299), .B(n1238), .Z(n1298) );
XOR2_X1 U1044 ( .A(G125), .B(G140), .Z(n1238) );
NOR2_X1 U1045 ( .A1(G146), .A2(KEYINPUT57), .ZN(n1299) );
XOR2_X1 U1046 ( .A(n1300), .B(n1301), .Z(n1297) );
NOR2_X1 U1047 ( .A1(KEYINPUT62), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1048 ( .A(n1303), .B(n1304), .Z(n1302) );
NAND2_X1 U1049 ( .A1(KEYINPUT20), .A2(n1268), .ZN(n1304) );
INV_X1 U1050 ( .A(G137), .ZN(n1268) );
NAND2_X1 U1051 ( .A1(n1256), .A2(G221), .ZN(n1303) );
AND2_X1 U1052 ( .A1(G234), .A2(n1011), .ZN(n1256) );
INV_X1 U1053 ( .A(G953), .ZN(n1011) );
NAND2_X1 U1054 ( .A1(n1305), .A2(n1306), .ZN(n1300) );
NAND2_X1 U1055 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1056 ( .A1(KEYINPUT50), .A2(n1309), .ZN(n1308) );
NAND2_X1 U1057 ( .A1(KEYINPUT63), .A2(G110), .ZN(n1309) );
INV_X1 U1058 ( .A(n1310), .ZN(n1307) );
NAND2_X1 U1059 ( .A1(n1311), .A2(n1312), .ZN(n1305) );
INV_X1 U1060 ( .A(G110), .ZN(n1312) );
NAND2_X1 U1061 ( .A1(KEYINPUT63), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1062 ( .A1(KEYINPUT50), .A2(n1310), .ZN(n1313) );
XOR2_X1 U1063 ( .A(G119), .B(G128), .Z(n1310) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1280), .ZN(n1131) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1248), .ZN(n1280) );
INV_X1 U1066 ( .A(G902), .ZN(n1248) );
endmodule


