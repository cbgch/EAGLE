//Key = 0101011110111110110110101101010011010100010000001001011001001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291;

XOR2_X1 U717 ( .A(n994), .B(n995), .Z(G9) );
NOR2_X1 U718 ( .A1(KEYINPUT9), .A2(n996), .ZN(n995) );
NAND4_X1 U719 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(G75) );
NAND4_X1 U720 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n999) );
NOR4_X1 U721 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
XNOR2_X1 U722 ( .A(KEYINPUT39), .B(n1009), .ZN(n1008) );
XOR2_X1 U723 ( .A(KEYINPUT36), .B(n1010), .Z(n1007) );
XNOR2_X1 U724 ( .A(n1011), .B(n1012), .ZN(n1006) );
NOR3_X1 U725 ( .A1(n1013), .A2(KEYINPUT56), .A3(G902), .ZN(n1011) );
NOR2_X1 U726 ( .A1(n1014), .A2(n1015), .ZN(n1003) );
XNOR2_X1 U727 ( .A(G469), .B(n1016), .ZN(n1002) );
NAND2_X1 U728 ( .A1(KEYINPUT33), .A2(n1017), .ZN(n1016) );
XNOR2_X1 U729 ( .A(KEYINPUT3), .B(n1018), .ZN(n1001) );
NAND2_X1 U730 ( .A1(n1019), .A2(n1020), .ZN(n998) );
NAND2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND4_X1 U732 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NAND2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND2_X1 U734 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U736 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U737 ( .A1(n1035), .A2(n1036), .ZN(n1027) );
NAND2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U739 ( .A1(n1014), .A2(n1018), .ZN(n1038) );
XOR2_X1 U740 ( .A(KEYINPUT10), .B(n1039), .Z(n1037) );
NAND3_X1 U741 ( .A1(n1035), .A2(n1040), .A3(n1029), .ZN(n1021) );
NAND3_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND3_X1 U743 ( .A1(n1024), .A2(n1044), .A3(n1026), .ZN(n1042) );
OR2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U745 ( .A1(n1023), .A2(n1024), .A3(n1015), .ZN(n1041) );
INV_X1 U746 ( .A(n1047), .ZN(n1019) );
XOR2_X1 U747 ( .A(n1048), .B(n1049), .Z(G72) );
XOR2_X1 U748 ( .A(n1050), .B(n1051), .Z(n1049) );
AND2_X1 U749 ( .A1(n1052), .A2(n1000), .ZN(n1051) );
NOR2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
XOR2_X1 U751 ( .A(n1055), .B(n1056), .Z(n1054) );
NAND3_X1 U752 ( .A1(n1057), .A2(n1058), .A3(KEYINPUT12), .ZN(n1056) );
NAND2_X1 U753 ( .A1(KEYINPUT35), .A2(n1059), .ZN(n1058) );
XOR2_X1 U754 ( .A(n1060), .B(n1061), .Z(n1059) );
NAND3_X1 U755 ( .A1(n1061), .A2(n1060), .A3(n1062), .ZN(n1057) );
INV_X1 U756 ( .A(KEYINPUT35), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1063), .A2(n1064), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XOR2_X1 U759 ( .A(KEYINPUT30), .B(G125), .Z(n1065) );
XOR2_X1 U760 ( .A(KEYINPUT13), .B(n1067), .Z(n1063) );
NOR2_X1 U761 ( .A1(G125), .A2(n1066), .ZN(n1067) );
NOR2_X1 U762 ( .A1(G900), .A2(n1000), .ZN(n1053) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1000), .ZN(n1048) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1068) );
XOR2_X1 U765 ( .A(n1069), .B(n1070), .Z(G69) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1000), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U768 ( .A(KEYINPUT16), .B(G224), .Z(n1073) );
NAND2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND2_X1 U772 ( .A1(KEYINPUT47), .A2(n1080), .ZN(n1079) );
INV_X1 U773 ( .A(n1081), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1000), .ZN(n1078) );
OR3_X1 U775 ( .A1(n1081), .A2(KEYINPUT47), .A3(n1077), .ZN(n1074) );
NAND2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U777 ( .A1(G953), .A2(n1072), .ZN(n1083) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(n1082) );
XNOR2_X1 U779 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND2_X1 U780 ( .A1(KEYINPUT60), .A2(n1088), .ZN(n1087) );
NAND2_X1 U781 ( .A1(KEYINPUT53), .A2(n1089), .ZN(n1086) );
NOR3_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(G66) );
NOR3_X1 U783 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1092) );
AND2_X1 U784 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
INV_X1 U785 ( .A(KEYINPUT42), .ZN(n1093) );
XOR2_X1 U786 ( .A(n1013), .B(n1095), .Z(n1090) );
NOR2_X1 U787 ( .A1(n1012), .A2(n1096), .ZN(n1095) );
NOR2_X1 U788 ( .A1(n1094), .A2(n1097), .ZN(G63) );
XOR2_X1 U789 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U790 ( .A1(n1100), .A2(n1101), .A3(G478), .ZN(n1098) );
XNOR2_X1 U791 ( .A(KEYINPUT62), .B(n1102), .ZN(n1100) );
NOR2_X1 U792 ( .A1(n1094), .A2(n1103), .ZN(G60) );
XOR2_X1 U793 ( .A(n1104), .B(n1105), .Z(n1103) );
AND2_X1 U794 ( .A1(G475), .A2(n1106), .ZN(n1104) );
XOR2_X1 U795 ( .A(G104), .B(n1107), .Z(G6) );
NOR2_X1 U796 ( .A1(n1094), .A2(n1108), .ZN(G57) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U799 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1112) );
XOR2_X1 U800 ( .A(n1113), .B(n1114), .Z(n1109) );
AND2_X1 U801 ( .A1(G472), .A2(n1106), .ZN(n1114) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(n1113) );
NAND2_X1 U803 ( .A1(KEYINPUT57), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U804 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1094), .A2(n1120), .ZN(G54) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U807 ( .A(n1119), .B(n1123), .Z(n1122) );
XOR2_X1 U808 ( .A(n1124), .B(n1125), .Z(n1121) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
AND2_X1 U810 ( .A1(G469), .A2(n1106), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1128), .A2(KEYINPUT41), .ZN(n1126) );
XNOR2_X1 U812 ( .A(n1129), .B(KEYINPUT5), .ZN(n1128) );
NAND2_X1 U813 ( .A1(KEYINPUT19), .A2(n1130), .ZN(n1124) );
NOR2_X1 U814 ( .A1(n1094), .A2(n1131), .ZN(G51) );
XNOR2_X1 U815 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR4_X1 U816 ( .A1(n1134), .A2(n1135), .A3(KEYINPUT0), .A4(n1136), .ZN(n1133) );
NOR2_X1 U817 ( .A1(KEYINPUT22), .A2(n1137), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1102), .A2(n1101), .ZN(n1137) );
INV_X1 U819 ( .A(n997), .ZN(n1101) );
AND2_X1 U820 ( .A1(n1096), .A2(KEYINPUT22), .ZN(n1134) );
INV_X1 U821 ( .A(n1106), .ZN(n1096) );
NOR2_X1 U822 ( .A1(n1102), .A2(n997), .ZN(n1106) );
NOR2_X1 U823 ( .A1(n1052), .A2(n1077), .ZN(n997) );
NAND2_X1 U824 ( .A1(n1138), .A2(n1139), .ZN(n1077) );
NOR4_X1 U825 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n994), .ZN(n1139) );
AND2_X1 U826 ( .A1(n1045), .A2(n1143), .ZN(n994) );
NOR4_X1 U827 ( .A1(n1107), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1138) );
NOR3_X1 U828 ( .A1(n1043), .A2(n1147), .A3(n1031), .ZN(n1146) );
AND2_X1 U829 ( .A1(n1046), .A2(n1143), .ZN(n1107) );
AND3_X1 U830 ( .A1(n1148), .A2(n1035), .A3(n1149), .ZN(n1143) );
NAND4_X1 U831 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1052) );
NOR4_X1 U832 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR3_X1 U833 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
INV_X1 U834 ( .A(n1046), .ZN(n1160) );
XOR2_X1 U835 ( .A(KEYINPUT32), .B(n1029), .Z(n1158) );
INV_X1 U836 ( .A(n1161), .ZN(n1155) );
NOR2_X1 U837 ( .A1(n1162), .A2(n1163), .ZN(n1152) );
NOR2_X1 U838 ( .A1(n1000), .A2(G952), .ZN(n1094) );
XOR2_X1 U839 ( .A(G146), .B(n1162), .Z(G48) );
AND3_X1 U840 ( .A1(n1164), .A2(n1039), .A3(n1046), .ZN(n1162) );
XNOR2_X1 U841 ( .A(n1150), .B(n1165), .ZN(G45) );
NOR2_X1 U842 ( .A1(KEYINPUT50), .A2(n1166), .ZN(n1165) );
NAND4_X1 U843 ( .A1(n1167), .A2(n1039), .A3(n1168), .A4(n1169), .ZN(n1150) );
XNOR2_X1 U844 ( .A(n1066), .B(n1154), .ZN(G42) );
AND3_X1 U845 ( .A1(n1170), .A2(n1148), .A3(n1029), .ZN(n1154) );
XOR2_X1 U846 ( .A(G137), .B(n1171), .Z(G39) );
NOR2_X1 U847 ( .A1(KEYINPUT34), .A2(n1161), .ZN(n1171) );
NAND3_X1 U848 ( .A1(n1029), .A2(n1164), .A3(n1023), .ZN(n1161) );
XNOR2_X1 U849 ( .A(G134), .B(n1172), .ZN(G36) );
NAND2_X1 U850 ( .A1(KEYINPUT48), .A2(n1156), .ZN(n1172) );
AND2_X1 U851 ( .A1(n1173), .A2(n1045), .ZN(n1156) );
XNOR2_X1 U852 ( .A(G131), .B(n1174), .ZN(G33) );
NAND2_X1 U853 ( .A1(n1173), .A2(n1046), .ZN(n1174) );
AND2_X1 U854 ( .A1(n1029), .A2(n1167), .ZN(n1173) );
INV_X1 U855 ( .A(n1159), .ZN(n1167) );
NAND3_X1 U856 ( .A1(n1148), .A2(n1175), .A3(n1176), .ZN(n1159) );
NOR2_X1 U857 ( .A1(n1177), .A2(n1014), .ZN(n1029) );
XNOR2_X1 U858 ( .A(G128), .B(n1151), .ZN(G30) );
NAND3_X1 U859 ( .A1(n1045), .A2(n1039), .A3(n1164), .ZN(n1151) );
AND4_X1 U860 ( .A1(n1034), .A2(n1148), .A3(n1005), .A4(n1175), .ZN(n1164) );
XOR2_X1 U861 ( .A(n1178), .B(n1179), .Z(G3) );
NOR4_X1 U862 ( .A1(n1180), .A2(n1031), .A3(n1043), .A4(n1181), .ZN(n1179) );
XOR2_X1 U863 ( .A(KEYINPUT7), .B(n1039), .Z(n1181) );
INV_X1 U864 ( .A(n1182), .ZN(n1180) );
NAND2_X1 U865 ( .A1(KEYINPUT1), .A2(n1183), .ZN(n1178) );
NAND3_X1 U866 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(G27) );
NAND2_X1 U867 ( .A1(n1163), .A2(n1187), .ZN(n1186) );
NAND3_X1 U868 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NAND2_X1 U869 ( .A1(KEYINPUT23), .A2(n1191), .ZN(n1190) );
NAND2_X1 U870 ( .A1(KEYINPUT21), .A2(G125), .ZN(n1189) );
NAND2_X1 U871 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
INV_X1 U872 ( .A(KEYINPUT21), .ZN(n1193) );
NAND2_X1 U873 ( .A1(G125), .A2(n1194), .ZN(n1192) );
NAND2_X1 U874 ( .A1(KEYINPUT45), .A2(n1195), .ZN(n1194) );
INV_X1 U875 ( .A(n1196), .ZN(n1163) );
NAND4_X1 U876 ( .A1(n1196), .A2(n1191), .A3(G125), .A4(n1195), .ZN(n1185) );
INV_X1 U877 ( .A(KEYINPUT23), .ZN(n1195) );
INV_X1 U878 ( .A(KEYINPUT45), .ZN(n1191) );
NAND2_X1 U879 ( .A1(KEYINPUT23), .A2(n1197), .ZN(n1184) );
NAND2_X1 U880 ( .A1(G125), .A2(n1198), .ZN(n1197) );
NAND2_X1 U881 ( .A1(KEYINPUT45), .A2(n1196), .ZN(n1198) );
NAND4_X1 U882 ( .A1(n1170), .A2(n1039), .A3(n1024), .A4(n1026), .ZN(n1196) );
AND4_X1 U883 ( .A1(n1033), .A2(n1046), .A3(n1034), .A4(n1175), .ZN(n1170) );
NAND2_X1 U884 ( .A1(n1047), .A2(n1199), .ZN(n1175) );
NAND4_X1 U885 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1201), .ZN(n1199) );
INV_X1 U886 ( .A(G900), .ZN(n1201) );
XOR2_X1 U887 ( .A(n1142), .B(n1202), .Z(G24) );
NOR2_X1 U888 ( .A1(KEYINPUT2), .A2(n1203), .ZN(n1202) );
AND4_X1 U889 ( .A1(n1204), .A2(n1035), .A3(n1168), .A4(n1169), .ZN(n1142) );
AND2_X1 U890 ( .A1(n1033), .A2(n1205), .ZN(n1035) );
INV_X1 U891 ( .A(n1005), .ZN(n1033) );
XOR2_X1 U892 ( .A(G119), .B(n1145), .Z(G21) );
AND4_X1 U893 ( .A1(n1204), .A2(n1023), .A3(n1034), .A4(n1005), .ZN(n1145) );
XOR2_X1 U894 ( .A(G116), .B(n1141), .Z(G18) );
AND3_X1 U895 ( .A1(n1176), .A2(n1045), .A3(n1204), .ZN(n1141) );
AND2_X1 U896 ( .A1(n1009), .A2(n1168), .ZN(n1045) );
XOR2_X1 U897 ( .A(G113), .B(n1144), .Z(G15) );
AND3_X1 U898 ( .A1(n1046), .A2(n1176), .A3(n1204), .ZN(n1144) );
AND3_X1 U899 ( .A1(n1024), .A2(n1026), .A3(n1149), .ZN(n1204) );
INV_X1 U900 ( .A(n1147), .ZN(n1149) );
XNOR2_X1 U901 ( .A(n1206), .B(KEYINPUT61), .ZN(n1024) );
INV_X1 U902 ( .A(n1031), .ZN(n1176) );
NAND2_X1 U903 ( .A1(n1005), .A2(n1205), .ZN(n1031) );
XNOR2_X1 U904 ( .A(n1034), .B(KEYINPUT38), .ZN(n1205) );
NOR2_X1 U905 ( .A1(n1168), .A2(n1009), .ZN(n1046) );
INV_X1 U906 ( .A(n1169), .ZN(n1009) );
XOR2_X1 U907 ( .A(G110), .B(n1140), .Z(G12) );
NOR4_X1 U908 ( .A1(n1043), .A2(n1147), .A3(n1005), .A4(n1207), .ZN(n1140) );
INV_X1 U909 ( .A(n1034), .ZN(n1207) );
XOR2_X1 U910 ( .A(n1208), .B(n1209), .Z(n1034) );
XOR2_X1 U911 ( .A(KEYINPUT37), .B(n1210), .Z(n1209) );
NOR2_X1 U912 ( .A1(G902), .A2(n1013), .ZN(n1210) );
XOR2_X1 U913 ( .A(n1211), .B(n1212), .Z(n1013) );
XOR2_X1 U914 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U915 ( .A(n1215), .B(G119), .Z(n1214) );
NAND2_X1 U916 ( .A1(G221), .A2(n1216), .ZN(n1215) );
INV_X1 U917 ( .A(n1217), .ZN(n1216) );
XNOR2_X1 U918 ( .A(G128), .B(KEYINPUT54), .ZN(n1213) );
XOR2_X1 U919 ( .A(n1218), .B(n1219), .Z(n1211) );
XOR2_X1 U920 ( .A(n1129), .B(n1220), .Z(n1219) );
XNOR2_X1 U921 ( .A(G110), .B(n1066), .ZN(n1129) );
NAND2_X1 U922 ( .A1(KEYINPUT29), .A2(n1221), .ZN(n1208) );
INV_X1 U923 ( .A(n1012), .ZN(n1221) );
NAND2_X1 U924 ( .A1(G217), .A2(n1222), .ZN(n1012) );
XNOR2_X1 U925 ( .A(n1223), .B(G472), .ZN(n1005) );
NAND2_X1 U926 ( .A1(n1224), .A2(n1102), .ZN(n1223) );
XOR2_X1 U927 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U928 ( .A(n1116), .B(n1119), .Z(n1226) );
AND2_X1 U929 ( .A1(G210), .A2(n1227), .ZN(n1116) );
XOR2_X1 U930 ( .A(n1228), .B(n1229), .Z(n1225) );
XNOR2_X1 U931 ( .A(n1183), .B(n1230), .ZN(n1229) );
NOR2_X1 U932 ( .A1(KEYINPUT40), .A2(n1231), .ZN(n1230) );
XOR2_X1 U933 ( .A(n1111), .B(KEYINPUT25), .Z(n1231) );
XOR2_X1 U934 ( .A(n1232), .B(G119), .Z(n1111) );
INV_X1 U935 ( .A(G101), .ZN(n1183) );
NOR2_X1 U936 ( .A1(n1233), .A2(KEYINPUT49), .ZN(n1228) );
NAND2_X1 U937 ( .A1(n1039), .A2(n1182), .ZN(n1147) );
NAND2_X1 U938 ( .A1(n1047), .A2(n1234), .ZN(n1182) );
NAND4_X1 U939 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1072), .ZN(n1234) );
INV_X1 U940 ( .A(G898), .ZN(n1072) );
NAND3_X1 U941 ( .A1(n1200), .A2(n1000), .A3(G952), .ZN(n1047) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1200) );
NOR2_X1 U943 ( .A1(n1018), .A2(n1014), .ZN(n1039) );
AND2_X1 U944 ( .A1(G214), .A2(n1235), .ZN(n1014) );
INV_X1 U945 ( .A(n1177), .ZN(n1018) );
XOR2_X1 U946 ( .A(n1236), .B(n1136), .Z(n1177) );
NAND2_X1 U947 ( .A1(G210), .A2(n1235), .ZN(n1136) );
NAND2_X1 U948 ( .A1(n1102), .A2(n1237), .ZN(n1235) );
INV_X1 U949 ( .A(G237), .ZN(n1237) );
NAND2_X1 U950 ( .A1(n1238), .A2(n1102), .ZN(n1236) );
XNOR2_X1 U951 ( .A(KEYINPUT59), .B(n1239), .ZN(n1238) );
INV_X1 U952 ( .A(n1132), .ZN(n1239) );
XNOR2_X1 U953 ( .A(n1240), .B(n1241), .ZN(n1132) );
XOR2_X1 U954 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U955 ( .A(n1233), .B(G125), .ZN(n1243) );
INV_X1 U956 ( .A(n1118), .ZN(n1233) );
NAND2_X1 U957 ( .A1(n1244), .A2(n1245), .ZN(n1118) );
NAND2_X1 U958 ( .A1(G128), .A2(n1246), .ZN(n1245) );
XOR2_X1 U959 ( .A(KEYINPUT8), .B(n1247), .Z(n1244) );
NOR2_X1 U960 ( .A1(G128), .A2(n1246), .ZN(n1247) );
INV_X1 U961 ( .A(n1248), .ZN(n1246) );
NAND2_X1 U962 ( .A1(n1249), .A2(G224), .ZN(n1242) );
XNOR2_X1 U963 ( .A(G953), .B(KEYINPUT15), .ZN(n1249) );
XNOR2_X1 U964 ( .A(n1250), .B(n1088), .ZN(n1240) );
XNOR2_X1 U965 ( .A(G110), .B(G122), .ZN(n1088) );
XOR2_X1 U966 ( .A(n1084), .B(n1089), .Z(n1250) );
XNOR2_X1 U967 ( .A(n1232), .B(n1251), .ZN(n1089) );
NOR2_X1 U968 ( .A1(G119), .A2(KEYINPUT26), .ZN(n1251) );
XNOR2_X1 U969 ( .A(G113), .B(n1252), .ZN(n1232) );
XOR2_X1 U970 ( .A(KEYINPUT6), .B(G116), .Z(n1252) );
XNOR2_X1 U971 ( .A(n1130), .B(KEYINPUT4), .ZN(n1084) );
NAND2_X1 U972 ( .A1(n1023), .A2(n1148), .ZN(n1043) );
NOR2_X1 U973 ( .A1(n1206), .A2(n1015), .ZN(n1148) );
INV_X1 U974 ( .A(n1026), .ZN(n1015) );
NAND2_X1 U975 ( .A1(G221), .A2(n1222), .ZN(n1026) );
NAND2_X1 U976 ( .A1(n1253), .A2(G234), .ZN(n1222) );
XNOR2_X1 U977 ( .A(G902), .B(KEYINPUT43), .ZN(n1253) );
XNOR2_X1 U978 ( .A(G469), .B(n1254), .ZN(n1206) );
NOR2_X1 U979 ( .A1(KEYINPUT18), .A2(n1017), .ZN(n1254) );
NAND2_X1 U980 ( .A1(n1255), .A2(n1102), .ZN(n1017) );
XOR2_X1 U981 ( .A(n1256), .B(n1257), .Z(n1255) );
XNOR2_X1 U982 ( .A(n1123), .B(n1130), .ZN(n1257) );
XOR2_X1 U983 ( .A(G101), .B(n1258), .Z(n1130) );
XNOR2_X1 U984 ( .A(n996), .B(G104), .ZN(n1258) );
XNOR2_X1 U985 ( .A(n1259), .B(n1061), .ZN(n1123) );
XNOR2_X1 U986 ( .A(n1260), .B(n1261), .ZN(n1061) );
NOR2_X1 U987 ( .A1(KEYINPUT52), .A2(n1248), .ZN(n1261) );
XOR2_X1 U988 ( .A(G146), .B(n1166), .Z(n1248) );
INV_X1 U989 ( .A(G143), .ZN(n1166) );
NAND2_X1 U990 ( .A1(G227), .A2(n1000), .ZN(n1259) );
XOR2_X1 U991 ( .A(n1262), .B(n1263), .Z(n1256) );
XNOR2_X1 U992 ( .A(n1066), .B(n1264), .ZN(n1263) );
NOR2_X1 U993 ( .A1(G110), .A2(KEYINPUT31), .ZN(n1264) );
INV_X1 U994 ( .A(G140), .ZN(n1066) );
NAND2_X1 U995 ( .A1(KEYINPUT24), .A2(n1119), .ZN(n1262) );
XOR2_X1 U996 ( .A(n1265), .B(n1060), .Z(n1119) );
XOR2_X1 U997 ( .A(n1266), .B(n1220), .Z(n1060) );
XOR2_X1 U998 ( .A(G137), .B(KEYINPUT17), .Z(n1220) );
XNOR2_X1 U999 ( .A(G131), .B(G134), .ZN(n1266) );
XNOR2_X1 U1000 ( .A(KEYINPUT63), .B(KEYINPUT58), .ZN(n1265) );
NOR2_X1 U1001 ( .A1(n1169), .A2(n1168), .ZN(n1023) );
XNOR2_X1 U1002 ( .A(n1010), .B(KEYINPUT14), .ZN(n1168) );
XNOR2_X1 U1003 ( .A(n1267), .B(G478), .ZN(n1010) );
NAND2_X1 U1004 ( .A1(n1099), .A2(n1102), .ZN(n1267) );
INV_X1 U1005 ( .A(G902), .ZN(n1102) );
XOR2_X1 U1006 ( .A(n1268), .B(n1269), .Z(n1099) );
XNOR2_X1 U1007 ( .A(n996), .B(n1270), .ZN(n1269) );
XNOR2_X1 U1008 ( .A(n1203), .B(G116), .ZN(n1270) );
INV_X1 U1009 ( .A(G122), .ZN(n1203) );
INV_X1 U1010 ( .A(G107), .ZN(n996) );
XOR2_X1 U1011 ( .A(n1271), .B(n1272), .Z(n1268) );
NOR3_X1 U1012 ( .A1(n1273), .A2(KEYINPUT44), .A3(n1217), .ZN(n1272) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1000), .ZN(n1217) );
INV_X1 U1014 ( .A(G953), .ZN(n1000) );
INV_X1 U1015 ( .A(G217), .ZN(n1273) );
NAND3_X1 U1016 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1271) );
OR2_X1 U1017 ( .A1(n1277), .A2(KEYINPUT51), .ZN(n1276) );
OR3_X1 U1018 ( .A1(n1278), .A2(n1279), .A3(G134), .ZN(n1275) );
INV_X1 U1019 ( .A(KEYINPUT51), .ZN(n1278) );
NAND2_X1 U1020 ( .A1(G134), .A2(n1279), .ZN(n1274) );
NAND2_X1 U1021 ( .A1(KEYINPUT20), .A2(n1277), .ZN(n1279) );
XNOR2_X1 U1022 ( .A(G143), .B(n1260), .ZN(n1277) );
INV_X1 U1023 ( .A(G128), .ZN(n1260) );
XNOR2_X1 U1024 ( .A(n1280), .B(G475), .ZN(n1169) );
OR2_X1 U1025 ( .A1(n1105), .A2(G902), .ZN(n1280) );
XNOR2_X1 U1026 ( .A(n1281), .B(n1282), .ZN(n1105) );
XOR2_X1 U1027 ( .A(n1283), .B(n1218), .Z(n1282) );
XNOR2_X1 U1028 ( .A(G146), .B(G125), .ZN(n1218) );
NAND2_X1 U1029 ( .A1(KEYINPUT27), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1030 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U1031 ( .A(G131), .B(G143), .ZN(n1286) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1227), .ZN(n1285) );
NOR2_X1 U1033 ( .A1(G953), .A2(G237), .ZN(n1227) );
XOR2_X1 U1034 ( .A(n1287), .B(n1288), .Z(n1281) );
NOR2_X1 U1035 ( .A1(KEYINPUT28), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U1036 ( .A(G113), .B(G122), .ZN(n1289) );
XNOR2_X1 U1037 ( .A(G104), .B(n1290), .ZN(n1287) );
NOR2_X1 U1038 ( .A1(KEYINPUT55), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U1039 ( .A(G140), .B(KEYINPUT11), .ZN(n1291) );
endmodule


