//Key = 0111001011000101001101000000110001111001010010011000000010000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;

XNOR2_X1 U806 ( .A(G107), .B(n1135), .ZN(G9) );
NOR2_X1 U807 ( .A1(n1136), .A2(n1137), .ZN(G75) );
NOR4_X1 U808 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
NOR2_X1 U809 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
AND4_X1 U810 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1142) );
AND2_X1 U811 ( .A1(n1148), .A2(n1149), .ZN(n1144) );
XNOR2_X1 U812 ( .A(KEYINPUT18), .B(n1150), .ZN(n1139) );
NAND3_X1 U813 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1138) );
NAND2_X1 U814 ( .A1(n1148), .A2(n1154), .ZN(n1153) );
NAND2_X1 U815 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND3_X1 U816 ( .A1(n1157), .A2(n1158), .A3(n1146), .ZN(n1156) );
NAND2_X1 U817 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1161), .ZN(n1160) );
OR2_X1 U819 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U820 ( .A1(n1145), .A2(n1164), .ZN(n1159) );
NAND2_X1 U821 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U822 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND3_X1 U823 ( .A1(n1145), .A2(n1169), .A3(n1149), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U825 ( .A1(n1146), .A2(n1172), .ZN(n1171) );
NAND2_X1 U826 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U827 ( .A1(n1147), .A2(n1143), .ZN(n1174) );
INV_X1 U828 ( .A(KEYINPUT51), .ZN(n1143) );
NAND2_X1 U829 ( .A1(n1157), .A2(n1175), .ZN(n1170) );
NAND2_X1 U830 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U831 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
INV_X1 U832 ( .A(n1180), .ZN(n1148) );
NOR3_X1 U833 ( .A1(n1181), .A2(G953), .A3(G952), .ZN(n1136) );
INV_X1 U834 ( .A(n1151), .ZN(n1181) );
NAND4_X1 U835 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1151) );
NOR4_X1 U836 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
XOR2_X1 U837 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U838 ( .A(n1192), .B(n1193), .ZN(n1188) );
XOR2_X1 U839 ( .A(G469), .B(n1194), .Z(n1187) );
XNOR2_X1 U840 ( .A(KEYINPUT37), .B(n1195), .ZN(n1186) );
NOR3_X1 U841 ( .A1(n1178), .A2(n1167), .A3(n1196), .ZN(n1184) );
INV_X1 U842 ( .A(n1197), .ZN(n1196) );
XOR2_X1 U843 ( .A(n1198), .B(n1199), .Z(G72) );
XOR2_X1 U844 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U845 ( .A1(G953), .A2(n1202), .ZN(n1201) );
NAND2_X1 U846 ( .A1(G900), .A2(G227), .ZN(n1202) );
NAND2_X1 U847 ( .A1(n1203), .A2(n1204), .ZN(n1200) );
NAND2_X1 U848 ( .A1(G953), .A2(n1205), .ZN(n1204) );
XOR2_X1 U849 ( .A(n1206), .B(n1207), .Z(n1203) );
XOR2_X1 U850 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U851 ( .A(G131), .B(G134), .ZN(n1209) );
NAND2_X1 U852 ( .A1(KEYINPUT9), .A2(n1210), .ZN(n1208) );
XNOR2_X1 U853 ( .A(n1211), .B(n1212), .ZN(n1206) );
NOR2_X1 U854 ( .A1(n1213), .A2(G953), .ZN(n1198) );
XOR2_X1 U855 ( .A(n1214), .B(n1215), .Z(G69) );
NOR2_X1 U856 ( .A1(n1216), .A2(n1152), .ZN(n1215) );
AND2_X1 U857 ( .A1(G224), .A2(G898), .ZN(n1216) );
NAND3_X1 U858 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1214) );
OR2_X1 U859 ( .A1(n1220), .A2(KEYINPUT2), .ZN(n1219) );
NAND3_X1 U860 ( .A1(KEYINPUT2), .A2(n1220), .A3(n1221), .ZN(n1218) );
NOR2_X1 U861 ( .A1(G953), .A2(n1222), .ZN(n1220) );
NAND2_X1 U862 ( .A1(n1223), .A2(n1224), .ZN(n1217) );
INV_X1 U863 ( .A(n1221), .ZN(n1224) );
XNOR2_X1 U864 ( .A(n1225), .B(n1226), .ZN(n1221) );
XNOR2_X1 U865 ( .A(n1227), .B(n1228), .ZN(n1225) );
NAND2_X1 U866 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
NAND2_X1 U867 ( .A1(G898), .A2(G953), .ZN(n1230) );
NAND2_X1 U868 ( .A1(n1222), .A2(n1152), .ZN(n1229) );
NOR2_X1 U869 ( .A1(n1231), .A2(n1232), .ZN(G66) );
XOR2_X1 U870 ( .A(n1233), .B(n1234), .Z(n1232) );
NAND2_X1 U871 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
NOR2_X1 U872 ( .A1(n1231), .A2(n1237), .ZN(G63) );
NOR3_X1 U873 ( .A1(n1193), .A2(n1238), .A3(n1239), .ZN(n1237) );
AND3_X1 U874 ( .A1(n1240), .A2(G478), .A3(n1235), .ZN(n1239) );
NOR2_X1 U875 ( .A1(n1241), .A2(n1240), .ZN(n1238) );
NOR2_X1 U876 ( .A1(n1242), .A2(n1192), .ZN(n1241) );
NOR2_X1 U877 ( .A1(n1150), .A2(n1141), .ZN(n1242) );
NOR2_X1 U878 ( .A1(n1231), .A2(n1243), .ZN(G60) );
XOR2_X1 U879 ( .A(n1244), .B(n1245), .Z(n1243) );
AND2_X1 U880 ( .A1(G475), .A2(n1235), .ZN(n1245) );
NAND2_X1 U881 ( .A1(KEYINPUT21), .A2(n1246), .ZN(n1244) );
XOR2_X1 U882 ( .A(KEYINPUT40), .B(n1247), .Z(n1246) );
XNOR2_X1 U883 ( .A(G104), .B(n1248), .ZN(G6) );
NOR3_X1 U884 ( .A1(n1231), .A2(n1249), .A3(n1250), .ZN(G57) );
NOR2_X1 U885 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U886 ( .A(n1253), .ZN(n1252) );
NOR2_X1 U887 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
AND2_X1 U888 ( .A1(KEYINPUT57), .A2(n1256), .ZN(n1255) );
NOR3_X1 U889 ( .A1(KEYINPUT57), .A2(KEYINPUT17), .A3(n1256), .ZN(n1254) );
NOR2_X1 U890 ( .A1(n1257), .A2(n1253), .ZN(n1249) );
XNOR2_X1 U891 ( .A(n1258), .B(n1259), .ZN(n1253) );
XOR2_X1 U892 ( .A(n1260), .B(n1261), .Z(n1258) );
NOR3_X1 U893 ( .A1(n1262), .A2(KEYINPUT31), .A3(n1263), .ZN(n1261) );
NAND2_X1 U894 ( .A1(n1264), .A2(n1265), .ZN(n1260) );
NAND3_X1 U895 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1265) );
NAND2_X1 U896 ( .A1(KEYINPUT42), .A2(n1269), .ZN(n1267) );
NAND2_X1 U897 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
INV_X1 U898 ( .A(KEYINPUT42), .ZN(n1271) );
NAND2_X1 U899 ( .A1(n1272), .A2(n1270), .ZN(n1264) );
NAND2_X1 U900 ( .A1(KEYINPUT35), .A2(n1269), .ZN(n1270) );
NOR2_X1 U901 ( .A1(KEYINPUT17), .A2(n1256), .ZN(n1257) );
XNOR2_X1 U902 ( .A(n1273), .B(n1274), .ZN(n1256) );
NOR2_X1 U903 ( .A1(KEYINPUT60), .A2(n1275), .ZN(n1274) );
NOR2_X1 U904 ( .A1(n1231), .A2(n1276), .ZN(G54) );
XNOR2_X1 U905 ( .A(n1277), .B(n1278), .ZN(n1276) );
XOR2_X1 U906 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U907 ( .A1(KEYINPUT30), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U908 ( .A(n1269), .B(n1282), .ZN(n1281) );
NOR2_X1 U909 ( .A1(KEYINPUT12), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U910 ( .A(n1284), .B(n1285), .ZN(n1283) );
XNOR2_X1 U911 ( .A(KEYINPUT15), .B(n1212), .ZN(n1285) );
NAND2_X1 U912 ( .A1(n1235), .A2(G469), .ZN(n1279) );
NOR2_X1 U913 ( .A1(n1231), .A2(n1286), .ZN(G51) );
XOR2_X1 U914 ( .A(n1287), .B(n1288), .Z(n1286) );
XNOR2_X1 U915 ( .A(KEYINPUT6), .B(n1289), .ZN(n1288) );
XOR2_X1 U916 ( .A(n1290), .B(n1291), .Z(n1287) );
NAND3_X1 U917 ( .A1(n1235), .A2(n1190), .A3(KEYINPUT61), .ZN(n1290) );
INV_X1 U918 ( .A(n1262), .ZN(n1235) );
NAND2_X1 U919 ( .A1(G902), .A2(n1292), .ZN(n1262) );
NAND2_X1 U920 ( .A1(n1213), .A2(n1222), .ZN(n1292) );
INV_X1 U921 ( .A(n1150), .ZN(n1222) );
NAND4_X1 U922 ( .A1(n1293), .A2(n1248), .A3(n1294), .A4(n1295), .ZN(n1150) );
AND4_X1 U923 ( .A1(n1135), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1295) );
NAND3_X1 U924 ( .A1(n1157), .A2(n1299), .A3(n1163), .ZN(n1135) );
AND2_X1 U925 ( .A1(n1300), .A2(n1301), .ZN(n1294) );
NAND3_X1 U926 ( .A1(n1157), .A2(n1299), .A3(n1162), .ZN(n1248) );
NAND2_X1 U927 ( .A1(n1302), .A2(n1303), .ZN(n1293) );
XOR2_X1 U928 ( .A(n1304), .B(KEYINPUT28), .Z(n1302) );
INV_X1 U929 ( .A(n1141), .ZN(n1213) );
NAND4_X1 U930 ( .A1(n1305), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(n1141) );
AND4_X1 U931 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1308) );
OR2_X1 U932 ( .A1(n1313), .A2(n1176), .ZN(n1307) );
NAND3_X1 U933 ( .A1(n1314), .A2(n1315), .A3(n1147), .ZN(n1305) );
NAND2_X1 U934 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND3_X1 U935 ( .A1(n1318), .A2(n1319), .A3(n1303), .ZN(n1317) );
NAND2_X1 U936 ( .A1(n1162), .A2(n1146), .ZN(n1316) );
NOR2_X1 U937 ( .A1(n1152), .A2(G952), .ZN(n1231) );
NAND3_X1 U938 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(G48) );
NAND2_X1 U939 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND3_X1 U940 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1324) );
NAND2_X1 U941 ( .A1(KEYINPUT59), .A2(n1328), .ZN(n1327) );
OR2_X1 U942 ( .A1(n1329), .A2(KEYINPUT47), .ZN(n1326) );
NAND2_X1 U943 ( .A1(KEYINPUT47), .A2(n1330), .ZN(n1325) );
NAND2_X1 U944 ( .A1(G146), .A2(n1331), .ZN(n1330) );
NAND2_X1 U945 ( .A1(KEYINPUT23), .A2(n1332), .ZN(n1331) );
INV_X1 U946 ( .A(n1306), .ZN(n1323) );
NAND4_X1 U947 ( .A1(n1306), .A2(n1328), .A3(G146), .A4(n1332), .ZN(n1321) );
INV_X1 U948 ( .A(KEYINPUT59), .ZN(n1332) );
INV_X1 U949 ( .A(KEYINPUT23), .ZN(n1328) );
NAND2_X1 U950 ( .A1(KEYINPUT59), .A2(n1333), .ZN(n1320) );
NAND2_X1 U951 ( .A1(G146), .A2(n1334), .ZN(n1333) );
NAND2_X1 U952 ( .A1(KEYINPUT23), .A2(n1306), .ZN(n1334) );
NAND3_X1 U953 ( .A1(n1335), .A2(n1303), .A3(n1162), .ZN(n1306) );
XNOR2_X1 U954 ( .A(G143), .B(n1336), .ZN(G45) );
NAND4_X1 U955 ( .A1(n1337), .A2(n1338), .A3(n1147), .A4(n1339), .ZN(n1336) );
NOR3_X1 U956 ( .A1(n1176), .A2(n1340), .A3(n1182), .ZN(n1339) );
OR2_X1 U957 ( .A1(n1314), .A2(KEYINPUT22), .ZN(n1338) );
NAND2_X1 U958 ( .A1(KEYINPUT22), .A2(n1341), .ZN(n1337) );
NAND2_X1 U959 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U960 ( .A(G140), .B(n1344), .Z(G42) );
NOR2_X1 U961 ( .A1(KEYINPUT58), .A2(n1312), .ZN(n1344) );
NAND4_X1 U962 ( .A1(n1162), .A2(n1345), .A3(n1146), .A4(n1314), .ZN(n1312) );
XNOR2_X1 U963 ( .A(G137), .B(n1311), .ZN(G39) );
NAND3_X1 U964 ( .A1(n1146), .A2(n1335), .A3(n1145), .ZN(n1311) );
XNOR2_X1 U965 ( .A(G134), .B(n1310), .ZN(G36) );
NAND4_X1 U966 ( .A1(n1147), .A2(n1146), .A3(n1314), .A4(n1163), .ZN(n1310) );
XNOR2_X1 U967 ( .A(G131), .B(n1346), .ZN(G33) );
NAND4_X1 U968 ( .A1(n1162), .A2(n1147), .A3(n1314), .A4(n1347), .ZN(n1346) );
XOR2_X1 U969 ( .A(KEYINPUT20), .B(n1146), .Z(n1347) );
AND2_X1 U970 ( .A1(n1348), .A2(n1179), .ZN(n1146) );
XNOR2_X1 U971 ( .A(KEYINPUT16), .B(n1178), .ZN(n1348) );
XNOR2_X1 U972 ( .A(G128), .B(n1309), .ZN(G30) );
NAND3_X1 U973 ( .A1(n1163), .A2(n1303), .A3(n1335), .ZN(n1309) );
AND3_X1 U974 ( .A1(n1349), .A2(n1350), .A3(n1314), .ZN(n1335) );
NOR2_X1 U975 ( .A1(n1165), .A2(n1342), .ZN(n1314) );
INV_X1 U976 ( .A(n1351), .ZN(n1342) );
INV_X1 U977 ( .A(n1343), .ZN(n1165) );
XNOR2_X1 U978 ( .A(G101), .B(n1301), .ZN(G3) );
NAND3_X1 U979 ( .A1(n1147), .A2(n1299), .A3(n1145), .ZN(n1301) );
AND3_X1 U980 ( .A1(n1343), .A2(n1352), .A3(n1303), .ZN(n1299) );
XOR2_X1 U981 ( .A(G125), .B(n1353), .Z(G27) );
NOR2_X1 U982 ( .A1(n1354), .A2(n1313), .ZN(n1353) );
NAND4_X1 U983 ( .A1(n1149), .A2(n1162), .A3(n1345), .A4(n1351), .ZN(n1313) );
NAND2_X1 U984 ( .A1(n1180), .A2(n1355), .ZN(n1351) );
NAND4_X1 U985 ( .A1(G953), .A2(G902), .A3(n1356), .A4(n1205), .ZN(n1355) );
INV_X1 U986 ( .A(G900), .ZN(n1205) );
XNOR2_X1 U987 ( .A(n1303), .B(KEYINPUT54), .ZN(n1354) );
NAND2_X1 U988 ( .A1(n1357), .A2(n1358), .ZN(G24) );
NAND2_X1 U989 ( .A1(G122), .A2(n1359), .ZN(n1358) );
NAND2_X1 U990 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U991 ( .A1(KEYINPUT55), .A2(n1362), .ZN(n1361) );
INV_X1 U992 ( .A(n1363), .ZN(n1362) );
XOR2_X1 U993 ( .A(n1300), .B(KEYINPUT44), .Z(n1360) );
OR3_X1 U994 ( .A1(n1363), .A2(KEYINPUT55), .A3(G122), .ZN(n1357) );
XNOR2_X1 U995 ( .A(n1300), .B(KEYINPUT19), .ZN(n1363) );
NAND4_X1 U996 ( .A1(n1364), .A2(n1157), .A3(n1318), .A4(n1319), .ZN(n1300) );
NOR2_X1 U997 ( .A1(n1365), .A2(n1350), .ZN(n1157) );
XNOR2_X1 U998 ( .A(G119), .B(n1298), .ZN(G21) );
NAND4_X1 U999 ( .A1(n1364), .A2(n1145), .A3(n1349), .A4(n1350), .ZN(n1298) );
INV_X1 U1000 ( .A(n1366), .ZN(n1350) );
XNOR2_X1 U1001 ( .A(G116), .B(n1297), .ZN(G18) );
NAND3_X1 U1002 ( .A1(n1147), .A2(n1163), .A3(n1364), .ZN(n1297) );
NOR2_X1 U1003 ( .A1(n1318), .A2(n1340), .ZN(n1163) );
INV_X1 U1004 ( .A(n1319), .ZN(n1340) );
XNOR2_X1 U1005 ( .A(G113), .B(n1296), .ZN(G15) );
NAND3_X1 U1006 ( .A1(n1162), .A2(n1147), .A3(n1364), .ZN(n1296) );
AND3_X1 U1007 ( .A1(n1303), .A2(n1352), .A3(n1149), .ZN(n1364) );
AND2_X1 U1008 ( .A1(n1367), .A2(n1168), .ZN(n1149) );
XNOR2_X1 U1009 ( .A(KEYINPUT45), .B(n1167), .ZN(n1367) );
NOR2_X1 U1010 ( .A1(n1365), .A2(n1366), .ZN(n1147) );
NOR2_X1 U1011 ( .A1(n1319), .A2(n1182), .ZN(n1162) );
INV_X1 U1012 ( .A(n1318), .ZN(n1182) );
XNOR2_X1 U1013 ( .A(n1228), .B(n1368), .ZN(G12) );
NOR2_X1 U1014 ( .A1(n1176), .A2(n1304), .ZN(n1368) );
NAND4_X1 U1015 ( .A1(n1345), .A2(n1145), .A3(n1343), .A4(n1352), .ZN(n1304) );
NAND2_X1 U1016 ( .A1(n1180), .A2(n1369), .ZN(n1352) );
NAND4_X1 U1017 ( .A1(G953), .A2(G902), .A3(n1356), .A4(n1370), .ZN(n1369) );
INV_X1 U1018 ( .A(G898), .ZN(n1370) );
NAND3_X1 U1019 ( .A1(n1356), .A2(n1152), .A3(G952), .ZN(n1180) );
NAND2_X1 U1020 ( .A1(G237), .A2(G234), .ZN(n1356) );
NOR2_X1 U1021 ( .A1(n1371), .A2(n1168), .ZN(n1343) );
XOR2_X1 U1022 ( .A(G469), .B(n1372), .Z(n1168) );
NOR2_X1 U1023 ( .A1(n1194), .A2(KEYINPUT7), .ZN(n1372) );
AND2_X1 U1024 ( .A1(n1373), .A2(n1374), .ZN(n1194) );
XOR2_X1 U1025 ( .A(n1375), .B(n1376), .Z(n1373) );
XNOR2_X1 U1026 ( .A(n1377), .B(n1378), .ZN(n1376) );
INV_X1 U1027 ( .A(n1277), .ZN(n1378) );
XNOR2_X1 U1028 ( .A(n1379), .B(n1380), .ZN(n1277) );
XNOR2_X1 U1029 ( .A(G140), .B(n1228), .ZN(n1380) );
NAND2_X1 U1030 ( .A1(G227), .A2(n1152), .ZN(n1379) );
NOR3_X1 U1031 ( .A1(n1381), .A2(n1382), .A3(n1383), .ZN(n1377) );
NOR2_X1 U1032 ( .A1(n1384), .A2(n1284), .ZN(n1383) );
NOR2_X1 U1033 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
XOR2_X1 U1034 ( .A(KEYINPUT52), .B(n1387), .Z(n1385) );
NOR3_X1 U1035 ( .A1(n1388), .A2(n1387), .A3(n1386), .ZN(n1382) );
INV_X1 U1036 ( .A(n1284), .ZN(n1388) );
NAND2_X1 U1037 ( .A1(n1389), .A2(n1390), .ZN(n1284) );
NAND2_X1 U1038 ( .A1(G101), .A2(n1391), .ZN(n1390) );
NAND2_X1 U1039 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND3_X1 U1040 ( .A1(n1392), .A2(n1393), .A3(n1275), .ZN(n1389) );
NAND2_X1 U1041 ( .A1(G104), .A2(n1394), .ZN(n1393) );
XNOR2_X1 U1042 ( .A(KEYINPUT48), .B(n1395), .ZN(n1392) );
NAND2_X1 U1043 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
XNOR2_X1 U1044 ( .A(KEYINPUT43), .B(n1394), .ZN(n1396) );
AND2_X1 U1045 ( .A1(n1386), .A2(n1387), .ZN(n1381) );
XNOR2_X1 U1046 ( .A(n1212), .B(KEYINPUT33), .ZN(n1387) );
NAND2_X1 U1047 ( .A1(n1398), .A2(n1399), .ZN(n1212) );
OR2_X1 U1048 ( .A1(n1400), .A2(KEYINPUT11), .ZN(n1399) );
NAND2_X1 U1049 ( .A1(KEYINPUT11), .A2(n1401), .ZN(n1398) );
NAND2_X1 U1050 ( .A1(n1402), .A2(n1403), .ZN(n1401) );
OR2_X1 U1051 ( .A1(n1404), .A2(G128), .ZN(n1403) );
INV_X1 U1052 ( .A(KEYINPUT29), .ZN(n1386) );
XNOR2_X1 U1053 ( .A(n1269), .B(KEYINPUT62), .ZN(n1375) );
XOR2_X1 U1054 ( .A(KEYINPUT45), .B(n1167), .Z(n1371) );
AND2_X1 U1055 ( .A1(G221), .A2(n1405), .ZN(n1167) );
NOR2_X1 U1056 ( .A1(n1319), .A2(n1318), .ZN(n1145) );
XNOR2_X1 U1057 ( .A(n1406), .B(G475), .ZN(n1318) );
NAND2_X1 U1058 ( .A1(n1247), .A2(n1374), .ZN(n1406) );
XNOR2_X1 U1059 ( .A(n1407), .B(n1408), .ZN(n1247) );
XOR2_X1 U1060 ( .A(n1409), .B(n1410), .Z(n1408) );
XNOR2_X1 U1061 ( .A(n1411), .B(G131), .ZN(n1410) );
XNOR2_X1 U1062 ( .A(KEYINPUT49), .B(n1329), .ZN(n1409) );
XOR2_X1 U1063 ( .A(n1412), .B(n1226), .Z(n1407) );
XOR2_X1 U1064 ( .A(G122), .B(n1413), .Z(n1226) );
XOR2_X1 U1065 ( .A(n1414), .B(n1415), .Z(n1412) );
NOR2_X1 U1066 ( .A1(KEYINPUT38), .A2(n1211), .ZN(n1415) );
NAND3_X1 U1067 ( .A1(n1416), .A2(n1152), .A3(G214), .ZN(n1414) );
NAND3_X1 U1068 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1319) );
OR2_X1 U1069 ( .A1(n1193), .A2(KEYINPUT56), .ZN(n1419) );
NAND3_X1 U1070 ( .A1(KEYINPUT56), .A2(n1193), .A3(n1192), .ZN(n1418) );
INV_X1 U1071 ( .A(G478), .ZN(n1192) );
NAND2_X1 U1072 ( .A1(G478), .A2(n1420), .ZN(n1417) );
NAND2_X1 U1073 ( .A1(KEYINPUT56), .A2(n1421), .ZN(n1420) );
XOR2_X1 U1074 ( .A(KEYINPUT25), .B(n1193), .Z(n1421) );
NOR2_X1 U1075 ( .A1(n1240), .A2(G902), .ZN(n1193) );
XNOR2_X1 U1076 ( .A(n1422), .B(n1423), .ZN(n1240) );
XOR2_X1 U1077 ( .A(n1424), .B(n1425), .Z(n1423) );
XNOR2_X1 U1078 ( .A(n1426), .B(G122), .ZN(n1425) );
XNOR2_X1 U1079 ( .A(KEYINPUT5), .B(n1427), .ZN(n1424) );
INV_X1 U1080 ( .A(G134), .ZN(n1427) );
XOR2_X1 U1081 ( .A(n1428), .B(n1429), .Z(n1422) );
XNOR2_X1 U1082 ( .A(G116), .B(n1394), .ZN(n1429) );
XOR2_X1 U1083 ( .A(n1430), .B(n1431), .Z(n1428) );
NOR2_X1 U1084 ( .A1(G143), .A2(KEYINPUT0), .ZN(n1431) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1432), .ZN(n1430) );
INV_X1 U1086 ( .A(n1173), .ZN(n1345) );
NAND2_X1 U1087 ( .A1(n1366), .A2(n1349), .ZN(n1173) );
XNOR2_X1 U1088 ( .A(n1365), .B(KEYINPUT13), .ZN(n1349) );
NAND2_X1 U1089 ( .A1(n1195), .A2(n1197), .ZN(n1365) );
NAND3_X1 U1090 ( .A1(n1433), .A2(n1374), .A3(n1234), .ZN(n1197) );
NAND2_X1 U1091 ( .A1(n1236), .A2(n1434), .ZN(n1195) );
NAND2_X1 U1092 ( .A1(n1234), .A2(n1374), .ZN(n1434) );
XOR2_X1 U1093 ( .A(n1435), .B(n1436), .Z(n1234) );
XNOR2_X1 U1094 ( .A(G137), .B(n1437), .ZN(n1436) );
NAND2_X1 U1095 ( .A1(G221), .A2(n1432), .ZN(n1437) );
AND2_X1 U1096 ( .A1(G234), .A2(n1152), .ZN(n1432) );
NAND2_X1 U1097 ( .A1(n1438), .A2(n1439), .ZN(n1435) );
NAND2_X1 U1098 ( .A1(n1440), .A2(n1441), .ZN(n1439) );
XOR2_X1 U1099 ( .A(KEYINPUT3), .B(n1442), .Z(n1441) );
XNOR2_X1 U1100 ( .A(n1443), .B(n1444), .ZN(n1440) );
NAND2_X1 U1101 ( .A1(n1445), .A2(n1446), .ZN(n1438) );
XNOR2_X1 U1102 ( .A(n1211), .B(n1443), .ZN(n1446) );
XNOR2_X1 U1103 ( .A(n1447), .B(KEYINPUT24), .ZN(n1443) );
NAND2_X1 U1104 ( .A1(KEYINPUT8), .A2(G146), .ZN(n1447) );
INV_X1 U1105 ( .A(n1444), .ZN(n1211) );
XOR2_X1 U1106 ( .A(G125), .B(G140), .Z(n1444) );
XNOR2_X1 U1107 ( .A(n1442), .B(KEYINPUT34), .ZN(n1445) );
XNOR2_X1 U1108 ( .A(n1448), .B(n1449), .ZN(n1442) );
NOR2_X1 U1109 ( .A1(KEYINPUT50), .A2(G119), .ZN(n1449) );
XNOR2_X1 U1110 ( .A(G110), .B(G128), .ZN(n1448) );
INV_X1 U1111 ( .A(n1433), .ZN(n1236) );
NAND2_X1 U1112 ( .A1(G217), .A2(n1405), .ZN(n1433) );
NAND2_X1 U1113 ( .A1(G234), .A2(n1374), .ZN(n1405) );
XOR2_X1 U1114 ( .A(n1183), .B(KEYINPUT63), .Z(n1366) );
XNOR2_X1 U1115 ( .A(n1450), .B(n1263), .ZN(n1183) );
INV_X1 U1116 ( .A(G472), .ZN(n1263) );
NAND2_X1 U1117 ( .A1(n1374), .A2(n1451), .ZN(n1450) );
NAND2_X1 U1118 ( .A1(n1452), .A2(n1453), .ZN(n1451) );
NAND3_X1 U1119 ( .A1(n1454), .A2(n1273), .A3(n1455), .ZN(n1453) );
XNOR2_X1 U1120 ( .A(KEYINPUT53), .B(n1456), .ZN(n1455) );
XOR2_X1 U1121 ( .A(KEYINPUT39), .B(n1457), .Z(n1454) );
NAND3_X1 U1122 ( .A1(n1458), .A2(n1459), .A3(n1460), .ZN(n1452) );
NAND2_X1 U1123 ( .A1(n1461), .A2(n1273), .ZN(n1460) );
NAND2_X1 U1124 ( .A1(n1462), .A2(n1456), .ZN(n1461) );
INV_X1 U1125 ( .A(n1463), .ZN(n1456) );
XNOR2_X1 U1126 ( .A(KEYINPUT39), .B(n1457), .ZN(n1462) );
OR3_X1 U1127 ( .A1(n1273), .A2(n1464), .A3(n1463), .ZN(n1459) );
NAND3_X1 U1128 ( .A1(n1416), .A2(n1152), .A3(G210), .ZN(n1273) );
NAND2_X1 U1129 ( .A1(n1464), .A2(n1463), .ZN(n1458) );
NAND2_X1 U1130 ( .A1(n1465), .A2(n1466), .ZN(n1463) );
NAND2_X1 U1131 ( .A1(n1467), .A2(n1259), .ZN(n1466) );
XOR2_X1 U1132 ( .A(KEYINPUT36), .B(n1468), .Z(n1465) );
NOR2_X1 U1133 ( .A1(n1467), .A2(n1259), .ZN(n1468) );
XNOR2_X1 U1134 ( .A(G113), .B(n1469), .ZN(n1259) );
AND2_X1 U1135 ( .A1(n1470), .A2(n1268), .ZN(n1467) );
NAND2_X1 U1136 ( .A1(n1272), .A2(n1269), .ZN(n1268) );
INV_X1 U1137 ( .A(n1471), .ZN(n1269) );
INV_X1 U1138 ( .A(n1400), .ZN(n1272) );
XOR2_X1 U1139 ( .A(n1472), .B(KEYINPUT32), .Z(n1470) );
NAND2_X1 U1140 ( .A1(n1400), .A2(n1471), .ZN(n1472) );
NAND2_X1 U1141 ( .A1(n1473), .A2(n1474), .ZN(n1471) );
NAND2_X1 U1142 ( .A1(G131), .A2(n1475), .ZN(n1474) );
XOR2_X1 U1143 ( .A(n1476), .B(KEYINPUT46), .Z(n1473) );
OR2_X1 U1144 ( .A1(n1475), .A2(G131), .ZN(n1476) );
XNOR2_X1 U1145 ( .A(G134), .B(n1210), .ZN(n1475) );
INV_X1 U1146 ( .A(G137), .ZN(n1210) );
NAND2_X1 U1147 ( .A1(n1457), .A2(n1477), .ZN(n1464) );
INV_X1 U1148 ( .A(KEYINPUT53), .ZN(n1477) );
XNOR2_X1 U1149 ( .A(n1275), .B(KEYINPUT41), .ZN(n1457) );
INV_X1 U1150 ( .A(G101), .ZN(n1275) );
INV_X1 U1151 ( .A(n1303), .ZN(n1176) );
NOR2_X1 U1152 ( .A1(n1478), .A2(n1179), .ZN(n1303) );
XOR2_X1 U1153 ( .A(n1190), .B(n1479), .Z(n1179) );
NOR2_X1 U1154 ( .A1(n1191), .A2(KEYINPUT27), .ZN(n1479) );
AND2_X1 U1155 ( .A1(n1480), .A2(n1374), .ZN(n1191) );
XNOR2_X1 U1156 ( .A(n1291), .B(n1481), .ZN(n1480) );
NOR2_X1 U1157 ( .A1(KEYINPUT14), .A2(n1289), .ZN(n1481) );
NAND2_X1 U1158 ( .A1(G224), .A2(n1152), .ZN(n1289) );
INV_X1 U1159 ( .A(G953), .ZN(n1152) );
XNOR2_X1 U1160 ( .A(n1482), .B(n1483), .ZN(n1291) );
XOR2_X1 U1161 ( .A(n1484), .B(n1485), .Z(n1483) );
XOR2_X1 U1162 ( .A(KEYINPUT1), .B(G125), .Z(n1485) );
NOR2_X1 U1163 ( .A1(KEYINPUT26), .A2(n1486), .ZN(n1484) );
XNOR2_X1 U1164 ( .A(G110), .B(G122), .ZN(n1486) );
XOR2_X1 U1165 ( .A(n1487), .B(n1413), .Z(n1482) );
XNOR2_X1 U1166 ( .A(G113), .B(n1397), .ZN(n1413) );
INV_X1 U1167 ( .A(G104), .ZN(n1397) );
XNOR2_X1 U1168 ( .A(n1227), .B(n1400), .ZN(n1487) );
NAND3_X1 U1169 ( .A1(n1488), .A2(n1489), .A3(n1402), .ZN(n1400) );
NAND2_X1 U1170 ( .A1(n1404), .A2(G128), .ZN(n1402) );
NOR2_X1 U1171 ( .A1(n1411), .A2(G146), .ZN(n1404) );
NAND3_X1 U1172 ( .A1(n1426), .A2(n1411), .A3(n1329), .ZN(n1489) );
INV_X1 U1173 ( .A(G146), .ZN(n1329) );
INV_X1 U1174 ( .A(G128), .ZN(n1426) );
NAND2_X1 U1175 ( .A1(n1490), .A2(G146), .ZN(n1488) );
XNOR2_X1 U1176 ( .A(n1411), .B(G128), .ZN(n1490) );
INV_X1 U1177 ( .A(G143), .ZN(n1411) );
XOR2_X1 U1178 ( .A(n1491), .B(n1492), .Z(n1227) );
XNOR2_X1 U1179 ( .A(KEYINPUT10), .B(n1394), .ZN(n1492) );
INV_X1 U1180 ( .A(G107), .ZN(n1394) );
XNOR2_X1 U1181 ( .A(G101), .B(n1493), .ZN(n1491) );
NOR2_X1 U1182 ( .A1(KEYINPUT4), .A2(n1469), .ZN(n1493) );
XNOR2_X1 U1183 ( .A(G116), .B(G119), .ZN(n1469) );
AND2_X1 U1184 ( .A1(G210), .A2(n1494), .ZN(n1190) );
XOR2_X1 U1185 ( .A(KEYINPUT16), .B(n1178), .Z(n1478) );
AND2_X1 U1186 ( .A1(G214), .A2(n1494), .ZN(n1178) );
NAND2_X1 U1187 ( .A1(n1374), .A2(n1416), .ZN(n1494) );
INV_X1 U1188 ( .A(G237), .ZN(n1416) );
INV_X1 U1189 ( .A(G902), .ZN(n1374) );
INV_X1 U1190 ( .A(G110), .ZN(n1228) );
endmodule


