//Key = 1110010110111110000010110011101010001000010000101000110011011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306;

XNOR2_X1 U711 ( .A(n985), .B(n986), .ZN(G9) );
INV_X1 U712 ( .A(G107), .ZN(n985) );
NOR2_X1 U713 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U714 ( .A1(G953), .A2(n989), .A3(n990), .A4(n991), .ZN(n988) );
NOR2_X1 U715 ( .A1(n992), .A2(n993), .ZN(n990) );
NOR2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR3_X1 U717 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NOR2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR3_X1 U719 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n999) );
INV_X1 U720 ( .A(KEYINPUT23), .ZN(n1001) );
NOR3_X1 U721 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n994) );
NOR2_X1 U722 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR3_X1 U723 ( .A1(n998), .A2(n1008), .A3(n1009), .ZN(n1007) );
NOR3_X1 U724 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1009) );
NOR2_X1 U725 ( .A1(n1013), .A2(n1014), .ZN(n1008) );
NOR2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NOR2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U728 ( .A1(n1002), .A2(n996), .ZN(n1006) );
INV_X1 U729 ( .A(n1019), .ZN(n996) );
NOR4_X1 U730 ( .A1(n1020), .A2(n1004), .A3(n1021), .A4(n1022), .ZN(n1002) );
NOR2_X1 U731 ( .A1(n998), .A2(KEYINPUT23), .ZN(n1020) );
INV_X1 U732 ( .A(n1023), .ZN(n998) );
INV_X1 U733 ( .A(n1024), .ZN(n1003) );
NOR3_X1 U734 ( .A1(n989), .A2(G953), .A3(G952), .ZN(n987) );
AND4_X1 U735 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n989) );
NOR4_X1 U736 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NOR3_X1 U737 ( .A1(n1004), .A2(n1033), .A3(n1034), .ZN(n1027) );
NAND2_X1 U738 ( .A1(n1035), .A2(n1036), .ZN(n1026) );
XOR2_X1 U739 ( .A(n1037), .B(KEYINPUT17), .Z(n1035) );
XNOR2_X1 U740 ( .A(KEYINPUT59), .B(n1038), .ZN(n1025) );
XOR2_X1 U741 ( .A(n1039), .B(n1040), .Z(G72) );
NOR2_X1 U742 ( .A1(KEYINPUT15), .A2(n1041), .ZN(n1040) );
XOR2_X1 U743 ( .A(n1042), .B(n1043), .Z(n1041) );
NAND2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U745 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XOR2_X1 U746 ( .A(n1048), .B(KEYINPUT39), .Z(n1046) );
XNOR2_X1 U747 ( .A(KEYINPUT46), .B(n1049), .ZN(n1044) );
NAND2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1042) );
NAND2_X1 U749 ( .A1(G953), .A2(n1052), .ZN(n1051) );
XOR2_X1 U750 ( .A(n1053), .B(n1054), .Z(n1050) );
XNOR2_X1 U751 ( .A(n1055), .B(KEYINPUT52), .ZN(n1054) );
NAND2_X1 U752 ( .A1(KEYINPUT48), .A2(n1056), .ZN(n1055) );
XNOR2_X1 U753 ( .A(n1057), .B(n1058), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1059), .B(n1060), .ZN(n1058) );
NAND3_X1 U755 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1059) );
OR2_X1 U756 ( .A1(n1064), .A2(KEYINPUT36), .ZN(n1063) );
NAND3_X1 U757 ( .A1(KEYINPUT36), .A2(n1064), .A3(G137), .ZN(n1062) );
NAND2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1067), .A2(KEYINPUT36), .ZN(n1065) );
XNOR2_X1 U760 ( .A(n1068), .B(n1064), .ZN(n1067) );
XNOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT51), .ZN(n1068) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1039) );
NAND2_X1 U763 ( .A1(G900), .A2(G227), .ZN(n1070) );
INV_X1 U764 ( .A(n1071), .ZN(n1069) );
XOR2_X1 U765 ( .A(n1072), .B(n1073), .Z(G69) );
NOR2_X1 U766 ( .A1(n1074), .A2(n1071), .ZN(n1073) );
XOR2_X1 U767 ( .A(G953), .B(KEYINPUT56), .Z(n1071) );
NOR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1072) );
OR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U771 ( .A(n1081), .B(KEYINPUT31), .Z(n1077) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1079), .ZN(n1081) );
NAND3_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1079) );
NAND2_X1 U774 ( .A1(G953), .A2(n1076), .ZN(n1084) );
OR2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1087), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U778 ( .A1(KEYINPUT53), .A2(n1086), .ZN(n1089) );
OR2_X1 U779 ( .A1(KEYINPUT19), .A2(n1090), .ZN(n1086) );
OR2_X1 U780 ( .A1(n1090), .A2(KEYINPUT53), .ZN(n1088) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U782 ( .A(G107), .B(KEYINPUT50), .ZN(n1091) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1085) );
XNOR2_X1 U784 ( .A(G110), .B(KEYINPUT11), .ZN(n1093) );
NOR2_X1 U785 ( .A1(G953), .A2(n1095), .ZN(n1080) );
NOR3_X1 U786 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(G66) );
AND2_X1 U787 ( .A1(KEYINPUT57), .A2(n1099), .ZN(n1098) );
NOR3_X1 U788 ( .A1(KEYINPUT57), .A2(n1049), .A3(n1100), .ZN(n1097) );
INV_X1 U789 ( .A(G952), .ZN(n1100) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(G63) );
XNOR2_X1 U793 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1109), .A2(n1104), .ZN(n1108) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1049), .ZN(n1105) );
XNOR2_X1 U796 ( .A(G952), .B(KEYINPUT5), .ZN(n1110) );
NOR2_X1 U797 ( .A1(n1099), .A2(n1111), .ZN(G60) );
XOR2_X1 U798 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1104), .ZN(n1112) );
XOR2_X1 U800 ( .A(G104), .B(n1115), .Z(G6) );
NOR2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(G57) );
XOR2_X1 U802 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
OR2_X1 U804 ( .A1(n1122), .A2(KEYINPUT32), .ZN(n1121) );
XOR2_X1 U805 ( .A(n1123), .B(n1124), .Z(n1120) );
NOR2_X1 U806 ( .A1(n1125), .A2(n1104), .ZN(n1124) );
NAND2_X1 U807 ( .A1(KEYINPUT32), .A2(n1122), .ZN(n1123) );
NAND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U810 ( .A(KEYINPUT0), .B(n1130), .Z(n1126) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1128), .ZN(n1130) );
XNOR2_X1 U812 ( .A(n1131), .B(n1132), .ZN(n1128) );
NOR2_X1 U813 ( .A1(G952), .A2(n1133), .ZN(n1116) );
XNOR2_X1 U814 ( .A(G953), .B(KEYINPUT16), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1099), .A2(n1134), .ZN(G54) );
XOR2_X1 U816 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U817 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U818 ( .A1(KEYINPUT20), .A2(n1139), .ZN(n1138) );
NAND3_X1 U819 ( .A1(n1140), .A2(n991), .A3(G469), .ZN(n1137) );
XNOR2_X1 U820 ( .A(KEYINPUT24), .B(n1141), .ZN(n1140) );
NOR2_X1 U821 ( .A1(n1099), .A2(n1142), .ZN(G51) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1104), .ZN(n1144) );
NAND2_X1 U824 ( .A1(G902), .A2(n991), .ZN(n1104) );
NAND3_X1 U825 ( .A1(n1095), .A2(n1048), .A3(n1047), .ZN(n991) );
AND4_X1 U826 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1047) );
NOR4_X1 U827 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
NAND2_X1 U828 ( .A1(n1154), .A2(n1155), .ZN(n1148) );
XOR2_X1 U829 ( .A(KEYINPUT62), .B(n1156), .Z(n1155) );
AND4_X1 U830 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1095) );
NOR4_X1 U831 ( .A1(n1115), .A2(n1161), .A3(n986), .A4(n1162), .ZN(n1160) );
NOR2_X1 U832 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U833 ( .A(KEYINPUT22), .B(n1165), .Z(n1164) );
INV_X1 U834 ( .A(n1000), .ZN(n1163) );
AND3_X1 U835 ( .A1(n1012), .A2(n1023), .A3(n1166), .ZN(n986) );
AND3_X1 U836 ( .A1(n1166), .A2(n1023), .A3(n1011), .ZN(n1115) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1168), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1170), .ZN(n1143) );
XOR2_X1 U839 ( .A(KEYINPUT34), .B(n1171), .Z(n1170) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
AND2_X1 U841 ( .A1(n1173), .A2(n1172), .ZN(n1169) );
XNOR2_X1 U842 ( .A(n1174), .B(n1175), .ZN(n1173) );
NAND3_X1 U843 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
OR2_X1 U844 ( .A1(n1132), .A2(KEYINPUT14), .ZN(n1178) );
NAND3_X1 U845 ( .A1(KEYINPUT14), .A2(n1132), .A3(G125), .ZN(n1177) );
NAND2_X1 U846 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1181), .A2(KEYINPUT14), .ZN(n1179) );
XNOR2_X1 U848 ( .A(n1182), .B(KEYINPUT58), .ZN(n1181) );
NOR2_X1 U849 ( .A1(n1049), .A2(G952), .ZN(n1099) );
XNOR2_X1 U850 ( .A(G146), .B(n1146), .ZN(G48) );
NAND3_X1 U851 ( .A1(n1156), .A2(n1011), .A3(n1183), .ZN(n1146) );
XOR2_X1 U852 ( .A(n1048), .B(n1184), .Z(G45) );
NAND2_X1 U853 ( .A1(KEYINPUT12), .A2(G143), .ZN(n1184) );
NAND4_X1 U854 ( .A1(n1183), .A2(n1021), .A3(n1032), .A4(n1185), .ZN(n1048) );
XOR2_X1 U855 ( .A(n1147), .B(n1186), .Z(G42) );
NAND2_X1 U856 ( .A1(KEYINPUT41), .A2(G140), .ZN(n1186) );
NAND3_X1 U857 ( .A1(n1022), .A2(n1011), .A3(n1187), .ZN(n1147) );
XNOR2_X1 U858 ( .A(G137), .B(n1188), .ZN(G39) );
NAND2_X1 U859 ( .A1(n1154), .A2(n1156), .ZN(n1188) );
AND2_X1 U860 ( .A1(n1189), .A2(n1187), .ZN(n1154) );
XNOR2_X1 U861 ( .A(G134), .B(n1190), .ZN(G36) );
NOR2_X1 U862 ( .A1(n1152), .A2(KEYINPUT9), .ZN(n1190) );
AND3_X1 U863 ( .A1(n1021), .A2(n1012), .A3(n1187), .ZN(n1152) );
XOR2_X1 U864 ( .A(n1151), .B(n1191), .Z(G33) );
NOR2_X1 U865 ( .A1(KEYINPUT43), .A2(n1060), .ZN(n1191) );
AND2_X1 U866 ( .A1(n1192), .A2(n1187), .ZN(n1151) );
AND3_X1 U867 ( .A1(n1024), .A2(n1193), .A3(n1194), .ZN(n1187) );
NOR3_X1 U868 ( .A1(n1004), .A2(n1017), .A3(n1033), .ZN(n1194) );
NAND3_X1 U869 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(G30) );
NAND2_X1 U870 ( .A1(KEYINPUT47), .A2(n1198), .ZN(n1197) );
NAND3_X1 U871 ( .A1(n1153), .A2(n1199), .A3(n1200), .ZN(n1196) );
INV_X1 U872 ( .A(n1198), .ZN(n1153) );
NAND2_X1 U873 ( .A1(G128), .A2(n1201), .ZN(n1195) );
NAND2_X1 U874 ( .A1(n1202), .A2(n1199), .ZN(n1201) );
INV_X1 U875 ( .A(KEYINPUT47), .ZN(n1199) );
XNOR2_X1 U876 ( .A(KEYINPUT29), .B(n1198), .ZN(n1202) );
NAND3_X1 U877 ( .A1(n1156), .A2(n1012), .A3(n1183), .ZN(n1198) );
AND4_X1 U878 ( .A1(n1000), .A2(n1193), .A3(n1018), .A4(n1203), .ZN(n1183) );
XNOR2_X1 U879 ( .A(G101), .B(n1157), .ZN(G3) );
NAND3_X1 U880 ( .A1(n1021), .A2(n1166), .A3(n1189), .ZN(n1157) );
XNOR2_X1 U881 ( .A(G125), .B(n1204), .ZN(G27) );
NOR2_X1 U882 ( .A1(n1150), .A2(KEYINPUT40), .ZN(n1204) );
AND4_X1 U883 ( .A1(n1000), .A2(n1193), .A3(n1013), .A4(n1205), .ZN(n1150) );
AND2_X1 U884 ( .A1(n1011), .A2(n1022), .ZN(n1205) );
NAND2_X1 U885 ( .A1(n993), .A2(n1206), .ZN(n1193) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1207), .A4(n1052), .ZN(n1206) );
INV_X1 U887 ( .A(G900), .ZN(n1052) );
XNOR2_X1 U888 ( .A(G122), .B(n1158), .ZN(G24) );
NAND4_X1 U889 ( .A1(n1208), .A2(n1023), .A3(n1032), .A4(n1185), .ZN(n1158) );
NOR2_X1 U890 ( .A1(n1031), .A2(n1209), .ZN(n1023) );
XNOR2_X1 U891 ( .A(G119), .B(n1210), .ZN(G21) );
NAND3_X1 U892 ( .A1(n1165), .A2(n1000), .A3(KEYINPUT7), .ZN(n1210) );
AND3_X1 U893 ( .A1(n1156), .A2(n1211), .A3(n1019), .ZN(n1165) );
NOR2_X1 U894 ( .A1(n1016), .A2(n1010), .ZN(n1019) );
INV_X1 U895 ( .A(n1189), .ZN(n1016) );
NOR2_X1 U896 ( .A1(n1212), .A2(n1213), .ZN(n1156) );
XNOR2_X1 U897 ( .A(G116), .B(n1214), .ZN(G18) );
NOR2_X1 U898 ( .A1(n1168), .A2(KEYINPUT55), .ZN(n1214) );
AND3_X1 U899 ( .A1(n1021), .A2(n1012), .A3(n1208), .ZN(n1168) );
NOR2_X1 U900 ( .A1(n1185), .A2(n1215), .ZN(n1012) );
INV_X1 U901 ( .A(n1032), .ZN(n1215) );
XNOR2_X1 U902 ( .A(n1216), .B(n1217), .ZN(G15) );
NAND2_X1 U903 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND4_X1 U904 ( .A1(n1220), .A2(n1010), .A3(n1192), .A4(n1221), .ZN(n1219) );
INV_X1 U905 ( .A(KEYINPUT26), .ZN(n1221) );
INV_X1 U906 ( .A(n1013), .ZN(n1010) );
NAND2_X1 U907 ( .A1(n1161), .A2(KEYINPUT26), .ZN(n1218) );
AND2_X1 U908 ( .A1(n1208), .A2(n1192), .ZN(n1161) );
AND2_X1 U909 ( .A1(n1021), .A2(n1011), .ZN(n1192) );
NOR2_X1 U910 ( .A1(n1032), .A2(n1038), .ZN(n1011) );
INV_X1 U911 ( .A(n1185), .ZN(n1038) );
NOR2_X1 U912 ( .A1(n1209), .A2(n1213), .ZN(n1021) );
INV_X1 U913 ( .A(n1031), .ZN(n1213) );
INV_X1 U914 ( .A(n1212), .ZN(n1209) );
AND2_X1 U915 ( .A1(n1013), .A2(n1220), .ZN(n1208) );
NOR2_X1 U916 ( .A1(n1203), .A2(n1033), .ZN(n1013) );
INV_X1 U917 ( .A(n1018), .ZN(n1033) );
XOR2_X1 U918 ( .A(G110), .B(n1167), .Z(G12) );
AND3_X1 U919 ( .A1(n1022), .A2(n1166), .A3(n1189), .ZN(n1167) );
NOR2_X1 U920 ( .A1(n1032), .A2(n1185), .ZN(n1189) );
XOR2_X1 U921 ( .A(n1222), .B(n1114), .Z(n1185) );
INV_X1 U922 ( .A(G475), .ZN(n1114) );
OR2_X1 U923 ( .A1(n1113), .A2(G902), .ZN(n1222) );
XNOR2_X1 U924 ( .A(n1223), .B(n1224), .ZN(n1113) );
XOR2_X1 U925 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U926 ( .A(n1217), .B(G104), .ZN(n1226) );
XNOR2_X1 U927 ( .A(n1227), .B(G131), .ZN(n1225) );
XNOR2_X1 U928 ( .A(n1228), .B(n1094), .ZN(n1223) );
INV_X1 U929 ( .A(n1229), .ZN(n1094) );
XOR2_X1 U930 ( .A(n1230), .B(n1231), .Z(n1228) );
AND2_X1 U931 ( .A1(G214), .A2(n1232), .ZN(n1231) );
NAND2_X1 U932 ( .A1(n1233), .A2(KEYINPUT63), .ZN(n1230) );
XOR2_X1 U933 ( .A(n1053), .B(G146), .Z(n1233) );
XNOR2_X1 U934 ( .A(G125), .B(n1234), .ZN(n1053) );
XOR2_X1 U935 ( .A(n1235), .B(n1109), .Z(n1032) );
INV_X1 U936 ( .A(G478), .ZN(n1109) );
NAND2_X1 U937 ( .A1(n1107), .A2(n1141), .ZN(n1235) );
XNOR2_X1 U938 ( .A(n1236), .B(n1237), .ZN(n1107) );
XNOR2_X1 U939 ( .A(n1238), .B(n1229), .ZN(n1237) );
NAND3_X1 U940 ( .A1(G217), .A2(n1239), .A3(KEYINPUT27), .ZN(n1238) );
XOR2_X1 U941 ( .A(n1240), .B(n1241), .Z(n1236) );
XNOR2_X1 U942 ( .A(n1242), .B(G107), .ZN(n1241) );
NAND2_X1 U943 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
OR2_X1 U944 ( .A1(n1245), .A2(n1064), .ZN(n1244) );
XOR2_X1 U945 ( .A(n1246), .B(KEYINPUT44), .Z(n1243) );
NAND2_X1 U946 ( .A1(n1245), .A2(n1064), .ZN(n1246) );
XOR2_X1 U947 ( .A(n1247), .B(n1200), .Z(n1245) );
NAND2_X1 U948 ( .A1(KEYINPUT28), .A2(n1227), .ZN(n1247) );
INV_X1 U949 ( .A(G143), .ZN(n1227) );
AND3_X1 U950 ( .A1(n1018), .A2(n1203), .A3(n1220), .ZN(n1166) );
AND2_X1 U951 ( .A1(n1000), .A2(n1211), .ZN(n1220) );
NAND2_X1 U952 ( .A1(n993), .A2(n1248), .ZN(n1211) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1207), .A4(n1076), .ZN(n1248) );
INV_X1 U954 ( .A(G898), .ZN(n1076) );
NAND3_X1 U955 ( .A1(n1207), .A2(n1049), .A3(G952), .ZN(n993) );
NAND2_X1 U956 ( .A1(G237), .A2(G234), .ZN(n1207) );
NOR2_X1 U957 ( .A1(n1024), .A2(n1004), .ZN(n1000) );
AND2_X1 U958 ( .A1(G214), .A2(n1249), .ZN(n1004) );
XOR2_X1 U959 ( .A(n1030), .B(KEYINPUT10), .Z(n1024) );
XOR2_X1 U960 ( .A(n1250), .B(n1145), .Z(n1030) );
NAND2_X1 U961 ( .A1(G210), .A2(n1249), .ZN(n1145) );
NAND2_X1 U962 ( .A1(n1251), .A2(n1141), .ZN(n1249) );
INV_X1 U963 ( .A(G237), .ZN(n1251) );
NAND2_X1 U964 ( .A1(n1252), .A2(n1141), .ZN(n1250) );
XOR2_X1 U965 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U966 ( .A(n1180), .B(n1175), .ZN(n1254) );
NOR2_X1 U967 ( .A1(n1075), .A2(G953), .ZN(n1175) );
INV_X1 U968 ( .A(G224), .ZN(n1075) );
XNOR2_X1 U969 ( .A(n1132), .B(n1172), .ZN(n1253) );
XOR2_X1 U970 ( .A(n1255), .B(n1092), .Z(n1172) );
XNOR2_X1 U971 ( .A(n1256), .B(n1257), .ZN(n1092) );
XNOR2_X1 U972 ( .A(n1258), .B(n1259), .ZN(n1257) );
NOR2_X1 U973 ( .A1(G104), .A2(KEYINPUT3), .ZN(n1259) );
NAND2_X1 U974 ( .A1(KEYINPUT30), .A2(n1260), .ZN(n1258) );
XNOR2_X1 U975 ( .A(n1242), .B(n1261), .ZN(n1260) );
XNOR2_X1 U976 ( .A(KEYINPUT33), .B(n1262), .ZN(n1261) );
INV_X1 U977 ( .A(G116), .ZN(n1242) );
XNOR2_X1 U978 ( .A(G101), .B(G113), .ZN(n1256) );
XNOR2_X1 U979 ( .A(n1263), .B(n1229), .ZN(n1255) );
XOR2_X1 U980 ( .A(G122), .B(KEYINPUT45), .Z(n1229) );
INV_X1 U981 ( .A(n1182), .ZN(n1132) );
INV_X1 U982 ( .A(n1017), .ZN(n1203) );
NOR2_X1 U983 ( .A1(n1264), .A2(n1034), .ZN(n1017) );
NOR2_X1 U984 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
AND2_X1 U985 ( .A1(n1037), .A2(n1036), .ZN(n1264) );
NAND2_X1 U986 ( .A1(n1265), .A2(n1141), .ZN(n1036) );
XNOR2_X1 U987 ( .A(n1135), .B(n1139), .ZN(n1265) );
XNOR2_X1 U988 ( .A(n1234), .B(KEYINPUT21), .ZN(n1139) );
XNOR2_X1 U989 ( .A(n1266), .B(n1267), .ZN(n1135) );
XOR2_X1 U990 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U991 ( .A(G104), .B(n1270), .ZN(n1269) );
AND2_X1 U992 ( .A1(n1049), .A2(G227), .ZN(n1270) );
NAND2_X1 U993 ( .A1(KEYINPUT60), .A2(n1271), .ZN(n1268) );
XNOR2_X1 U994 ( .A(n1272), .B(n1273), .ZN(n1266) );
INV_X1 U995 ( .A(n1057), .ZN(n1273) );
XOR2_X1 U996 ( .A(G128), .B(n1274), .Z(n1057) );
NOR2_X1 U997 ( .A1(KEYINPUT6), .A2(n1275), .ZN(n1274) );
XNOR2_X1 U998 ( .A(G143), .B(G146), .ZN(n1275) );
XOR2_X1 U999 ( .A(n1131), .B(n1263), .Z(n1272) );
XOR2_X1 U1000 ( .A(G107), .B(G110), .Z(n1263) );
XNOR2_X1 U1001 ( .A(G469), .B(KEYINPUT1), .ZN(n1037) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1276), .ZN(n1018) );
NOR2_X1 U1003 ( .A1(n1212), .A2(n1031), .ZN(n1022) );
XOR2_X1 U1004 ( .A(n1277), .B(n1125), .Z(n1031) );
INV_X1 U1005 ( .A(G472), .ZN(n1125) );
NAND2_X1 U1006 ( .A1(n1278), .A2(n1141), .ZN(n1277) );
XOR2_X1 U1007 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U1008 ( .A(n1119), .B(n1182), .ZN(n1280) );
XOR2_X1 U1009 ( .A(G143), .B(n1281), .Z(n1182) );
XOR2_X1 U1010 ( .A(n1282), .B(n1271), .Z(n1119) );
INV_X1 U1011 ( .A(G101), .ZN(n1271) );
NAND2_X1 U1012 ( .A1(n1232), .A2(G210), .ZN(n1282) );
NOR2_X1 U1013 ( .A1(G953), .A2(G237), .ZN(n1232) );
XOR2_X1 U1014 ( .A(n1283), .B(n1284), .Z(n1279) );
NOR2_X1 U1015 ( .A1(KEYINPUT25), .A2(n1131), .ZN(n1284) );
XOR2_X1 U1016 ( .A(n1285), .B(n1286), .Z(n1131) );
XNOR2_X1 U1017 ( .A(KEYINPUT18), .B(n1066), .ZN(n1286) );
XNOR2_X1 U1018 ( .A(n1287), .B(n1064), .ZN(n1285) );
INV_X1 U1019 ( .A(G134), .ZN(n1064) );
NAND2_X1 U1020 ( .A1(KEYINPUT61), .A2(n1060), .ZN(n1287) );
INV_X1 U1021 ( .A(G131), .ZN(n1060) );
XNOR2_X1 U1022 ( .A(n1129), .B(KEYINPUT2), .ZN(n1283) );
AND2_X1 U1023 ( .A1(n1288), .A2(n1289), .ZN(n1129) );
NAND2_X1 U1024 ( .A1(n1290), .A2(n1217), .ZN(n1289) );
INV_X1 U1025 ( .A(G113), .ZN(n1217) );
XOR2_X1 U1026 ( .A(n1291), .B(KEYINPUT8), .Z(n1290) );
XOR2_X1 U1027 ( .A(n1292), .B(KEYINPUT35), .Z(n1288) );
NAND2_X1 U1028 ( .A1(G113), .A2(n1291), .ZN(n1292) );
NAND2_X1 U1029 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
OR2_X1 U1030 ( .A1(n1295), .A2(n1262), .ZN(n1294) );
XOR2_X1 U1031 ( .A(n1296), .B(KEYINPUT4), .Z(n1293) );
NAND2_X1 U1032 ( .A1(n1295), .A2(n1262), .ZN(n1296) );
INV_X1 U1033 ( .A(G119), .ZN(n1262) );
XOR2_X1 U1034 ( .A(G116), .B(KEYINPUT49), .Z(n1295) );
XOR2_X1 U1035 ( .A(n1029), .B(KEYINPUT13), .Z(n1212) );
XOR2_X1 U1036 ( .A(n1297), .B(n1103), .Z(n1029) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1276), .ZN(n1103) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1141), .ZN(n1276) );
NAND2_X1 U1039 ( .A1(n1101), .A2(n1141), .ZN(n1297) );
INV_X1 U1040 ( .A(G902), .ZN(n1141) );
XNOR2_X1 U1041 ( .A(n1298), .B(n1299), .ZN(n1101) );
XNOR2_X1 U1042 ( .A(n1066), .B(n1300), .ZN(n1299) );
NOR2_X1 U1043 ( .A1(KEYINPUT38), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1044 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1045 ( .A(n1304), .B(n1281), .Z(n1303) );
XNOR2_X1 U1046 ( .A(n1200), .B(G146), .ZN(n1281) );
INV_X1 U1047 ( .A(G128), .ZN(n1200) );
NOR2_X1 U1048 ( .A1(KEYINPUT42), .A2(n1305), .ZN(n1304) );
INV_X1 U1049 ( .A(n1234), .ZN(n1305) );
XOR2_X1 U1050 ( .A(G140), .B(KEYINPUT37), .Z(n1234) );
XNOR2_X1 U1051 ( .A(G110), .B(n1306), .ZN(n1302) );
XNOR2_X1 U1052 ( .A(n1180), .B(G119), .ZN(n1306) );
INV_X1 U1053 ( .A(G125), .ZN(n1180) );
INV_X1 U1054 ( .A(G137), .ZN(n1066) );
NAND2_X1 U1055 ( .A1(n1239), .A2(G221), .ZN(n1298) );
AND2_X1 U1056 ( .A1(G234), .A2(n1049), .ZN(n1239) );
INV_X1 U1057 ( .A(G953), .ZN(n1049) );
endmodule


