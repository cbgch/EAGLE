//Key = 0101001100111111011011111101011010010000011111101011000110011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352;

XNOR2_X1 U727 ( .A(G107), .B(n1021), .ZN(G9) );
NAND2_X1 U728 ( .A1(KEYINPUT13), .A2(n1022), .ZN(n1021) );
NOR2_X1 U729 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR4_X1 U730 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
INV_X1 U731 ( .A(G952), .ZN(n1027) );
XOR2_X1 U732 ( .A(KEYINPUT31), .B(n1029), .Z(n1026) );
NOR4_X1 U733 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
NAND2_X1 U734 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NAND3_X1 U735 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1025) );
NAND2_X1 U736 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U737 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U738 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NAND2_X1 U739 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NAND2_X1 U740 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
OR2_X1 U741 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U742 ( .A1(n1052), .A2(n1053), .ZN(n1046) );
NAND3_X1 U743 ( .A1(n1053), .A2(n1054), .A3(n1048), .ZN(n1041) );
NAND3_X1 U744 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U745 ( .A1(n1045), .A2(n1058), .ZN(n1057) );
NAND3_X1 U746 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1056) );
XNOR2_X1 U747 ( .A(KEYINPUT0), .B(n1032), .ZN(n1059) );
INV_X1 U748 ( .A(n1045), .ZN(n1032) );
NAND2_X1 U749 ( .A1(n1043), .A2(n1062), .ZN(n1055) );
NAND2_X1 U750 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U751 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U752 ( .A(n1033), .ZN(n1039) );
NOR3_X1 U753 ( .A1(n1067), .A2(G953), .A3(n1068), .ZN(n1023) );
INV_X1 U754 ( .A(n1036), .ZN(n1068) );
NAND4_X1 U755 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1036) );
NOR4_X1 U756 ( .A1(n1065), .A2(n1061), .A3(n1073), .A4(n1074), .ZN(n1072) );
NOR2_X1 U757 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
AND2_X1 U758 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U759 ( .A1(n1079), .A2(n1080), .ZN(n1071) );
XNOR2_X1 U760 ( .A(n1081), .B(n1082), .ZN(n1080) );
XNOR2_X1 U761 ( .A(G475), .B(n1083), .ZN(n1079) );
XOR2_X1 U762 ( .A(n1084), .B(G469), .Z(n1070) );
XOR2_X1 U763 ( .A(n1085), .B(KEYINPUT61), .Z(n1069) );
XNOR2_X1 U764 ( .A(G952), .B(KEYINPUT60), .ZN(n1067) );
XOR2_X1 U765 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U766 ( .A1(n1088), .A2(G953), .ZN(n1087) );
NOR2_X1 U767 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
AND2_X1 U768 ( .A1(n1037), .A2(n1091), .ZN(n1090) );
NOR3_X1 U769 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1089) );
NOR2_X1 U770 ( .A1(n1091), .A2(n1095), .ZN(n1094) );
NOR2_X1 U771 ( .A1(G227), .A2(n1096), .ZN(n1093) );
NOR2_X1 U772 ( .A1(n1091), .A2(n1037), .ZN(n1096) );
XOR2_X1 U773 ( .A(n1097), .B(n1098), .Z(n1091) );
XNOR2_X1 U774 ( .A(G131), .B(n1099), .ZN(n1098) );
NAND2_X1 U775 ( .A1(KEYINPUT62), .A2(n1100), .ZN(n1099) );
XOR2_X1 U776 ( .A(n1101), .B(n1102), .Z(n1097) );
XOR2_X1 U777 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U778 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U779 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U780 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U781 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U782 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U783 ( .A(n1111), .B(n1112), .Z(n1108) );
XNOR2_X1 U784 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND2_X1 U785 ( .A1(KEYINPUT6), .A2(n1115), .ZN(n1114) );
NAND2_X1 U786 ( .A1(KEYINPUT20), .A2(n1116), .ZN(n1113) );
NOR2_X1 U787 ( .A1(n1117), .A2(G953), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U789 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND3_X1 U790 ( .A1(G902), .A2(n1122), .A3(G217), .ZN(n1120) );
XNOR2_X1 U791 ( .A(KEYINPUT44), .B(n1028), .ZN(n1122) );
NOR3_X1 U792 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(G63) );
NOR3_X1 U793 ( .A1(n1126), .A2(G953), .A3(G952), .ZN(n1125) );
AND2_X1 U794 ( .A1(n1126), .A2(n1118), .ZN(n1124) );
INV_X1 U795 ( .A(KEYINPUT40), .ZN(n1126) );
NOR3_X1 U796 ( .A1(n1082), .A2(n1127), .A3(n1128), .ZN(n1123) );
AND3_X1 U797 ( .A1(n1129), .A2(G478), .A3(n1130), .ZN(n1128) );
NOR2_X1 U798 ( .A1(n1131), .A2(n1129), .ZN(n1127) );
NOR2_X1 U799 ( .A1(n1132), .A2(n1081), .ZN(n1131) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1133), .ZN(G60) );
NOR3_X1 U801 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR3_X1 U802 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR2_X1 U803 ( .A1(n1140), .A2(n1141), .ZN(n1135) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1138), .ZN(n1141) );
XNOR2_X1 U805 ( .A(G104), .B(n1142), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1118), .A2(n1143), .ZN(G57) );
XNOR2_X1 U807 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U808 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U809 ( .A(n1148), .B(KEYINPUT27), .Z(n1147) );
NAND2_X1 U810 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U811 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
AND2_X1 U812 ( .A1(n1130), .A2(G472), .ZN(n1149) );
NOR2_X1 U813 ( .A1(n1118), .A2(n1151), .ZN(G54) );
XOR2_X1 U814 ( .A(n1152), .B(n1153), .Z(n1151) );
AND2_X1 U815 ( .A1(G469), .A2(n1130), .ZN(n1153) );
NAND2_X1 U816 ( .A1(n1154), .A2(KEYINPUT30), .ZN(n1152) );
XOR2_X1 U817 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U818 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U819 ( .A(G140), .B(G110), .Z(n1158) );
XNOR2_X1 U820 ( .A(n1159), .B(n1160), .ZN(n1155) );
NOR2_X1 U821 ( .A1(KEYINPUT47), .A2(n1161), .ZN(n1160) );
XOR2_X1 U822 ( .A(n1162), .B(KEYINPUT54), .Z(n1161) );
NOR2_X1 U823 ( .A1(n1118), .A2(n1163), .ZN(G51) );
XOR2_X1 U824 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U825 ( .A1(n1076), .A2(n1139), .ZN(n1165) );
INV_X1 U826 ( .A(n1130), .ZN(n1139) );
NOR2_X1 U827 ( .A1(n1077), .A2(n1132), .ZN(n1130) );
INV_X1 U828 ( .A(n1028), .ZN(n1132) );
NAND2_X1 U829 ( .A1(n1117), .A2(n1088), .ZN(n1028) );
AND4_X1 U830 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1088) );
AND4_X1 U831 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NOR2_X1 U832 ( .A1(n1174), .A2(n1175), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
INV_X1 U834 ( .A(KEYINPUT11), .ZN(n1176) );
NOR2_X1 U835 ( .A1(KEYINPUT11), .A2(n1178), .ZN(n1174) );
NAND4_X1 U836 ( .A1(n1179), .A2(n1043), .A3(n1180), .A4(n1063), .ZN(n1178) );
INV_X1 U837 ( .A(n1181), .ZN(n1063) );
NAND2_X1 U838 ( .A1(n1182), .A2(n1183), .ZN(n1166) );
NAND2_X1 U839 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
AND2_X1 U840 ( .A1(n1186), .A2(n1187), .ZN(n1117) );
AND4_X1 U841 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR4_X1 U842 ( .A1(n1192), .A2(n1193), .A3(n1022), .A4(n1194), .ZN(n1186) );
AND3_X1 U843 ( .A1(n1050), .A2(n1048), .A3(n1195), .ZN(n1022) );
INV_X1 U844 ( .A(n1142), .ZN(n1193) );
NAND3_X1 U845 ( .A1(n1195), .A2(n1048), .A3(n1051), .ZN(n1142) );
INV_X1 U846 ( .A(n1196), .ZN(n1192) );
NOR2_X1 U847 ( .A1(n1197), .A2(n1198), .ZN(n1164) );
XOR2_X1 U848 ( .A(n1199), .B(KEYINPUT23), .Z(n1198) );
NAND2_X1 U849 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NOR2_X1 U850 ( .A1(n1200), .A2(n1201), .ZN(n1197) );
XOR2_X1 U851 ( .A(n1202), .B(n1203), .Z(n1200) );
XOR2_X1 U852 ( .A(KEYINPUT50), .B(KEYINPUT33), .Z(n1203) );
XNOR2_X1 U853 ( .A(n1204), .B(n1205), .ZN(n1202) );
NOR2_X1 U854 ( .A1(n1037), .A2(G952), .ZN(n1118) );
XNOR2_X1 U855 ( .A(G146), .B(n1170), .ZN(G48) );
NAND3_X1 U856 ( .A1(n1051), .A2(n1206), .A3(n1207), .ZN(n1170) );
XNOR2_X1 U857 ( .A(G143), .B(n1167), .ZN(G45) );
OR4_X1 U858 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1206), .ZN(n1167) );
XNOR2_X1 U859 ( .A(G140), .B(n1173), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1045), .A2(n1182), .A3(n1179), .ZN(n1173) );
XNOR2_X1 U861 ( .A(G137), .B(n1211), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
INV_X1 U863 ( .A(n1184), .ZN(n1214) );
NAND3_X1 U864 ( .A1(n1035), .A2(n1215), .A3(n1045), .ZN(n1184) );
OR2_X1 U865 ( .A1(n1182), .A2(KEYINPUT63), .ZN(n1213) );
NAND2_X1 U866 ( .A1(KEYINPUT63), .A2(n1216), .ZN(n1212) );
XNOR2_X1 U867 ( .A(G134), .B(n1217), .ZN(G36) );
NAND3_X1 U868 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
INV_X1 U869 ( .A(n1185), .ZN(n1220) );
NAND3_X1 U870 ( .A1(n1052), .A2(n1050), .A3(n1045), .ZN(n1185) );
OR2_X1 U871 ( .A1(n1182), .A2(KEYINPUT2), .ZN(n1219) );
NAND2_X1 U872 ( .A1(KEYINPUT2), .A2(n1216), .ZN(n1218) );
NAND2_X1 U873 ( .A1(n1221), .A2(n1058), .ZN(n1216) );
INV_X1 U874 ( .A(n1180), .ZN(n1221) );
XNOR2_X1 U875 ( .A(G131), .B(n1172), .ZN(G33) );
NAND4_X1 U876 ( .A1(n1045), .A2(n1182), .A3(n1052), .A4(n1051), .ZN(n1172) );
NOR2_X1 U877 ( .A1(n1222), .A2(n1065), .ZN(n1045) );
XOR2_X1 U878 ( .A(G128), .B(n1223), .Z(G30) );
NOR2_X1 U879 ( .A1(KEYINPUT19), .A2(n1171), .ZN(n1223) );
NAND3_X1 U880 ( .A1(n1050), .A2(n1206), .A3(n1207), .ZN(n1171) );
INV_X1 U881 ( .A(n1209), .ZN(n1207) );
NAND3_X1 U882 ( .A1(n1181), .A2(n1215), .A3(n1182), .ZN(n1209) );
AND2_X1 U883 ( .A1(n1058), .A2(n1180), .ZN(n1182) );
XNOR2_X1 U884 ( .A(G101), .B(n1196), .ZN(G3) );
NAND3_X1 U885 ( .A1(n1195), .A2(n1053), .A3(n1052), .ZN(n1196) );
XNOR2_X1 U886 ( .A(G125), .B(n1177), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1179), .A2(n1043), .A3(n1181), .A4(n1180), .ZN(n1177) );
NAND2_X1 U888 ( .A1(n1033), .A2(n1224), .ZN(n1180) );
NAND4_X1 U889 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1092), .ZN(n1224) );
INV_X1 U890 ( .A(G900), .ZN(n1092) );
AND3_X1 U891 ( .A1(n1034), .A2(n1206), .A3(n1051), .ZN(n1179) );
XOR2_X1 U892 ( .A(G122), .B(n1226), .Z(G24) );
NOR2_X1 U893 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U894 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
INV_X1 U895 ( .A(KEYINPUT34), .ZN(n1230) );
NOR2_X1 U896 ( .A1(n1231), .A2(n1181), .ZN(n1229) );
AND2_X1 U897 ( .A1(n1232), .A2(n1033), .ZN(n1231) );
NOR2_X1 U898 ( .A1(n1194), .A2(n1233), .ZN(n1227) );
AND2_X1 U899 ( .A1(n1234), .A2(KEYINPUT34), .ZN(n1233) );
AND2_X1 U900 ( .A1(n1234), .A2(n1235), .ZN(n1194) );
NOR4_X1 U901 ( .A1(n1208), .A2(n1030), .A3(n1210), .A4(n1074), .ZN(n1234) );
INV_X1 U902 ( .A(n1048), .ZN(n1074) );
NOR2_X1 U903 ( .A1(n1206), .A2(n1215), .ZN(n1048) );
XNOR2_X1 U904 ( .A(G119), .B(n1191), .ZN(G21) );
NAND3_X1 U905 ( .A1(n1035), .A2(n1215), .A3(n1236), .ZN(n1191) );
XNOR2_X1 U906 ( .A(n1190), .B(n1237), .ZN(G18) );
NOR2_X1 U907 ( .A1(KEYINPUT36), .A2(n1238), .ZN(n1237) );
NAND3_X1 U908 ( .A1(n1236), .A2(n1050), .A3(n1052), .ZN(n1190) );
XNOR2_X1 U909 ( .A(G113), .B(n1189), .ZN(G15) );
NAND3_X1 U910 ( .A1(n1236), .A2(n1051), .A3(n1052), .ZN(n1189) );
NOR2_X1 U911 ( .A1(n1206), .A2(n1034), .ZN(n1052) );
AND2_X1 U912 ( .A1(n1239), .A2(n1240), .ZN(n1051) );
XNOR2_X1 U913 ( .A(KEYINPUT35), .B(n1210), .ZN(n1239) );
AND2_X1 U914 ( .A1(n1043), .A2(n1235), .ZN(n1236) );
INV_X1 U915 ( .A(n1030), .ZN(n1043) );
NAND2_X1 U916 ( .A1(n1060), .A2(n1241), .ZN(n1030) );
XNOR2_X1 U917 ( .A(G110), .B(n1188), .ZN(G12) );
NAND3_X1 U918 ( .A1(n1034), .A2(n1195), .A3(n1035), .ZN(n1188) );
AND2_X1 U919 ( .A1(n1053), .A2(n1206), .ZN(n1035) );
NAND3_X1 U920 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1206) );
OR2_X1 U921 ( .A1(n1245), .A2(n1121), .ZN(n1244) );
NAND3_X1 U922 ( .A1(n1121), .A2(n1245), .A3(n1077), .ZN(n1243) );
NAND2_X1 U923 ( .A1(G217), .A2(n1246), .ZN(n1245) );
XOR2_X1 U924 ( .A(n1247), .B(n1248), .Z(n1121) );
XOR2_X1 U925 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U926 ( .A(n1251), .B(G110), .ZN(n1250) );
XOR2_X1 U927 ( .A(KEYINPUT37), .B(KEYINPUT24), .Z(n1249) );
XNOR2_X1 U928 ( .A(n1102), .B(n1252), .ZN(n1247) );
XOR2_X1 U929 ( .A(n1253), .B(n1254), .Z(n1252) );
NAND2_X1 U930 ( .A1(n1255), .A2(G221), .ZN(n1254) );
NAND2_X1 U931 ( .A1(KEYINPUT12), .A2(n1256), .ZN(n1253) );
XOR2_X1 U932 ( .A(G128), .B(G119), .Z(n1256) );
XOR2_X1 U933 ( .A(G137), .B(n1257), .Z(n1102) );
NAND2_X1 U934 ( .A1(G217), .A2(G902), .ZN(n1242) );
NAND2_X1 U935 ( .A1(n1258), .A2(n1259), .ZN(n1053) );
NAND2_X1 U936 ( .A1(n1050), .A2(n1260), .ZN(n1259) );
INV_X1 U937 ( .A(KEYINPUT35), .ZN(n1260) );
NOR2_X1 U938 ( .A1(n1210), .A2(n1240), .ZN(n1050) );
INV_X1 U939 ( .A(n1208), .ZN(n1240) );
NAND3_X1 U940 ( .A1(n1210), .A2(n1208), .A3(KEYINPUT35), .ZN(n1258) );
XOR2_X1 U941 ( .A(n1261), .B(n1083), .Z(n1208) );
INV_X1 U942 ( .A(n1134), .ZN(n1083) );
NOR2_X1 U943 ( .A1(n1140), .A2(G902), .ZN(n1134) );
INV_X1 U944 ( .A(n1137), .ZN(n1140) );
NAND3_X1 U945 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1137) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U947 ( .A1(KEYINPUT15), .A2(n1267), .ZN(n1266) );
XOR2_X1 U948 ( .A(KEYINPUT58), .B(n1268), .Z(n1267) );
XOR2_X1 U949 ( .A(n1269), .B(n1270), .Z(n1265) );
OR2_X1 U950 ( .A1(n1268), .A2(KEYINPUT15), .ZN(n1263) );
NAND3_X1 U951 ( .A1(n1271), .A2(n1268), .A3(KEYINPUT15), .ZN(n1262) );
XOR2_X1 U952 ( .A(G104), .B(n1272), .Z(n1268) );
XNOR2_X1 U953 ( .A(G122), .B(n1273), .ZN(n1272) );
XNOR2_X1 U954 ( .A(n1269), .B(n1270), .ZN(n1271) );
XOR2_X1 U955 ( .A(G146), .B(n1274), .Z(n1270) );
NOR2_X1 U956 ( .A1(KEYINPUT9), .A2(n1257), .ZN(n1274) );
XOR2_X1 U957 ( .A(G125), .B(G140), .Z(n1257) );
NAND2_X1 U958 ( .A1(n1275), .A2(KEYINPUT10), .ZN(n1269) );
XOR2_X1 U959 ( .A(n1276), .B(n1277), .Z(n1275) );
AND2_X1 U960 ( .A1(G214), .A2(n1278), .ZN(n1277) );
XOR2_X1 U961 ( .A(n1279), .B(G143), .Z(n1276) );
NAND2_X1 U962 ( .A1(KEYINPUT48), .A2(n1280), .ZN(n1279) );
INV_X1 U963 ( .A(G131), .ZN(n1280) );
NAND2_X1 U964 ( .A1(KEYINPUT59), .A2(n1138), .ZN(n1261) );
INV_X1 U965 ( .A(G475), .ZN(n1138) );
XNOR2_X1 U966 ( .A(n1281), .B(n1082), .ZN(n1210) );
NOR2_X1 U967 ( .A1(n1129), .A2(G902), .ZN(n1082) );
XNOR2_X1 U968 ( .A(n1282), .B(n1283), .ZN(n1129) );
XNOR2_X1 U969 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND2_X1 U970 ( .A1(G217), .A2(n1255), .ZN(n1284) );
NOR2_X1 U971 ( .A1(n1246), .A2(G953), .ZN(n1255) );
INV_X1 U972 ( .A(G234), .ZN(n1246) );
XNOR2_X1 U973 ( .A(n1286), .B(n1100), .ZN(n1282) );
NAND2_X1 U974 ( .A1(KEYINPUT29), .A2(n1287), .ZN(n1286) );
XOR2_X1 U975 ( .A(G107), .B(n1288), .Z(n1287) );
NOR2_X1 U976 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U977 ( .A(n1291), .B(KEYINPUT3), .Z(n1290) );
NAND2_X1 U978 ( .A1(G122), .A2(n1292), .ZN(n1291) );
NOR2_X1 U979 ( .A1(G122), .A2(n1292), .ZN(n1289) );
XNOR2_X1 U980 ( .A(KEYINPUT41), .B(n1238), .ZN(n1292) );
NAND2_X1 U981 ( .A1(KEYINPUT18), .A2(n1081), .ZN(n1281) );
INV_X1 U982 ( .A(G478), .ZN(n1081) );
AND2_X1 U983 ( .A1(n1058), .A2(n1235), .ZN(n1195) );
AND2_X1 U984 ( .A1(n1181), .A2(n1293), .ZN(n1235) );
NAND2_X1 U985 ( .A1(n1033), .A2(n1232), .ZN(n1293) );
NAND4_X1 U986 ( .A1(n1294), .A2(G953), .A3(n1110), .A4(n1225), .ZN(n1232) );
XOR2_X1 U987 ( .A(KEYINPUT1), .B(G898), .Z(n1110) );
XNOR2_X1 U988 ( .A(G902), .B(KEYINPUT45), .ZN(n1294) );
NAND3_X1 U989 ( .A1(n1225), .A2(n1037), .A3(G952), .ZN(n1033) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U991 ( .A1(n1065), .A2(n1066), .ZN(n1181) );
INV_X1 U992 ( .A(n1222), .ZN(n1066) );
NAND2_X1 U993 ( .A1(n1295), .A2(n1085), .ZN(n1222) );
NAND3_X1 U994 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1085) );
NAND2_X1 U995 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U996 ( .A1(n1078), .A2(n1077), .ZN(n1297) );
XNOR2_X1 U997 ( .A(n1201), .B(n1298), .ZN(n1078) );
XOR2_X1 U998 ( .A(n1205), .B(n1299), .Z(n1298) );
NOR3_X1 U999 ( .A1(KEYINPUT16), .A2(n1300), .A3(n1301), .ZN(n1299) );
NOR3_X1 U1000 ( .A1(KEYINPUT55), .A2(G125), .A3(n1302), .ZN(n1301) );
INV_X1 U1001 ( .A(n1303), .ZN(n1302) );
NOR2_X1 U1002 ( .A1(n1204), .A2(n1304), .ZN(n1300) );
INV_X1 U1003 ( .A(KEYINPUT55), .ZN(n1304) );
XOR2_X1 U1004 ( .A(n1303), .B(G125), .Z(n1204) );
AND2_X1 U1005 ( .A1(G224), .A2(n1037), .ZN(n1205) );
INV_X1 U1006 ( .A(G953), .ZN(n1037) );
XNOR2_X1 U1007 ( .A(n1115), .B(n1305), .ZN(n1201) );
NOR2_X1 U1008 ( .A1(KEYINPUT38), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U1009 ( .A(n1111), .B(n1116), .ZN(n1306) );
XOR2_X1 U1010 ( .A(n1307), .B(n1308), .Z(n1116) );
XNOR2_X1 U1011 ( .A(G107), .B(n1309), .ZN(n1308) );
NAND2_X1 U1012 ( .A1(KEYINPUT22), .A2(n1310), .ZN(n1307) );
XNOR2_X1 U1013 ( .A(n1311), .B(n1273), .ZN(n1111) );
INV_X1 U1014 ( .A(G113), .ZN(n1273) );
NAND2_X1 U1015 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1016 ( .A(KEYINPUT49), .B(KEYINPUT42), .Z(n1312) );
XNOR2_X1 U1017 ( .A(G110), .B(G122), .ZN(n1115) );
INV_X1 U1018 ( .A(n1076), .ZN(n1296) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1314), .ZN(n1076) );
AND2_X1 U1020 ( .A1(G214), .A2(n1314), .ZN(n1065) );
NAND2_X1 U1021 ( .A1(n1315), .A2(n1077), .ZN(n1314) );
INV_X1 U1022 ( .A(G237), .ZN(n1315) );
NOR2_X1 U1023 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
INV_X1 U1024 ( .A(n1241), .ZN(n1061) );
NAND2_X1 U1025 ( .A1(n1316), .A2(G221), .ZN(n1241) );
XOR2_X1 U1026 ( .A(n1317), .B(KEYINPUT26), .Z(n1316) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1077), .ZN(n1317) );
XNOR2_X1 U1028 ( .A(n1084), .B(n1318), .ZN(n1060) );
NOR2_X1 U1029 ( .A1(G469), .A2(KEYINPUT8), .ZN(n1318) );
NAND3_X1 U1030 ( .A1(n1319), .A2(n1320), .A3(n1077), .ZN(n1084) );
NAND2_X1 U1031 ( .A1(KEYINPUT14), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U1032 ( .A(n1322), .B(n1323), .ZN(n1321) );
NAND2_X1 U1033 ( .A1(KEYINPUT56), .A2(n1324), .ZN(n1322) );
OR3_X1 U1034 ( .A1(n1323), .A2(n1324), .A3(KEYINPUT14), .ZN(n1319) );
XOR2_X1 U1035 ( .A(n1325), .B(n1326), .Z(n1324) );
NOR2_X1 U1036 ( .A1(KEYINPUT52), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1037 ( .A(n1328), .B(G140), .Z(n1327) );
NAND2_X1 U1038 ( .A1(KEYINPUT7), .A2(G110), .ZN(n1328) );
XNOR2_X1 U1039 ( .A(n1157), .B(KEYINPUT21), .ZN(n1325) );
NOR2_X1 U1040 ( .A1(n1095), .A2(G953), .ZN(n1157) );
INV_X1 U1041 ( .A(G227), .ZN(n1095) );
XOR2_X1 U1042 ( .A(n1329), .B(n1159), .Z(n1323) );
XOR2_X1 U1043 ( .A(n1330), .B(KEYINPUT25), .Z(n1159) );
XOR2_X1 U1044 ( .A(n1162), .B(KEYINPUT32), .Z(n1329) );
XOR2_X1 U1045 ( .A(n1331), .B(n1332), .Z(n1162) );
XNOR2_X1 U1046 ( .A(n1310), .B(G101), .ZN(n1332) );
INV_X1 U1047 ( .A(G104), .ZN(n1310) );
XOR2_X1 U1048 ( .A(n1101), .B(n1333), .Z(n1331) );
NOR2_X1 U1049 ( .A1(G107), .A2(KEYINPUT57), .ZN(n1333) );
XOR2_X1 U1050 ( .A(n1334), .B(G128), .Z(n1101) );
NAND2_X1 U1051 ( .A1(n1335), .A2(KEYINPUT51), .ZN(n1334) );
XNOR2_X1 U1052 ( .A(G143), .B(n1336), .ZN(n1335) );
NOR2_X1 U1053 ( .A1(KEYINPUT53), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1054 ( .A(KEYINPUT4), .B(n1251), .ZN(n1337) );
INV_X1 U1055 ( .A(G146), .ZN(n1251) );
INV_X1 U1056 ( .A(n1215), .ZN(n1034) );
XNOR2_X1 U1057 ( .A(n1338), .B(G472), .ZN(n1215) );
NAND2_X1 U1058 ( .A1(n1339), .A2(n1077), .ZN(n1338) );
INV_X1 U1059 ( .A(G902), .ZN(n1077) );
XOR2_X1 U1060 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1061 ( .A(KEYINPUT43), .B(KEYINPUT17), .Z(n1341) );
XNOR2_X1 U1062 ( .A(n1342), .B(n1150), .ZN(n1340) );
XOR2_X1 U1063 ( .A(n1343), .B(n1344), .Z(n1150) );
XNOR2_X1 U1064 ( .A(n1345), .B(n1303), .ZN(n1344) );
XOR2_X1 U1065 ( .A(G146), .B(n1285), .Z(n1303) );
XOR2_X1 U1066 ( .A(G128), .B(G143), .Z(n1285) );
INV_X1 U1067 ( .A(n1330), .ZN(n1345) );
XNOR2_X1 U1068 ( .A(n1346), .B(n1347), .ZN(n1330) );
XNOR2_X1 U1069 ( .A(n1100), .B(n1348), .ZN(n1347) );
NOR2_X1 U1070 ( .A1(G131), .A2(KEYINPUT39), .ZN(n1348) );
INV_X1 U1071 ( .A(G134), .ZN(n1100) );
XNOR2_X1 U1072 ( .A(G137), .B(KEYINPUT28), .ZN(n1346) );
XOR2_X1 U1073 ( .A(n1349), .B(n1313), .Z(n1343) );
XNOR2_X1 U1074 ( .A(G119), .B(n1238), .ZN(n1313) );
INV_X1 U1075 ( .A(G116), .ZN(n1238) );
XNOR2_X1 U1076 ( .A(G113), .B(KEYINPUT5), .ZN(n1349) );
NAND2_X1 U1077 ( .A1(KEYINPUT46), .A2(n1144), .ZN(n1342) );
AND2_X1 U1078 ( .A1(n1350), .A2(n1351), .ZN(n1144) );
NAND2_X1 U1079 ( .A1(n1352), .A2(n1309), .ZN(n1351) );
INV_X1 U1080 ( .A(G101), .ZN(n1309) );
NAND2_X1 U1081 ( .A1(n1278), .A2(G210), .ZN(n1352) );
NAND3_X1 U1082 ( .A1(n1278), .A2(G210), .A3(G101), .ZN(n1350) );
NOR2_X1 U1083 ( .A1(G953), .A2(G237), .ZN(n1278) );
endmodule


