//Key = 0000011000111000110010010100101110000100110010001011110100011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416;

XOR2_X1 U772 ( .A(n1057), .B(n1058), .Z(G9) );
NOR2_X1 U773 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U774 ( .A(n1061), .B(KEYINPUT56), .Z(n1059) );
NAND2_X1 U775 ( .A1(KEYINPUT52), .A2(n1062), .ZN(n1057) );
INV_X1 U776 ( .A(G107), .ZN(n1062) );
NAND4_X1 U777 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(G75) );
NAND3_X1 U778 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
INV_X1 U779 ( .A(G952), .ZN(n1068) );
OR2_X1 U780 ( .A1(n1067), .A2(n1069), .ZN(n1065) );
INV_X1 U781 ( .A(KEYINPUT53), .ZN(n1069) );
NAND2_X1 U782 ( .A1(G952), .A2(n1070), .ZN(n1063) );
NAND3_X1 U783 ( .A1(n1071), .A2(n1067), .A3(n1072), .ZN(n1070) );
INV_X1 U784 ( .A(n1073), .ZN(n1072) );
NAND4_X1 U785 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1067) );
NOR3_X1 U786 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
XOR2_X1 U787 ( .A(n1081), .B(n1082), .Z(n1079) );
XOR2_X1 U788 ( .A(KEYINPUT17), .B(G469), .Z(n1082) );
NAND3_X1 U789 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1078) );
NAND2_X1 U790 ( .A1(G472), .A2(n1086), .ZN(n1085) );
NOR3_X1 U791 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1076) );
NOR2_X1 U792 ( .A1(KEYINPUT21), .A2(n1090), .ZN(n1089) );
NOR2_X1 U793 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND2_X1 U794 ( .A1(n1086), .A2(KEYINPUT34), .ZN(n1092) );
NOR3_X1 U795 ( .A1(KEYINPUT34), .A2(G472), .A3(n1086), .ZN(n1091) );
NOR2_X1 U796 ( .A1(n1093), .A2(n1094), .ZN(n1088) );
INV_X1 U797 ( .A(KEYINPUT21), .ZN(n1094) );
NOR2_X1 U798 ( .A1(G472), .A2(n1095), .ZN(n1093) );
XOR2_X1 U799 ( .A(n1086), .B(KEYINPUT34), .Z(n1095) );
XNOR2_X1 U800 ( .A(n1096), .B(n1097), .ZN(n1087) );
NOR2_X1 U801 ( .A1(KEYINPUT58), .A2(n1098), .ZN(n1097) );
NAND2_X1 U802 ( .A1(n1099), .A2(n1100), .ZN(n1071) );
NAND2_X1 U803 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND3_X1 U804 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NAND3_X1 U805 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1104) );
NAND2_X1 U806 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U807 ( .A1(n1111), .A2(n1112), .ZN(n1106) );
NAND2_X1 U808 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U809 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND3_X1 U810 ( .A1(n1111), .A2(n1117), .A3(n1109), .ZN(n1101) );
NAND2_X1 U811 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U812 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
OR2_X1 U813 ( .A1(n1083), .A2(n1105), .ZN(n1121) );
NAND2_X1 U814 ( .A1(n1123), .A2(n1083), .ZN(n1120) );
NAND2_X1 U815 ( .A1(n1105), .A2(n1124), .ZN(n1118) );
INV_X1 U816 ( .A(n1125), .ZN(n1099) );
XOR2_X1 U817 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U818 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U819 ( .A1(n1130), .A2(G953), .ZN(n1129) );
NAND3_X1 U820 ( .A1(n1131), .A2(n1132), .A3(KEYINPUT59), .ZN(n1128) );
NAND2_X1 U821 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XNOR2_X1 U822 ( .A(n1135), .B(n1136), .ZN(n1131) );
NAND2_X1 U823 ( .A1(KEYINPUT30), .A2(n1137), .ZN(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U825 ( .A(n1140), .B(G131), .Z(n1139) );
NAND2_X1 U826 ( .A1(KEYINPUT32), .A2(n1141), .ZN(n1140) );
NAND2_X1 U827 ( .A1(G953), .A2(n1142), .ZN(n1126) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1142) );
XOR2_X1 U829 ( .A(n1143), .B(n1144), .Z(G69) );
XOR2_X1 U830 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U831 ( .A1(n1147), .A2(n1064), .ZN(n1146) );
AND2_X1 U832 ( .A1(G224), .A2(G898), .ZN(n1147) );
NAND2_X1 U833 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
NAND2_X1 U834 ( .A1(n1064), .A2(n1150), .ZN(n1143) );
NAND2_X1 U835 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U836 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XOR2_X1 U837 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND4_X1 U838 ( .A1(n1157), .A2(G217), .A3(n1158), .A4(n1073), .ZN(n1155) );
XOR2_X1 U839 ( .A(n1159), .B(KEYINPUT8), .Z(n1157) );
NOR2_X1 U840 ( .A1(n1153), .A2(n1160), .ZN(G63) );
XNOR2_X1 U841 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U843 ( .A(G478), .ZN(n1163) );
NOR2_X1 U844 ( .A1(n1153), .A2(n1165), .ZN(G60) );
XOR2_X1 U845 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U846 ( .A1(n1168), .A2(n1164), .ZN(n1167) );
XOR2_X1 U847 ( .A(n1169), .B(n1170), .Z(G6) );
NOR2_X1 U848 ( .A1(n1153), .A2(n1171), .ZN(G57) );
XOR2_X1 U849 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND3_X1 U851 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
NAND2_X1 U852 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
INV_X1 U853 ( .A(KEYINPUT20), .ZN(n1180) );
NAND2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
XOR2_X1 U855 ( .A(KEYINPUT61), .B(n1183), .Z(n1181) );
NAND2_X1 U856 ( .A1(KEYINPUT20), .A2(n1184), .ZN(n1176) );
NAND2_X1 U857 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
OR3_X1 U858 ( .A1(n1187), .A2(n1188), .A3(KEYINPUT61), .ZN(n1186) );
NAND2_X1 U859 ( .A1(KEYINPUT61), .A2(n1188), .ZN(n1185) );
XOR2_X1 U860 ( .A(n1189), .B(n1190), .Z(n1172) );
XNOR2_X1 U861 ( .A(n1191), .B(n1192), .ZN(n1190) );
NOR2_X1 U862 ( .A1(KEYINPUT49), .A2(n1193), .ZN(n1191) );
XOR2_X1 U863 ( .A(KEYINPUT42), .B(n1194), .Z(n1193) );
NOR2_X1 U864 ( .A1(n1195), .A2(n1164), .ZN(n1189) );
INV_X1 U865 ( .A(G472), .ZN(n1195) );
NOR2_X1 U866 ( .A1(n1153), .A2(n1196), .ZN(G54) );
XOR2_X1 U867 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U868 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U869 ( .A1(n1201), .A2(n1164), .ZN(n1200) );
NAND2_X1 U870 ( .A1(KEYINPUT23), .A2(n1202), .ZN(n1199) );
XOR2_X1 U871 ( .A(n1203), .B(n1204), .Z(n1197) );
XOR2_X1 U872 ( .A(G140), .B(G110), .Z(n1204) );
NAND3_X1 U873 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1203) );
NAND2_X1 U874 ( .A1(n1208), .A2(n1183), .ZN(n1207) );
NAND2_X1 U875 ( .A1(KEYINPUT22), .A2(n1209), .ZN(n1206) );
NAND2_X1 U876 ( .A1(n1210), .A2(n1188), .ZN(n1209) );
XNOR2_X1 U877 ( .A(KEYINPUT45), .B(n1208), .ZN(n1210) );
NAND2_X1 U878 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
INV_X1 U879 ( .A(KEYINPUT22), .ZN(n1212) );
NAND2_X1 U880 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
OR3_X1 U881 ( .A1(n1208), .A2(n1183), .A3(KEYINPUT45), .ZN(n1214) );
NAND2_X1 U882 ( .A1(KEYINPUT45), .A2(n1208), .ZN(n1213) );
XNOR2_X1 U883 ( .A(n1215), .B(n1138), .ZN(n1208) );
NOR2_X1 U884 ( .A1(n1153), .A2(n1216), .ZN(G51) );
XOR2_X1 U885 ( .A(n1148), .B(n1217), .Z(n1216) );
XOR2_X1 U886 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR3_X1 U887 ( .A1(n1220), .A2(n1096), .A3(n1164), .ZN(n1219) );
NAND2_X1 U888 ( .A1(n1159), .A2(n1073), .ZN(n1164) );
NAND3_X1 U889 ( .A1(n1130), .A2(n1151), .A3(n1221), .ZN(n1073) );
XOR2_X1 U890 ( .A(n1152), .B(KEYINPUT35), .Z(n1221) );
AND4_X1 U891 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1151) );
NOR3_X1 U892 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1225) );
NOR2_X1 U893 ( .A1(n1061), .A2(n1060), .ZN(n1228) );
NAND3_X1 U894 ( .A1(n1229), .A2(n1230), .A3(n1111), .ZN(n1060) );
INV_X1 U895 ( .A(n1170), .ZN(n1227) );
NAND4_X1 U896 ( .A1(n1231), .A2(n1124), .A3(n1111), .A4(n1229), .ZN(n1170) );
NOR2_X1 U897 ( .A1(n1123), .A2(n1232), .ZN(n1226) );
NOR2_X1 U898 ( .A1(n1231), .A2(n1230), .ZN(n1123) );
AND4_X1 U899 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1130) );
AND4_X1 U900 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NAND2_X1 U901 ( .A1(n1241), .A2(n1242), .ZN(n1235) );
NAND2_X1 U902 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U903 ( .A(KEYINPUT6), .B(n1230), .Z(n1244) );
XOR2_X1 U904 ( .A(n1245), .B(KEYINPUT4), .Z(n1243) );
NAND3_X1 U905 ( .A1(n1246), .A2(n1124), .A3(n1109), .ZN(n1234) );
XOR2_X1 U906 ( .A(n1247), .B(KEYINPUT41), .Z(n1159) );
XOR2_X1 U907 ( .A(KEYINPUT63), .B(KEYINPUT27), .Z(n1220) );
NAND2_X1 U908 ( .A1(n1248), .A2(n1249), .ZN(n1218) );
NAND2_X1 U909 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
INV_X1 U910 ( .A(n1252), .ZN(n1248) );
NOR2_X1 U911 ( .A1(n1064), .A2(G952), .ZN(n1153) );
XOR2_X1 U912 ( .A(n1253), .B(n1240), .Z(G48) );
NAND3_X1 U913 ( .A1(n1231), .A2(n1080), .A3(n1254), .ZN(n1240) );
XNOR2_X1 U914 ( .A(G143), .B(n1239), .ZN(G45) );
NAND4_X1 U915 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1239) );
XNOR2_X1 U916 ( .A(G140), .B(n1258), .ZN(G42) );
NAND4_X1 U917 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1258) );
NOR2_X1 U918 ( .A1(n1061), .A2(n1245), .ZN(n1262) );
XOR2_X1 U919 ( .A(KEYINPUT29), .B(n1110), .Z(n1261) );
XOR2_X1 U920 ( .A(KEYINPUT54), .B(n1109), .Z(n1259) );
XNOR2_X1 U921 ( .A(G137), .B(n1238), .ZN(G39) );
NAND4_X1 U922 ( .A1(n1109), .A2(n1263), .A3(n1260), .A4(n1080), .ZN(n1238) );
XOR2_X1 U923 ( .A(n1264), .B(n1265), .Z(G36) );
NOR2_X1 U924 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U925 ( .A(n1268), .B(KEYINPUT51), .Z(n1264) );
XOR2_X1 U926 ( .A(G131), .B(n1269), .Z(G33) );
NOR2_X1 U927 ( .A1(n1245), .A2(n1267), .ZN(n1269) );
INV_X1 U928 ( .A(n1241), .ZN(n1267) );
NOR3_X1 U929 ( .A1(n1061), .A2(n1270), .A3(n1107), .ZN(n1241) );
NAND3_X1 U930 ( .A1(n1255), .A2(n1271), .A3(n1109), .ZN(n1107) );
NOR2_X1 U931 ( .A1(n1272), .A2(n1115), .ZN(n1109) );
INV_X1 U932 ( .A(n1084), .ZN(n1115) );
XOR2_X1 U933 ( .A(n1273), .B(n1274), .Z(G30) );
XOR2_X1 U934 ( .A(KEYINPUT26), .B(G128), .Z(n1274) );
NAND2_X1 U935 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
OR2_X1 U936 ( .A1(n1233), .A2(KEYINPUT36), .ZN(n1276) );
NAND3_X1 U937 ( .A1(n1230), .A2(n1080), .A3(n1254), .ZN(n1233) );
NOR4_X1 U938 ( .A1(n1061), .A2(n1113), .A3(n1277), .A4(n1270), .ZN(n1254) );
NAND4_X1 U939 ( .A1(n1278), .A2(n1230), .A3(n1279), .A4(KEYINPUT36), .ZN(n1275) );
NOR3_X1 U940 ( .A1(n1270), .A2(n1255), .A3(n1124), .ZN(n1279) );
INV_X1 U941 ( .A(n1260), .ZN(n1270) );
INV_X1 U942 ( .A(n1266), .ZN(n1230) );
NOR2_X1 U943 ( .A1(n1277), .A2(n1113), .ZN(n1278) );
XNOR2_X1 U944 ( .A(G101), .B(n1280), .ZN(G3) );
NAND2_X1 U945 ( .A1(KEYINPUT28), .A2(n1281), .ZN(n1280) );
INV_X1 U946 ( .A(n1152), .ZN(n1281) );
NAND3_X1 U947 ( .A1(n1229), .A2(n1255), .A3(n1263), .ZN(n1152) );
NOR3_X1 U948 ( .A1(n1061), .A2(n1277), .A3(n1282), .ZN(n1263) );
INV_X1 U949 ( .A(n1124), .ZN(n1061) );
NAND2_X1 U950 ( .A1(n1283), .A2(n1284), .ZN(G27) );
NAND2_X1 U951 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U952 ( .A1(G125), .A2(n1287), .ZN(n1283) );
NAND2_X1 U953 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U954 ( .A1(KEYINPUT46), .A2(n1290), .ZN(n1289) );
INV_X1 U955 ( .A(n1237), .ZN(n1290) );
OR2_X1 U956 ( .A1(n1285), .A2(KEYINPUT46), .ZN(n1288) );
NOR2_X1 U957 ( .A1(KEYINPUT2), .A2(n1237), .ZN(n1285) );
NAND3_X1 U958 ( .A1(n1103), .A2(n1291), .A3(n1246), .ZN(n1237) );
AND3_X1 U959 ( .A1(n1231), .A2(n1260), .A3(n1110), .ZN(n1246) );
NAND2_X1 U960 ( .A1(n1125), .A2(n1292), .ZN(n1260) );
NAND4_X1 U961 ( .A1(G902), .A2(n1133), .A3(n1293), .A4(n1134), .ZN(n1292) );
INV_X1 U962 ( .A(G900), .ZN(n1134) );
XOR2_X1 U963 ( .A(n1294), .B(n1224), .Z(G24) );
NAND3_X1 U964 ( .A1(n1103), .A2(n1111), .A3(n1295), .ZN(n1224) );
NOR3_X1 U965 ( .A1(n1296), .A2(n1074), .A3(n1075), .ZN(n1295) );
NOR2_X1 U966 ( .A1(n1080), .A2(n1271), .ZN(n1111) );
XNOR2_X1 U967 ( .A(G119), .B(n1222), .ZN(G21) );
NAND3_X1 U968 ( .A1(n1105), .A2(n1080), .A3(n1297), .ZN(n1222) );
XOR2_X1 U969 ( .A(G116), .B(n1298), .Z(G18) );
NOR2_X1 U970 ( .A1(n1266), .A2(n1232), .ZN(n1298) );
NAND2_X1 U971 ( .A1(n1074), .A2(n1256), .ZN(n1266) );
INV_X1 U972 ( .A(n1075), .ZN(n1256) );
XOR2_X1 U973 ( .A(G113), .B(n1299), .Z(G15) );
NOR2_X1 U974 ( .A1(n1232), .A2(n1300), .ZN(n1299) );
XOR2_X1 U975 ( .A(KEYINPUT48), .B(n1231), .Z(n1300) );
INV_X1 U976 ( .A(n1245), .ZN(n1231) );
NAND2_X1 U977 ( .A1(n1301), .A2(n1257), .ZN(n1245) );
INV_X1 U978 ( .A(n1074), .ZN(n1257) );
NAND2_X1 U979 ( .A1(n1297), .A2(n1255), .ZN(n1232) );
AND3_X1 U980 ( .A1(n1229), .A2(n1271), .A3(n1103), .ZN(n1297) );
AND2_X1 U981 ( .A1(n1122), .A2(n1083), .ZN(n1103) );
XOR2_X1 U982 ( .A(n1302), .B(n1223), .Z(G12) );
NAND4_X1 U983 ( .A1(n1105), .A2(n1110), .A3(n1124), .A4(n1229), .ZN(n1223) );
INV_X1 U984 ( .A(n1296), .ZN(n1229) );
NAND2_X1 U985 ( .A1(n1291), .A2(n1303), .ZN(n1296) );
NAND2_X1 U986 ( .A1(n1304), .A2(n1125), .ZN(n1303) );
NAND3_X1 U987 ( .A1(n1293), .A2(n1064), .A3(G952), .ZN(n1125) );
NAND3_X1 U988 ( .A1(G902), .A2(n1293), .A3(n1305), .ZN(n1304) );
INV_X1 U989 ( .A(n1149), .ZN(n1305) );
NAND2_X1 U990 ( .A1(n1133), .A2(n1306), .ZN(n1149) );
INV_X1 U991 ( .A(G898), .ZN(n1306) );
XOR2_X1 U992 ( .A(G953), .B(KEYINPUT3), .Z(n1133) );
NAND2_X1 U993 ( .A1(G237), .A2(G234), .ZN(n1293) );
INV_X1 U994 ( .A(n1113), .ZN(n1291) );
NAND2_X1 U995 ( .A1(n1272), .A2(n1084), .ZN(n1113) );
NAND2_X1 U996 ( .A1(n1307), .A2(G214), .ZN(n1084) );
XOR2_X1 U997 ( .A(n1308), .B(KEYINPUT14), .Z(n1307) );
INV_X1 U998 ( .A(n1116), .ZN(n1272) );
XNOR2_X1 U999 ( .A(n1098), .B(n1096), .ZN(n1116) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1308), .ZN(n1096) );
OR2_X1 U1001 ( .A1(G902), .A2(G237), .ZN(n1308) );
NAND2_X1 U1002 ( .A1(n1309), .A2(n1247), .ZN(n1098) );
XOR2_X1 U1003 ( .A(n1310), .B(n1311), .Z(n1309) );
NAND2_X1 U1004 ( .A1(KEYINPUT62), .A2(n1148), .ZN(n1311) );
XOR2_X1 U1005 ( .A(n1312), .B(n1313), .Z(n1148) );
XOR2_X1 U1006 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1007 ( .A(n1316), .B(KEYINPUT55), .Z(n1315) );
NAND2_X1 U1008 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1009 ( .A1(n1319), .A2(n1302), .ZN(n1318) );
NAND2_X1 U1010 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U1011 ( .A1(KEYINPUT25), .A2(n1294), .ZN(n1321) );
INV_X1 U1012 ( .A(G122), .ZN(n1294) );
NAND2_X1 U1013 ( .A1(G122), .A2(n1322), .ZN(n1317) );
NAND2_X1 U1014 ( .A1(KEYINPUT25), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1015 ( .A1(G110), .A2(n1320), .ZN(n1323) );
INV_X1 U1016 ( .A(KEYINPUT18), .ZN(n1320) );
NAND2_X1 U1017 ( .A1(n1324), .A2(n1325), .ZN(n1314) );
INV_X1 U1018 ( .A(G113), .ZN(n1325) );
XOR2_X1 U1019 ( .A(KEYINPUT39), .B(KEYINPUT31), .Z(n1324) );
XOR2_X1 U1020 ( .A(n1326), .B(n1327), .Z(n1312) );
XOR2_X1 U1021 ( .A(n1328), .B(n1329), .Z(n1327) );
NAND2_X1 U1022 ( .A1(n1330), .A2(n1331), .ZN(n1326) );
NAND2_X1 U1023 ( .A1(KEYINPUT5), .A2(n1332), .ZN(n1331) );
OR3_X1 U1024 ( .A1(n1169), .A2(G107), .A3(KEYINPUT5), .ZN(n1330) );
NAND2_X1 U1025 ( .A1(n1333), .A2(n1334), .ZN(n1310) );
NAND2_X1 U1026 ( .A1(n1250), .A2(n1335), .ZN(n1334) );
NAND2_X1 U1027 ( .A1(KEYINPUT11), .A2(G224), .ZN(n1335) );
NAND2_X1 U1028 ( .A1(n1252), .A2(KEYINPUT11), .ZN(n1333) );
NOR2_X1 U1029 ( .A1(n1251), .A2(n1250), .ZN(n1252) );
XOR2_X1 U1030 ( .A(G125), .B(n1187), .Z(n1250) );
NAND2_X1 U1031 ( .A1(G224), .A2(n1064), .ZN(n1251) );
NOR2_X1 U1032 ( .A1(n1336), .A2(n1122), .ZN(n1124) );
XOR2_X1 U1033 ( .A(n1201), .B(n1337), .Z(n1122) );
NOR2_X1 U1034 ( .A1(KEYINPUT33), .A2(n1081), .ZN(n1337) );
NAND2_X1 U1035 ( .A1(n1338), .A2(n1247), .ZN(n1081) );
XOR2_X1 U1036 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1037 ( .A(G140), .B(n1341), .Z(n1340) );
NOR2_X1 U1038 ( .A1(KEYINPUT15), .A2(n1302), .ZN(n1341) );
NAND2_X1 U1039 ( .A1(n1342), .A2(n1343), .ZN(n1339) );
NAND2_X1 U1040 ( .A1(n1344), .A2(n1183), .ZN(n1343) );
XOR2_X1 U1041 ( .A(KEYINPUT13), .B(n1345), .Z(n1344) );
NAND2_X1 U1042 ( .A1(n1346), .A2(n1188), .ZN(n1342) );
XNOR2_X1 U1043 ( .A(n1345), .B(KEYINPUT19), .ZN(n1346) );
XOR2_X1 U1044 ( .A(n1347), .B(n1202), .Z(n1345) );
NAND2_X1 U1045 ( .A1(G227), .A2(n1064), .ZN(n1202) );
INV_X1 U1046 ( .A(G953), .ZN(n1064) );
NAND2_X1 U1047 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1048 ( .A1(n1138), .A2(n1215), .ZN(n1349) );
XOR2_X1 U1049 ( .A(n1350), .B(KEYINPUT47), .Z(n1348) );
OR2_X1 U1050 ( .A1(n1215), .A2(n1138), .ZN(n1350) );
XNOR2_X1 U1051 ( .A(n1351), .B(n1352), .ZN(n1138) );
XNOR2_X1 U1052 ( .A(n1332), .B(n1175), .ZN(n1215) );
XOR2_X1 U1053 ( .A(n1169), .B(G107), .Z(n1332) );
INV_X1 U1054 ( .A(G469), .ZN(n1201) );
XOR2_X1 U1055 ( .A(KEYINPUT12), .B(n1083), .Z(n1336) );
NAND2_X1 U1056 ( .A1(G221), .A2(n1158), .ZN(n1083) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1247), .ZN(n1158) );
NOR2_X1 U1058 ( .A1(n1271), .A2(n1255), .ZN(n1110) );
INV_X1 U1059 ( .A(n1080), .ZN(n1255) );
NAND3_X1 U1060 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1080) );
OR2_X1 U1061 ( .A1(n1356), .A2(n1156), .ZN(n1355) );
NAND3_X1 U1062 ( .A1(n1156), .A2(n1356), .A3(n1247), .ZN(n1354) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1064 ( .A(n1358), .B(n1359), .ZN(n1156) );
XOR2_X1 U1065 ( .A(G110), .B(n1360), .Z(n1359) );
XOR2_X1 U1066 ( .A(G137), .B(G119), .Z(n1360) );
XOR2_X1 U1067 ( .A(n1361), .B(n1136), .Z(n1358) );
XOR2_X1 U1068 ( .A(n1362), .B(n1351), .Z(n1361) );
XOR2_X1 U1069 ( .A(n1363), .B(n1253), .Z(n1351) );
NAND2_X1 U1070 ( .A1(G221), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1071 ( .A1(G902), .A2(G217), .ZN(n1353) );
INV_X1 U1072 ( .A(n1277), .ZN(n1271) );
XOR2_X1 U1073 ( .A(n1086), .B(G472), .Z(n1277) );
NAND2_X1 U1074 ( .A1(n1365), .A2(n1247), .ZN(n1086) );
XOR2_X1 U1075 ( .A(n1366), .B(n1367), .Z(n1365) );
XOR2_X1 U1076 ( .A(n1192), .B(n1368), .Z(n1367) );
NAND2_X1 U1077 ( .A1(n1369), .A2(KEYINPUT16), .ZN(n1368) );
XOR2_X1 U1078 ( .A(n1370), .B(n1194), .Z(n1369) );
XOR2_X1 U1079 ( .A(G113), .B(n1329), .Z(n1194) );
XOR2_X1 U1080 ( .A(G116), .B(G119), .Z(n1329) );
NAND2_X1 U1081 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NAND2_X1 U1082 ( .A1(n1183), .A2(n1182), .ZN(n1372) );
INV_X1 U1083 ( .A(n1187), .ZN(n1182) );
XOR2_X1 U1084 ( .A(n1178), .B(KEYINPUT43), .Z(n1371) );
NAND2_X1 U1085 ( .A1(n1187), .A2(n1188), .ZN(n1178) );
INV_X1 U1086 ( .A(n1183), .ZN(n1188) );
XOR2_X1 U1087 ( .A(G131), .B(n1141), .Z(n1183) );
XOR2_X1 U1088 ( .A(G137), .B(n1268), .Z(n1141) );
XOR2_X1 U1089 ( .A(n1373), .B(G128), .Z(n1187) );
NAND3_X1 U1090 ( .A1(n1374), .A2(n1375), .A3(n1376), .ZN(n1373) );
NAND2_X1 U1091 ( .A1(n1352), .A2(n1253), .ZN(n1376) );
NAND2_X1 U1092 ( .A1(n1377), .A2(n1378), .ZN(n1375) );
INV_X1 U1093 ( .A(KEYINPUT10), .ZN(n1378) );
NAND2_X1 U1094 ( .A1(n1379), .A2(n1380), .ZN(n1377) );
XOR2_X1 U1095 ( .A(KEYINPUT37), .B(n1253), .Z(n1379) );
INV_X1 U1096 ( .A(G146), .ZN(n1253) );
NAND2_X1 U1097 ( .A1(KEYINPUT10), .A2(n1381), .ZN(n1374) );
NAND2_X1 U1098 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
OR2_X1 U1099 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1383) );
NAND3_X1 U1100 ( .A1(G146), .A2(n1380), .A3(KEYINPUT37), .ZN(n1382) );
NAND2_X1 U1101 ( .A1(G210), .A2(n1384), .ZN(n1192) );
NAND2_X1 U1102 ( .A1(KEYINPUT40), .A2(n1328), .ZN(n1366) );
INV_X1 U1103 ( .A(n1175), .ZN(n1328) );
XNOR2_X1 U1104 ( .A(G101), .B(KEYINPUT38), .ZN(n1175) );
INV_X1 U1105 ( .A(n1282), .ZN(n1105) );
NAND2_X1 U1106 ( .A1(n1301), .A2(n1074), .ZN(n1282) );
XOR2_X1 U1107 ( .A(n1168), .B(n1385), .Z(n1074) );
NOR2_X1 U1108 ( .A1(G902), .A2(n1166), .ZN(n1385) );
NAND2_X1 U1109 ( .A1(n1386), .A2(n1387), .ZN(n1166) );
NAND2_X1 U1110 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1111 ( .A1(n1390), .A2(n1391), .ZN(n1388) );
NAND2_X1 U1112 ( .A1(KEYINPUT50), .A2(n1392), .ZN(n1391) );
INV_X1 U1113 ( .A(KEYINPUT9), .ZN(n1390) );
NAND2_X1 U1114 ( .A1(n1393), .A2(n1394), .ZN(n1386) );
NAND2_X1 U1115 ( .A1(KEYINPUT50), .A2(n1395), .ZN(n1394) );
OR2_X1 U1116 ( .A1(n1389), .A2(KEYINPUT9), .ZN(n1395) );
NAND2_X1 U1117 ( .A1(n1396), .A2(n1397), .ZN(n1389) );
NAND2_X1 U1118 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
XOR2_X1 U1119 ( .A(KEYINPUT60), .B(n1400), .Z(n1396) );
NOR2_X1 U1120 ( .A1(n1398), .A2(n1399), .ZN(n1400) );
XOR2_X1 U1121 ( .A(G146), .B(n1136), .Z(n1399) );
XNOR2_X1 U1122 ( .A(n1286), .B(G140), .ZN(n1136) );
INV_X1 U1123 ( .A(G125), .ZN(n1286) );
XOR2_X1 U1124 ( .A(n1401), .B(n1402), .Z(n1398) );
XOR2_X1 U1125 ( .A(G131), .B(n1403), .Z(n1402) );
NOR2_X1 U1126 ( .A1(KEYINPUT1), .A2(n1404), .ZN(n1403) );
XOR2_X1 U1127 ( .A(KEYINPUT0), .B(n1352), .Z(n1404) );
NAND2_X1 U1128 ( .A1(G214), .A2(n1384), .ZN(n1401) );
NOR2_X1 U1129 ( .A1(G953), .A2(G237), .ZN(n1384) );
INV_X1 U1130 ( .A(n1392), .ZN(n1393) );
XOR2_X1 U1131 ( .A(n1169), .B(n1405), .Z(n1392) );
XOR2_X1 U1132 ( .A(G122), .B(G113), .Z(n1405) );
INV_X1 U1133 ( .A(G104), .ZN(n1169) );
INV_X1 U1134 ( .A(G475), .ZN(n1168) );
XOR2_X1 U1135 ( .A(n1075), .B(KEYINPUT24), .Z(n1301) );
XOR2_X1 U1136 ( .A(n1406), .B(G478), .Z(n1075) );
NAND2_X1 U1137 ( .A1(n1161), .A2(n1247), .ZN(n1406) );
INV_X1 U1138 ( .A(G902), .ZN(n1247) );
XNOR2_X1 U1139 ( .A(n1407), .B(n1408), .ZN(n1161) );
XOR2_X1 U1140 ( .A(G107), .B(n1409), .Z(n1408) );
XOR2_X1 U1141 ( .A(G122), .B(G116), .Z(n1409) );
XOR2_X1 U1142 ( .A(n1410), .B(n1411), .Z(n1407) );
AND3_X1 U1143 ( .A1(n1364), .A2(n1412), .A3(G217), .ZN(n1411) );
INV_X1 U1144 ( .A(KEYINPUT57), .ZN(n1412) );
NOR2_X1 U1145 ( .A1(n1357), .A2(G953), .ZN(n1364) );
INV_X1 U1146 ( .A(G234), .ZN(n1357) );
NAND2_X1 U1147 ( .A1(n1413), .A2(n1414), .ZN(n1410) );
NAND2_X1 U1148 ( .A1(n1415), .A2(n1268), .ZN(n1414) );
XOR2_X1 U1149 ( .A(KEYINPUT44), .B(n1416), .Z(n1413) );
NOR2_X1 U1150 ( .A1(n1415), .A2(n1268), .ZN(n1416) );
INV_X1 U1151 ( .A(G134), .ZN(n1268) );
XOR2_X1 U1152 ( .A(n1363), .B(n1352), .Z(n1415) );
INV_X1 U1153 ( .A(n1380), .ZN(n1352) );
XNOR2_X1 U1154 ( .A(G143), .B(KEYINPUT7), .ZN(n1380) );
INV_X1 U1155 ( .A(G128), .ZN(n1363) );
INV_X1 U1156 ( .A(G110), .ZN(n1302) );
endmodule


