//Key = 0011110011001011001101000101011101100000100010111100000010100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298;

XOR2_X1 U705 ( .A(G107), .B(n987), .Z(G9) );
NOR2_X1 U706 ( .A1(n988), .A2(n989), .ZN(G75) );
NOR4_X1 U707 ( .A1(n990), .A2(n991), .A3(G953), .A4(n992), .ZN(n989) );
NOR2_X1 U708 ( .A1(n993), .A2(n994), .ZN(n991) );
XOR2_X1 U709 ( .A(n995), .B(KEYINPUT52), .Z(n993) );
NAND4_X1 U710 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(n995) );
XOR2_X1 U711 ( .A(KEYINPUT37), .B(n1000), .Z(n999) );
NAND2_X1 U712 ( .A1(n1001), .A2(n1002), .ZN(n990) );
NAND2_X1 U713 ( .A1(n996), .A2(n1003), .ZN(n1002) );
NAND2_X1 U714 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U715 ( .A1(n1000), .A2(n1006), .ZN(n1005) );
NAND2_X1 U716 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U717 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND3_X1 U718 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NAND2_X1 U719 ( .A1(n1014), .A2(n997), .ZN(n1013) );
NAND2_X1 U720 ( .A1(n998), .A2(n1015), .ZN(n1011) );
NAND2_X1 U721 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
XOR2_X1 U722 ( .A(KEYINPUT27), .B(n1018), .Z(n1016) );
NAND4_X1 U723 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n998), .ZN(n1007) );
INV_X1 U724 ( .A(n1022), .ZN(n1020) );
XNOR2_X1 U725 ( .A(n997), .B(KEYINPUT56), .ZN(n1019) );
NAND4_X1 U726 ( .A1(n1009), .A2(n997), .A3(n998), .A4(n1023), .ZN(n1004) );
NAND2_X1 U727 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U728 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
INV_X1 U729 ( .A(n1028), .ZN(n996) );
NOR3_X1 U730 ( .A1(n992), .A2(G953), .A3(G952), .ZN(n988) );
AND4_X1 U731 ( .A1(n1029), .A2(n1022), .A3(n1030), .A4(n1031), .ZN(n992) );
NOR4_X1 U732 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
XOR2_X1 U733 ( .A(KEYINPUT54), .B(n1036), .Z(n1035) );
XOR2_X1 U734 ( .A(n1037), .B(n1038), .Z(n1032) );
XNOR2_X1 U735 ( .A(KEYINPUT35), .B(KEYINPUT30), .ZN(n1037) );
NOR3_X1 U736 ( .A1(n1027), .A2(n1039), .A3(n1040), .ZN(n1030) );
INV_X1 U737 ( .A(n1041), .ZN(n1040) );
XOR2_X1 U738 ( .A(n1042), .B(n1043), .Z(n1029) );
XNOR2_X1 U739 ( .A(G472), .B(KEYINPUT40), .ZN(n1043) );
XOR2_X1 U740 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U741 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
AND2_X1 U742 ( .A1(G227), .A2(G900), .ZN(n1046) );
NAND2_X1 U743 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NAND2_X1 U744 ( .A1(n1050), .A2(n1047), .ZN(n1049) );
XOR2_X1 U745 ( .A(n1051), .B(n1052), .Z(n1050) );
NAND3_X1 U746 ( .A1(n1053), .A2(n1052), .A3(G953), .ZN(n1048) );
XOR2_X1 U747 ( .A(n1054), .B(n1055), .Z(n1052) );
XOR2_X1 U748 ( .A(n1056), .B(n1057), .Z(n1055) );
XOR2_X1 U749 ( .A(n1058), .B(n1059), .Z(n1054) );
NOR2_X1 U750 ( .A1(G140), .A2(KEYINPUT57), .ZN(n1059) );
XOR2_X1 U751 ( .A(n1060), .B(n1061), .Z(n1058) );
NOR2_X1 U752 ( .A1(G131), .A2(KEYINPUT7), .ZN(n1061) );
XOR2_X1 U753 ( .A(n1062), .B(KEYINPUT61), .Z(n1053) );
XOR2_X1 U754 ( .A(n1063), .B(n1064), .Z(G69) );
AND2_X1 U755 ( .A1(n1065), .A2(n1047), .ZN(n1064) );
NAND2_X1 U756 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NAND2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U758 ( .A(n1070), .ZN(n1068) );
NAND2_X1 U759 ( .A1(n1071), .A2(n1070), .ZN(n1066) );
NAND2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XNOR2_X1 U761 ( .A(n1074), .B(n1075), .ZN(n1072) );
NAND2_X1 U762 ( .A1(n1073), .A2(n1069), .ZN(n1071) );
NAND2_X1 U763 ( .A1(G953), .A2(n1076), .ZN(n1069) );
INV_X1 U764 ( .A(G224), .ZN(n1076) );
INV_X1 U765 ( .A(n1077), .ZN(n1073) );
NOR2_X1 U766 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XNOR2_X1 U767 ( .A(n1080), .B(n1081), .ZN(n1079) );
NAND2_X1 U768 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
XOR2_X1 U769 ( .A(KEYINPUT39), .B(G217), .Z(n1083) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1084), .ZN(G63) );
NOR2_X1 U771 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U772 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U774 ( .A1(n1082), .A2(G478), .ZN(n1087) );
NOR2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1085) );
INV_X1 U776 ( .A(KEYINPUT41), .ZN(n1090) );
NOR2_X1 U777 ( .A1(n1078), .A2(n1091), .ZN(G60) );
XOR2_X1 U778 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND3_X1 U779 ( .A1(n1094), .A2(n1095), .A3(G475), .ZN(n1092) );
OR2_X1 U780 ( .A1(n1082), .A2(KEYINPUT51), .ZN(n1095) );
NAND2_X1 U781 ( .A1(KEYINPUT51), .A2(n1096), .ZN(n1094) );
NAND2_X1 U782 ( .A1(n1001), .A2(G902), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(G6) );
NAND2_X1 U784 ( .A1(G104), .A2(n1099), .ZN(n1098) );
NAND2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U787 ( .A(KEYINPUT58), .ZN(n1103) );
NAND2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
INV_X1 U789 ( .A(KEYINPUT50), .ZN(n1105) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1097) );
INV_X1 U791 ( .A(G104), .ZN(n1107) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND2_X1 U793 ( .A1(KEYINPUT58), .A2(n1102), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1104), .B(KEYINPUT44), .Z(n1102) );
NAND2_X1 U795 ( .A1(KEYINPUT50), .A2(n1104), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1078), .A2(n1110), .ZN(G57) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U798 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND3_X1 U799 ( .A1(n1082), .A2(G472), .A3(KEYINPUT49), .ZN(n1113) );
XOR2_X1 U800 ( .A(n1115), .B(n1116), .Z(n1111) );
XOR2_X1 U801 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U802 ( .A1(KEYINPUT8), .A2(n1119), .ZN(n1117) );
NAND2_X1 U803 ( .A1(KEYINPUT29), .A2(n1120), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1078), .A2(n1121), .ZN(G54) );
XOR2_X1 U805 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U807 ( .A1(KEYINPUT38), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U808 ( .A(n1127), .B(n1128), .ZN(n1126) );
NAND2_X1 U809 ( .A1(KEYINPUT19), .A2(n1129), .ZN(n1127) );
NAND2_X1 U810 ( .A1(n1082), .A2(G469), .ZN(n1124) );
NOR2_X1 U811 ( .A1(n1078), .A2(n1130), .ZN(G51) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND3_X1 U814 ( .A1(n1082), .A2(G210), .A3(KEYINPUT2), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1001), .ZN(n1082) );
NOR2_X1 U816 ( .A1(n1065), .A2(n1051), .ZN(n1001) );
NAND4_X1 U817 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1051) );
AND4_X1 U818 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
NAND2_X1 U819 ( .A1(n1009), .A2(n1144), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U821 ( .A(KEYINPUT15), .B(n1147), .ZN(n1145) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1136) );
INV_X1 U823 ( .A(n1150), .ZN(n1148) );
NAND4_X1 U824 ( .A1(n1151), .A2(n1104), .A3(n1152), .A4(n1153), .ZN(n1065) );
NOR4_X1 U825 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n987), .ZN(n1153) );
AND3_X1 U826 ( .A1(n998), .A2(n1157), .A3(n1018), .ZN(n987) );
AND2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NAND3_X1 U828 ( .A1(n998), .A2(n1157), .A3(n1160), .ZN(n1104) );
NAND3_X1 U829 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1151) );
XOR2_X1 U830 ( .A(KEYINPUT17), .B(n1000), .Z(n1162) );
NAND2_X1 U831 ( .A1(n1164), .A2(n1165), .ZN(n1133) );
XOR2_X1 U832 ( .A(n1166), .B(KEYINPUT55), .Z(n1164) );
NOR2_X1 U833 ( .A1(KEYINPUT43), .A2(n1167), .ZN(n1131) );
NOR2_X1 U834 ( .A1(n1047), .A2(G952), .ZN(n1078) );
XOR2_X1 U835 ( .A(n1168), .B(n1169), .Z(G48) );
NOR2_X1 U836 ( .A1(KEYINPUT10), .A2(n1170), .ZN(n1169) );
NOR3_X1 U837 ( .A1(n1150), .A2(n1171), .A3(n1172), .ZN(n1168) );
NOR2_X1 U838 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
INV_X1 U839 ( .A(KEYINPUT0), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1025), .A2(n1175), .ZN(n1173) );
NOR2_X1 U841 ( .A1(KEYINPUT0), .A2(n1149), .ZN(n1171) );
NAND4_X1 U842 ( .A1(n1176), .A2(n1160), .A3(n1177), .A4(n1033), .ZN(n1150) );
XOR2_X1 U843 ( .A(n1178), .B(n1137), .Z(G45) );
NAND3_X1 U844 ( .A1(n1149), .A2(n1014), .A3(n1179), .ZN(n1137) );
AND3_X1 U845 ( .A1(n1177), .A2(n1180), .A3(n1038), .ZN(n1179) );
XOR2_X1 U846 ( .A(n1181), .B(G140), .Z(G42) );
NAND2_X1 U847 ( .A1(KEYINPUT34), .A2(n1143), .ZN(n1181) );
NAND3_X1 U848 ( .A1(n1160), .A2(n1182), .A3(n1183), .ZN(n1143) );
XOR2_X1 U849 ( .A(n1142), .B(n1184), .Z(G39) );
NAND2_X1 U850 ( .A1(KEYINPUT4), .A2(G137), .ZN(n1184) );
NAND3_X1 U851 ( .A1(n1176), .A2(n997), .A3(n1183), .ZN(n1142) );
AND3_X1 U852 ( .A1(n1149), .A2(n1033), .A3(n1009), .ZN(n1183) );
INV_X1 U853 ( .A(n1185), .ZN(n1009) );
XOR2_X1 U854 ( .A(G134), .B(n1186), .Z(G36) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1185), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1146), .B(KEYINPUT28), .Z(n1187) );
NAND3_X1 U857 ( .A1(n1014), .A2(n1018), .A3(n1149), .ZN(n1146) );
XOR2_X1 U858 ( .A(G131), .B(n1188), .Z(G33) );
NOR2_X1 U859 ( .A1(n1185), .A2(n1147), .ZN(n1188) );
NAND2_X1 U860 ( .A1(n1149), .A2(n1163), .ZN(n1147) );
NAND2_X1 U861 ( .A1(n1021), .A2(n1022), .ZN(n1185) );
XOR2_X1 U862 ( .A(n1034), .B(KEYINPUT46), .Z(n1021) );
NAND2_X1 U863 ( .A1(n1189), .A2(n1190), .ZN(G30) );
NAND2_X1 U864 ( .A1(G128), .A2(n1141), .ZN(n1190) );
XOR2_X1 U865 ( .A(KEYINPUT47), .B(n1191), .Z(n1189) );
NOR2_X1 U866 ( .A1(G128), .A2(n1141), .ZN(n1191) );
NAND3_X1 U867 ( .A1(n1176), .A2(n1149), .A3(n1192), .ZN(n1141) );
AND3_X1 U868 ( .A1(n1018), .A2(n1033), .A3(n1177), .ZN(n1192) );
NOR2_X1 U869 ( .A1(n1025), .A2(n1193), .ZN(n1149) );
XOR2_X1 U870 ( .A(n1156), .B(n1194), .Z(G3) );
NOR2_X1 U871 ( .A1(KEYINPUT23), .A2(n1120), .ZN(n1194) );
AND3_X1 U872 ( .A1(n997), .A2(n1157), .A3(n1014), .ZN(n1156) );
XOR2_X1 U873 ( .A(n1060), .B(n1140), .Z(G27) );
NAND4_X1 U874 ( .A1(n1000), .A2(n1177), .A3(n1160), .A4(n1195), .ZN(n1140) );
NOR3_X1 U875 ( .A1(n1196), .A2(n1197), .A3(n1193), .ZN(n1195) );
INV_X1 U876 ( .A(n1175), .ZN(n1193) );
NAND2_X1 U877 ( .A1(n1028), .A2(n1198), .ZN(n1175) );
NAND4_X1 U878 ( .A1(G953), .A2(G902), .A3(n1199), .A4(n1062), .ZN(n1198) );
INV_X1 U879 ( .A(G900), .ZN(n1062) );
XOR2_X1 U880 ( .A(n1159), .B(n1200), .Z(G24) );
XOR2_X1 U881 ( .A(KEYINPUT12), .B(G122), .Z(n1200) );
NAND4_X1 U882 ( .A1(n1201), .A2(n998), .A3(n1038), .A4(n1180), .ZN(n1159) );
NOR2_X1 U883 ( .A1(n1196), .A2(n1033), .ZN(n998) );
XNOR2_X1 U884 ( .A(G119), .B(n1158), .ZN(G21) );
NAND4_X1 U885 ( .A1(n1176), .A2(n1201), .A3(n997), .A4(n1033), .ZN(n1158) );
XNOR2_X1 U886 ( .A(n1155), .B(n1202), .ZN(G18) );
NAND2_X1 U887 ( .A1(KEYINPUT31), .A2(G116), .ZN(n1202) );
AND3_X1 U888 ( .A1(n1201), .A2(n1018), .A3(n1014), .ZN(n1155) );
NOR2_X1 U889 ( .A1(n1180), .A2(n1203), .ZN(n1018) );
XNOR2_X1 U890 ( .A(G113), .B(n1204), .ZN(G15) );
NAND2_X1 U891 ( .A1(n1163), .A2(n1201), .ZN(n1204) );
AND2_X1 U892 ( .A1(n1000), .A2(n1161), .ZN(n1201) );
INV_X1 U893 ( .A(n1205), .ZN(n1161) );
AND2_X1 U894 ( .A1(n1026), .A2(n1206), .ZN(n1000) );
XOR2_X1 U895 ( .A(n1207), .B(KEYINPUT13), .Z(n1026) );
AND2_X1 U896 ( .A1(n1160), .A2(n1014), .ZN(n1163) );
AND2_X1 U897 ( .A1(n1208), .A2(n1197), .ZN(n1014) );
INV_X1 U898 ( .A(n1033), .ZN(n1197) );
XOR2_X1 U899 ( .A(n1176), .B(KEYINPUT63), .Z(n1208) );
XOR2_X1 U900 ( .A(n1196), .B(KEYINPUT26), .Z(n1176) );
INV_X1 U901 ( .A(n1017), .ZN(n1160) );
NAND2_X1 U902 ( .A1(n1203), .A2(n1180), .ZN(n1017) );
XOR2_X1 U903 ( .A(G110), .B(n1154), .Z(G12) );
NOR2_X1 U904 ( .A1(n1012), .A2(n1209), .ZN(n1154) );
INV_X1 U905 ( .A(n1157), .ZN(n1209) );
NOR2_X1 U906 ( .A1(n1025), .A2(n1205), .ZN(n1157) );
NAND2_X1 U907 ( .A1(n1177), .A2(n1210), .ZN(n1205) );
NAND2_X1 U908 ( .A1(n1211), .A2(n1028), .ZN(n1210) );
NAND3_X1 U909 ( .A1(n1199), .A2(n1047), .A3(G952), .ZN(n1028) );
NAND3_X1 U910 ( .A1(G902), .A2(n1199), .A3(n1077), .ZN(n1211) );
NOR2_X1 U911 ( .A1(G898), .A2(n1047), .ZN(n1077) );
NAND2_X1 U912 ( .A1(G234), .A2(G237), .ZN(n1199) );
INV_X1 U913 ( .A(n994), .ZN(n1177) );
NAND2_X1 U914 ( .A1(n1034), .A2(n1022), .ZN(n994) );
NAND2_X1 U915 ( .A1(G214), .A2(n1212), .ZN(n1022) );
NAND2_X1 U916 ( .A1(n1213), .A2(n1135), .ZN(n1212) );
NAND2_X1 U917 ( .A1(n1214), .A2(n1215), .ZN(n1034) );
NAND2_X1 U918 ( .A1(G210), .A2(n1216), .ZN(n1215) );
NAND2_X1 U919 ( .A1(n1135), .A2(n1217), .ZN(n1216) );
OR2_X1 U920 ( .A1(n1213), .A2(n1218), .ZN(n1217) );
INV_X1 U921 ( .A(G237), .ZN(n1213) );
NAND3_X1 U922 ( .A1(n1219), .A2(n1135), .A3(n1218), .ZN(n1214) );
XNOR2_X1 U923 ( .A(n1220), .B(n1167), .ZN(n1218) );
XOR2_X1 U924 ( .A(n1074), .B(n1221), .Z(n1167) );
NOR2_X1 U925 ( .A1(KEYINPUT22), .A2(n1075), .ZN(n1221) );
XOR2_X1 U926 ( .A(n1222), .B(n1223), .Z(n1075) );
NAND2_X1 U927 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
NAND2_X1 U928 ( .A1(G113), .A2(n1226), .ZN(n1225) );
XOR2_X1 U929 ( .A(n1227), .B(KEYINPUT6), .Z(n1224) );
OR2_X1 U930 ( .A1(n1226), .A2(G113), .ZN(n1227) );
XNOR2_X1 U931 ( .A(G110), .B(G122), .ZN(n1074) );
XOR2_X1 U932 ( .A(n1228), .B(KEYINPUT1), .Z(n1220) );
NAND2_X1 U933 ( .A1(n1166), .A2(n1165), .ZN(n1228) );
NAND2_X1 U934 ( .A1(n1229), .A2(n1230), .ZN(n1165) );
NAND2_X1 U935 ( .A1(G224), .A2(n1047), .ZN(n1230) );
XOR2_X1 U936 ( .A(n1060), .B(n1231), .Z(n1229) );
NAND3_X1 U937 ( .A1(G224), .A2(n1047), .A3(n1232), .ZN(n1166) );
XOR2_X1 U938 ( .A(n1231), .B(G125), .Z(n1232) );
NAND2_X1 U939 ( .A1(G210), .A2(G237), .ZN(n1219) );
NAND2_X1 U940 ( .A1(n1233), .A2(n1036), .ZN(n1025) );
INV_X1 U941 ( .A(n1207), .ZN(n1036) );
XOR2_X1 U942 ( .A(n1234), .B(G469), .Z(n1207) );
NAND2_X1 U943 ( .A1(n1235), .A2(n1135), .ZN(n1234) );
XOR2_X1 U944 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U945 ( .A(KEYINPUT48), .B(n1238), .Z(n1237) );
NOR2_X1 U946 ( .A1(KEYINPUT32), .A2(n1128), .ZN(n1238) );
XNOR2_X1 U947 ( .A(n1122), .B(n1129), .ZN(n1236) );
XNOR2_X1 U948 ( .A(n1223), .B(n1057), .ZN(n1129) );
XOR2_X1 U949 ( .A(G128), .B(n1239), .Z(n1057) );
NOR2_X1 U950 ( .A1(KEYINPUT60), .A2(n1240), .ZN(n1239) );
XOR2_X1 U951 ( .A(n1170), .B(G143), .Z(n1240) );
XNOR2_X1 U952 ( .A(n1120), .B(n1241), .ZN(n1223) );
XOR2_X1 U953 ( .A(G107), .B(G104), .Z(n1241) );
XOR2_X1 U954 ( .A(n1242), .B(n1243), .Z(n1122) );
NAND2_X1 U955 ( .A1(G227), .A2(n1047), .ZN(n1242) );
XOR2_X1 U956 ( .A(KEYINPUT9), .B(n1027), .Z(n1233) );
INV_X1 U957 ( .A(n1206), .ZN(n1027) );
NAND2_X1 U958 ( .A1(G221), .A2(n1244), .ZN(n1206) );
NAND2_X1 U959 ( .A1(G234), .A2(n1135), .ZN(n1244) );
NAND3_X1 U960 ( .A1(n1182), .A2(n1033), .A3(n997), .ZN(n1012) );
NOR2_X1 U961 ( .A1(n1038), .A2(n1180), .ZN(n997) );
NAND2_X1 U962 ( .A1(n1245), .A2(n1041), .ZN(n1180) );
NAND2_X1 U963 ( .A1(G475), .A2(n1246), .ZN(n1041) );
NAND2_X1 U964 ( .A1(n1093), .A2(n1247), .ZN(n1246) );
XOR2_X1 U965 ( .A(KEYINPUT33), .B(n1039), .Z(n1245) );
AND3_X1 U966 ( .A1(n1247), .A2(n1248), .A3(n1093), .ZN(n1039) );
XOR2_X1 U967 ( .A(n1249), .B(n1250), .Z(n1093) );
XOR2_X1 U968 ( .A(G122), .B(G104), .Z(n1250) );
XNOR2_X1 U969 ( .A(n1251), .B(n1252), .ZN(n1249) );
NOR2_X1 U970 ( .A1(G113), .A2(KEYINPUT59), .ZN(n1252) );
NOR2_X1 U971 ( .A1(KEYINPUT53), .A2(n1253), .ZN(n1251) );
XOR2_X1 U972 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U973 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U974 ( .A1(KEYINPUT45), .A2(n1258), .ZN(n1257) );
XOR2_X1 U975 ( .A(G140), .B(n1259), .Z(n1258) );
NAND2_X1 U976 ( .A1(G214), .A2(n1260), .ZN(n1256) );
XOR2_X1 U977 ( .A(G131), .B(n1178), .Z(n1254) );
INV_X1 U978 ( .A(G475), .ZN(n1248) );
XOR2_X1 U979 ( .A(G902), .B(KEYINPUT18), .Z(n1247) );
INV_X1 U980 ( .A(n1203), .ZN(n1038) );
XOR2_X1 U981 ( .A(n1261), .B(G478), .Z(n1203) );
NAND2_X1 U982 ( .A1(n1089), .A2(n1135), .ZN(n1261) );
XNOR2_X1 U983 ( .A(n1262), .B(n1263), .ZN(n1089) );
NOR2_X1 U984 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U985 ( .A1(KEYINPUT25), .A2(n1266), .ZN(n1262) );
XOR2_X1 U986 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U987 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U988 ( .A(G107), .B(n1271), .Z(n1270) );
NOR2_X1 U989 ( .A1(G134), .A2(KEYINPUT62), .ZN(n1271) );
NOR2_X1 U990 ( .A1(G116), .A2(KEYINPUT36), .ZN(n1269) );
XOR2_X1 U991 ( .A(G122), .B(n1272), .Z(n1267) );
XOR2_X1 U992 ( .A(G143), .B(G128), .Z(n1272) );
NAND3_X1 U993 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1033) );
NAND2_X1 U994 ( .A1(n1276), .A2(n1081), .ZN(n1275) );
OR3_X1 U995 ( .A1(n1081), .A2(n1276), .A3(G902), .ZN(n1274) );
NOR2_X1 U996 ( .A1(n1265), .A2(G234), .ZN(n1276) );
INV_X1 U997 ( .A(G217), .ZN(n1265) );
XOR2_X1 U998 ( .A(n1277), .B(n1278), .Z(n1081) );
XNOR2_X1 U999 ( .A(n1259), .B(n1279), .ZN(n1278) );
XNOR2_X1 U1000 ( .A(n1243), .B(n1280), .ZN(n1279) );
NOR3_X1 U1001 ( .A1(n1281), .A2(KEYINPUT11), .A3(n1264), .ZN(n1280) );
NAND2_X1 U1002 ( .A1(G234), .A2(n1047), .ZN(n1264) );
INV_X1 U1003 ( .A(G221), .ZN(n1281) );
XOR2_X1 U1004 ( .A(G110), .B(G140), .Z(n1243) );
XOR2_X1 U1005 ( .A(n1060), .B(n1170), .Z(n1259) );
INV_X1 U1006 ( .A(G146), .ZN(n1170) );
INV_X1 U1007 ( .A(G125), .ZN(n1060) );
XOR2_X1 U1008 ( .A(n1282), .B(n1283), .Z(n1277) );
XOR2_X1 U1009 ( .A(G119), .B(n1284), .Z(n1283) );
NOR2_X1 U1010 ( .A1(G128), .A2(KEYINPUT24), .ZN(n1284) );
XNOR2_X1 U1011 ( .A(G137), .B(KEYINPUT14), .ZN(n1282) );
NAND2_X1 U1012 ( .A1(G217), .A2(G902), .ZN(n1273) );
INV_X1 U1013 ( .A(n1196), .ZN(n1182) );
NAND2_X1 U1014 ( .A1(n1285), .A2(n1286), .ZN(n1196) );
NAND2_X1 U1015 ( .A1(G472), .A2(n1042), .ZN(n1286) );
XOR2_X1 U1016 ( .A(n1287), .B(KEYINPUT42), .Z(n1285) );
OR2_X1 U1017 ( .A1(n1042), .A2(G472), .ZN(n1287) );
NAND2_X1 U1018 ( .A1(n1288), .A2(n1135), .ZN(n1042) );
INV_X1 U1019 ( .A(G902), .ZN(n1135) );
XOR2_X1 U1020 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1021 ( .A(n1114), .B(n1119), .Z(n1290) );
XOR2_X1 U1022 ( .A(n1231), .B(n1128), .Z(n1119) );
XNOR2_X1 U1023 ( .A(G131), .B(n1056), .ZN(n1128) );
XOR2_X1 U1024 ( .A(G134), .B(G137), .Z(n1056) );
XOR2_X1 U1025 ( .A(n1291), .B(n1292), .Z(n1231) );
NOR2_X1 U1026 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U1027 ( .A(n1295), .B(KEYINPUT21), .Z(n1294) );
NAND2_X1 U1028 ( .A1(n1296), .A2(n1178), .ZN(n1295) );
XOR2_X1 U1029 ( .A(KEYINPUT20), .B(n1297), .Z(n1296) );
NOR2_X1 U1030 ( .A1(n1178), .A2(n1297), .ZN(n1293) );
XOR2_X1 U1031 ( .A(G146), .B(KEYINPUT16), .Z(n1297) );
INV_X1 U1032 ( .A(G143), .ZN(n1178) );
XNOR2_X1 U1033 ( .A(G128), .B(KEYINPUT3), .ZN(n1291) );
XNOR2_X1 U1034 ( .A(G113), .B(n1226), .ZN(n1114) );
XOR2_X1 U1035 ( .A(G116), .B(G119), .Z(n1226) );
XOR2_X1 U1036 ( .A(n1120), .B(n1118), .Z(n1289) );
AND2_X1 U1037 ( .A1(G210), .A2(n1260), .ZN(n1118) );
AND2_X1 U1038 ( .A1(n1298), .A2(n1047), .ZN(n1260) );
INV_X1 U1039 ( .A(G953), .ZN(n1047) );
XOR2_X1 U1040 ( .A(KEYINPUT5), .B(G237), .Z(n1298) );
INV_X1 U1041 ( .A(G101), .ZN(n1120) );
endmodule


