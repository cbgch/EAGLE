//Key = 0000111010010001010110110000100111001010101101010111111011001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329;

XOR2_X1 U729 ( .A(G107), .B(n1006), .Z(G9) );
NOR2_X1 U730 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1009), .A2(n1010), .A3(G953), .A4(n1011), .ZN(n1008) );
NOR2_X1 U732 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U733 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR3_X1 U734 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR3_X1 U736 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR3_X1 U737 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1022) );
AND3_X1 U739 ( .A1(KEYINPUT53), .A2(n1027), .A3(n1029), .ZN(n1019) );
NOR4_X1 U740 ( .A1(n1030), .A2(n1021), .A3(n1031), .A4(n1024), .ZN(n1014) );
NOR2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U742 ( .A1(n1034), .A2(n1018), .ZN(n1033) );
NOR3_X1 U743 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
AND2_X1 U744 ( .A1(n1038), .A2(KEYINPUT27), .ZN(n1037) );
NOR3_X1 U745 ( .A1(KEYINPUT27), .A2(n1039), .A3(n1040), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1041), .A2(n1016), .ZN(n1032) );
NOR2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NAND3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1009) );
NAND2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
INV_X1 U751 ( .A(KEYINPUT53), .ZN(n1050) );
NAND4_X1 U752 ( .A1(n1051), .A2(n1038), .A3(n1052), .A4(n1029), .ZN(n1049) );
NOR2_X1 U753 ( .A1(n1018), .A2(n1031), .ZN(n1052) );
INV_X1 U754 ( .A(n1027), .ZN(n1031) );
INV_X1 U755 ( .A(n1053), .ZN(n1018) );
INV_X1 U756 ( .A(n1013), .ZN(n1051) );
NOR3_X1 U757 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U758 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1011) );
NOR4_X1 U759 ( .A1(n1058), .A2(n1059), .A3(n1024), .A4(n1060), .ZN(n1057) );
XNOR2_X1 U760 ( .A(n1061), .B(n1062), .ZN(n1060) );
XOR2_X1 U761 ( .A(n1063), .B(KEYINPUT12), .Z(n1062) );
XOR2_X1 U762 ( .A(n1064), .B(KEYINPUT50), .Z(n1058) );
NOR3_X1 U763 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1056) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1055) );
XOR2_X1 U765 ( .A(KEYINPUT61), .B(n1070), .Z(n1054) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1073), .B(KEYINPUT33), .Z(n1072) );
NAND2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XNOR2_X1 U769 ( .A(KEYINPUT17), .B(n1076), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1076), .ZN(n1071) );
INV_X1 U771 ( .A(n1077), .ZN(n1074) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR3_X1 U775 ( .A1(KEYINPUT59), .A2(n1084), .A3(n1085), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U777 ( .A(n1088), .ZN(n1087) );
NOR2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NOR2_X1 U779 ( .A1(G900), .A2(n1081), .ZN(n1089) );
NOR2_X1 U780 ( .A1(n1090), .A2(n1088), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1088) );
XOR2_X1 U782 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U783 ( .A(G134), .B(KEYINPUT60), .ZN(n1094) );
NAND2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U785 ( .A1(G140), .A2(n1097), .ZN(n1096) );
XOR2_X1 U786 ( .A(KEYINPUT51), .B(n1098), .Z(n1095) );
NOR2_X1 U787 ( .A1(G140), .A2(n1097), .ZN(n1098) );
XOR2_X1 U788 ( .A(n1099), .B(n1100), .Z(n1091) );
AND2_X1 U789 ( .A1(n1101), .A2(n1081), .ZN(n1090) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U791 ( .A(n1104), .ZN(n1103) );
NAND3_X1 U792 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G69) );
XOR2_X1 U793 ( .A(n1108), .B(KEYINPUT34), .Z(n1107) );
NAND3_X1 U794 ( .A1(n1109), .A2(n1110), .A3(G953), .ZN(n1108) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1109) );
NAND2_X1 U796 ( .A1(n1111), .A2(n1081), .ZN(n1106) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND3_X1 U798 ( .A1(n1113), .A2(G224), .A3(G953), .ZN(n1105) );
INV_X1 U799 ( .A(n1110), .ZN(n1113) );
NAND3_X1 U800 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1110) );
NAND2_X1 U801 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
XNOR2_X1 U803 ( .A(n1120), .B(n1121), .ZN(n1118) );
XNOR2_X1 U804 ( .A(KEYINPUT8), .B(KEYINPUT62), .ZN(n1120) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1114) );
INV_X1 U806 ( .A(n1119), .ZN(n1122) );
XOR2_X1 U807 ( .A(n1123), .B(KEYINPUT25), .Z(n1119) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U810 ( .A1(n1076), .A2(n1128), .ZN(n1127) );
NOR2_X1 U811 ( .A1(n1124), .A2(n1129), .ZN(G63) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U813 ( .A1(n1063), .A2(n1128), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1132), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1133), .B(n1134), .ZN(n1132) );
AND2_X1 U816 ( .A1(G475), .A2(n1135), .ZN(n1134) );
XNOR2_X1 U817 ( .A(G104), .B(n1136), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1124), .A2(n1137), .ZN(G57) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1128), .ZN(n1141) );
XNOR2_X1 U822 ( .A(G472), .B(KEYINPUT35), .ZN(n1142) );
NAND2_X1 U823 ( .A1(n1143), .A2(KEYINPUT20), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1144), .B(KEYINPUT11), .Z(n1143) );
NOR3_X1 U825 ( .A1(n1124), .A2(n1145), .A3(n1146), .ZN(G54) );
NOR2_X1 U826 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
AND2_X1 U828 ( .A1(n1151), .A2(KEYINPUT7), .ZN(n1150) );
NOR3_X1 U829 ( .A1(KEYINPUT7), .A2(n1151), .A3(n1152), .ZN(n1149) );
INV_X1 U830 ( .A(n1153), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n1154), .A2(n1153), .ZN(n1145) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1153) );
XOR2_X1 U833 ( .A(G143), .B(n1157), .Z(n1156) );
XOR2_X1 U834 ( .A(KEYINPUT9), .B(KEYINPUT41), .Z(n1157) );
XOR2_X1 U835 ( .A(n1158), .B(n1159), .Z(n1155) );
XNOR2_X1 U836 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1151), .A2(n1152), .ZN(n1154) );
INV_X1 U838 ( .A(KEYINPUT5), .ZN(n1152) );
NAND2_X1 U839 ( .A1(n1135), .A2(G469), .ZN(n1151) );
INV_X1 U840 ( .A(n1128), .ZN(n1135) );
NOR2_X1 U841 ( .A1(n1081), .A2(G952), .ZN(n1124) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(G51) );
XOR2_X1 U843 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U844 ( .A1(n1166), .A2(n1128), .ZN(n1165) );
NAND2_X1 U845 ( .A1(G902), .A2(n1167), .ZN(n1128) );
NAND2_X1 U846 ( .A1(n1048), .A2(n1046), .ZN(n1167) );
XNOR2_X1 U847 ( .A(n1102), .B(KEYINPUT42), .ZN(n1046) );
NOR4_X1 U848 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1102) );
INV_X1 U849 ( .A(n1172), .ZN(n1170) );
NOR2_X1 U850 ( .A1(n1112), .A2(n1104), .ZN(n1048) );
NAND4_X1 U851 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1104) );
NAND4_X1 U852 ( .A1(n1177), .A2(n1136), .A3(n1178), .A4(n1179), .ZN(n1112) );
NOR4_X1 U853 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1006), .ZN(n1179) );
AND4_X1 U854 ( .A1(n1043), .A2(n1025), .A3(n1028), .A4(n1183), .ZN(n1006) );
INV_X1 U855 ( .A(n1184), .ZN(n1183) );
NAND2_X1 U856 ( .A1(n1035), .A2(n1185), .ZN(n1178) );
NAND2_X1 U857 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U858 ( .A(n1188), .B(KEYINPUT18), .ZN(n1187) );
XOR2_X1 U859 ( .A(n1189), .B(KEYINPUT13), .Z(n1186) );
NAND4_X1 U860 ( .A1(n1190), .A2(n1191), .A3(n1028), .A4(n1192), .ZN(n1136) );
AND2_X1 U861 ( .A1(n1043), .A2(n1193), .ZN(n1192) );
NAND3_X1 U862 ( .A1(n1053), .A2(n1194), .A3(n1026), .ZN(n1177) );
NOR2_X1 U863 ( .A1(n1195), .A2(n1196), .ZN(n1164) );
XOR2_X1 U864 ( .A(KEYINPUT26), .B(n1197), .Z(n1196) );
NOR2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
AND2_X1 U866 ( .A1(n1199), .A2(n1198), .ZN(n1195) );
XNOR2_X1 U867 ( .A(n1200), .B(n1201), .ZN(n1199) );
NAND2_X1 U868 ( .A1(KEYINPUT63), .A2(n1202), .ZN(n1200) );
NOR2_X1 U869 ( .A1(G952), .A2(n1203), .ZN(n1162) );
XOR2_X1 U870 ( .A(n1081), .B(KEYINPUT16), .Z(n1203) );
XNOR2_X1 U871 ( .A(G146), .B(n1204), .ZN(G48) );
NAND2_X1 U872 ( .A1(KEYINPUT49), .A2(n1169), .ZN(n1204) );
AND2_X1 U873 ( .A1(n1205), .A2(n1193), .ZN(n1169) );
XOR2_X1 U874 ( .A(n1206), .B(n1172), .Z(G45) );
NAND4_X1 U875 ( .A1(n1207), .A2(n1208), .A3(n1035), .A4(n1209), .ZN(n1172) );
XOR2_X1 U876 ( .A(n1210), .B(G140), .Z(G42) );
NAND3_X1 U877 ( .A1(n1211), .A2(n1212), .A3(KEYINPUT15), .ZN(n1210) );
NAND2_X1 U878 ( .A1(n1168), .A2(n1213), .ZN(n1212) );
INV_X1 U879 ( .A(KEYINPUT44), .ZN(n1213) );
NOR2_X1 U880 ( .A1(n1214), .A2(n1016), .ZN(n1168) );
INV_X1 U881 ( .A(n1038), .ZN(n1016) );
NAND3_X1 U882 ( .A1(n1038), .A2(n1214), .A3(KEYINPUT44), .ZN(n1211) );
NAND4_X1 U883 ( .A1(n1029), .A2(n1026), .A3(n1043), .A4(n1215), .ZN(n1214) );
XOR2_X1 U884 ( .A(G137), .B(n1171), .Z(G39) );
AND3_X1 U885 ( .A1(n1205), .A2(n1027), .A3(n1038), .ZN(n1171) );
XNOR2_X1 U886 ( .A(G134), .B(n1173), .ZN(G36) );
NAND3_X1 U887 ( .A1(n1208), .A2(n1025), .A3(n1038), .ZN(n1173) );
XNOR2_X1 U888 ( .A(G131), .B(n1174), .ZN(G33) );
NAND3_X1 U889 ( .A1(n1208), .A2(n1026), .A3(n1038), .ZN(n1174) );
NOR2_X1 U890 ( .A1(n1039), .A2(n1065), .ZN(n1038) );
INV_X1 U891 ( .A(n1040), .ZN(n1065) );
AND4_X1 U892 ( .A1(n1190), .A2(n1043), .A3(n1024), .A4(n1215), .ZN(n1208) );
NAND2_X1 U893 ( .A1(n1216), .A2(n1217), .ZN(G30) );
OR2_X1 U894 ( .A1(n1176), .A2(G128), .ZN(n1217) );
XOR2_X1 U895 ( .A(n1218), .B(KEYINPUT0), .Z(n1216) );
NAND2_X1 U896 ( .A1(G128), .A2(n1176), .ZN(n1218) );
NAND3_X1 U897 ( .A1(n1025), .A2(n1035), .A3(n1205), .ZN(n1176) );
AND4_X1 U898 ( .A1(n1043), .A2(n1024), .A3(n1021), .A4(n1215), .ZN(n1205) );
INV_X1 U899 ( .A(n1190), .ZN(n1021) );
XOR2_X1 U900 ( .A(G101), .B(n1182), .Z(G3) );
AND3_X1 U901 ( .A1(n1194), .A2(n1043), .A3(n1027), .ZN(n1182) );
XOR2_X1 U902 ( .A(n1097), .B(n1175), .Z(G27) );
NAND4_X1 U903 ( .A1(n1029), .A2(n1193), .A3(n1053), .A4(n1215), .ZN(n1175) );
NAND2_X1 U904 ( .A1(n1013), .A2(n1219), .ZN(n1215) );
NAND4_X1 U905 ( .A1(G902), .A2(n1220), .A3(n1221), .A4(n1083), .ZN(n1219) );
INV_X1 U906 ( .A(G900), .ZN(n1083) );
XOR2_X1 U907 ( .A(KEYINPUT29), .B(G953), .Z(n1220) );
AND2_X1 U908 ( .A1(n1026), .A2(n1035), .ZN(n1193) );
XOR2_X1 U909 ( .A(n1222), .B(n1181), .Z(G24) );
AND3_X1 U910 ( .A1(n1207), .A2(n1053), .A3(n1223), .ZN(n1181) );
NOR3_X1 U911 ( .A1(n1184), .A2(n1224), .A3(n1024), .ZN(n1223) );
NAND2_X1 U912 ( .A1(KEYINPUT31), .A2(n1225), .ZN(n1222) );
XNOR2_X1 U913 ( .A(G119), .B(n1226), .ZN(G21) );
NAND2_X1 U914 ( .A1(n1188), .A2(n1035), .ZN(n1226) );
AND3_X1 U915 ( .A1(n1027), .A2(n1053), .A3(n1227), .ZN(n1188) );
NOR3_X1 U916 ( .A1(n1028), .A2(n1228), .A3(n1190), .ZN(n1227) );
XOR2_X1 U917 ( .A(G116), .B(n1180), .Z(G18) );
AND3_X1 U918 ( .A1(n1194), .A2(n1025), .A3(n1053), .ZN(n1180) );
NOR2_X1 U919 ( .A1(n1207), .A2(n1224), .ZN(n1025) );
XOR2_X1 U920 ( .A(n1229), .B(n1230), .Z(G15) );
XOR2_X1 U921 ( .A(KEYINPUT23), .B(G113), .Z(n1230) );
NAND4_X1 U922 ( .A1(n1026), .A2(n1053), .A3(n1231), .A4(n1232), .ZN(n1229) );
OR2_X1 U923 ( .A1(n1194), .A2(KEYINPUT48), .ZN(n1232) );
NOR2_X1 U924 ( .A1(n1184), .A2(n1028), .ZN(n1194) );
NAND3_X1 U925 ( .A1(n1190), .A2(n1191), .A3(n1035), .ZN(n1184) );
NAND2_X1 U926 ( .A1(KEYINPUT48), .A2(n1233), .ZN(n1231) );
NAND4_X1 U927 ( .A1(n1228), .A2(n1035), .A3(n1190), .A4(n1024), .ZN(n1233) );
INV_X1 U928 ( .A(n1234), .ZN(n1035) );
INV_X1 U929 ( .A(n1191), .ZN(n1228) );
NOR2_X1 U930 ( .A1(n1044), .A2(n1067), .ZN(n1053) );
INV_X1 U931 ( .A(n1045), .ZN(n1067) );
AND2_X1 U932 ( .A1(n1224), .A2(n1207), .ZN(n1026) );
INV_X1 U933 ( .A(n1209), .ZN(n1224) );
XOR2_X1 U934 ( .A(n1235), .B(n1236), .Z(G12) );
XOR2_X1 U935 ( .A(KEYINPUT30), .B(G110), .Z(n1236) );
NOR2_X1 U936 ( .A1(n1234), .A2(n1189), .ZN(n1235) );
NAND4_X1 U937 ( .A1(n1029), .A2(n1027), .A3(n1043), .A4(n1191), .ZN(n1189) );
NAND2_X1 U938 ( .A1(n1013), .A2(n1237), .ZN(n1191) );
NAND4_X1 U939 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1117), .ZN(n1237) );
INV_X1 U940 ( .A(G898), .ZN(n1117) );
NAND3_X1 U941 ( .A1(n1221), .A2(n1081), .A3(G952), .ZN(n1013) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1221) );
AND2_X1 U943 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U944 ( .A1(G221), .A2(n1238), .ZN(n1045) );
XOR2_X1 U945 ( .A(n1064), .B(KEYINPUT47), .Z(n1044) );
XOR2_X1 U946 ( .A(n1239), .B(G469), .Z(n1064) );
NAND2_X1 U947 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U948 ( .A(n1242), .B(n1243), .Z(n1240) );
XNOR2_X1 U949 ( .A(n1244), .B(KEYINPUT46), .ZN(n1243) );
NAND2_X1 U950 ( .A1(n1245), .A2(KEYINPUT52), .ZN(n1244) );
XOR2_X1 U951 ( .A(n1161), .B(n1246), .Z(n1245) );
NOR2_X1 U952 ( .A1(KEYINPUT1), .A2(n1247), .ZN(n1246) );
XOR2_X1 U953 ( .A(KEYINPUT41), .B(G140), .Z(n1247) );
XNOR2_X1 U954 ( .A(G110), .B(n1248), .ZN(n1161) );
NOR2_X1 U955 ( .A1(G953), .A2(n1082), .ZN(n1248) );
INV_X1 U956 ( .A(G227), .ZN(n1082) );
XOR2_X1 U957 ( .A(n1158), .B(n1100), .Z(n1242) );
XOR2_X1 U958 ( .A(G146), .B(G143), .Z(n1100) );
XOR2_X1 U959 ( .A(n1249), .B(n1250), .Z(n1158) );
XOR2_X1 U960 ( .A(KEYINPUT37), .B(G104), .Z(n1250) );
XOR2_X1 U961 ( .A(n1251), .B(n1252), .Z(n1249) );
NOR2_X1 U962 ( .A1(n1209), .A2(n1207), .ZN(n1027) );
XNOR2_X1 U963 ( .A(n1059), .B(KEYINPUT54), .ZN(n1207) );
XNOR2_X1 U964 ( .A(n1253), .B(G475), .ZN(n1059) );
NAND2_X1 U965 ( .A1(n1241), .A2(n1133), .ZN(n1253) );
NAND2_X1 U966 ( .A1(n1254), .A2(n1255), .ZN(n1133) );
OR2_X1 U967 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U968 ( .A(n1258), .B(KEYINPUT10), .Z(n1254) );
NAND2_X1 U969 ( .A1(n1257), .A2(n1256), .ZN(n1258) );
XNOR2_X1 U970 ( .A(n1259), .B(n1260), .ZN(n1256) );
NOR2_X1 U971 ( .A1(G122), .A2(KEYINPUT39), .ZN(n1260) );
XNOR2_X1 U972 ( .A(G104), .B(G113), .ZN(n1259) );
XNOR2_X1 U973 ( .A(n1261), .B(n1262), .ZN(n1257) );
XOR2_X1 U974 ( .A(n1263), .B(G131), .Z(n1261) );
NAND2_X1 U975 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND4_X1 U976 ( .A1(G214), .A2(G143), .A3(n1266), .A4(n1081), .ZN(n1265) );
NAND2_X1 U977 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
NAND3_X1 U978 ( .A1(n1266), .A2(n1081), .A3(G214), .ZN(n1268) );
XOR2_X1 U979 ( .A(KEYINPUT19), .B(G143), .Z(n1267) );
NAND2_X1 U980 ( .A1(n1269), .A2(n1270), .ZN(n1209) );
NAND2_X1 U981 ( .A1(n1061), .A2(n1063), .ZN(n1270) );
XOR2_X1 U982 ( .A(KEYINPUT36), .B(n1271), .Z(n1269) );
NOR2_X1 U983 ( .A1(n1061), .A2(n1063), .ZN(n1271) );
INV_X1 U984 ( .A(G478), .ZN(n1063) );
NOR2_X1 U985 ( .A1(n1272), .A2(n1131), .ZN(n1061) );
XNOR2_X1 U986 ( .A(n1273), .B(n1274), .ZN(n1131) );
NOR2_X1 U987 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR2_X1 U988 ( .A1(KEYINPUT38), .A2(n1277), .ZN(n1276) );
AND2_X1 U989 ( .A1(KEYINPUT45), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U990 ( .A(n1278), .B(n1279), .ZN(n1277) );
XNOR2_X1 U991 ( .A(G107), .B(n1280), .ZN(n1279) );
NAND2_X1 U992 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U993 ( .A1(G128), .A2(n1283), .ZN(n1282) );
NAND2_X1 U994 ( .A1(KEYINPUT43), .A2(n1284), .ZN(n1283) );
NAND2_X1 U995 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1284) );
NAND2_X1 U996 ( .A1(n1285), .A2(n1206), .ZN(n1281) );
INV_X1 U997 ( .A(G143), .ZN(n1206) );
NAND2_X1 U998 ( .A1(KEYINPUT56), .A2(n1286), .ZN(n1285) );
NAND2_X1 U999 ( .A1(KEYINPUT43), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U1000 ( .A(G116), .B(n1288), .ZN(n1278) );
XOR2_X1 U1001 ( .A(G134), .B(G122), .Z(n1288) );
NAND2_X1 U1002 ( .A1(G217), .A2(n1289), .ZN(n1273) );
XOR2_X1 U1003 ( .A(KEYINPUT22), .B(n1241), .Z(n1272) );
NOR2_X1 U1004 ( .A1(n1024), .A2(n1190), .ZN(n1029) );
XOR2_X1 U1005 ( .A(n1076), .B(n1290), .Z(n1190) );
NOR2_X1 U1006 ( .A1(KEYINPUT2), .A2(n1077), .ZN(n1290) );
NAND2_X1 U1007 ( .A1(n1241), .A2(n1291), .ZN(n1077) );
INV_X1 U1008 ( .A(n1126), .ZN(n1291) );
XOR2_X1 U1009 ( .A(n1292), .B(n1293), .Z(n1126) );
XOR2_X1 U1010 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1011 ( .A(G119), .B(G110), .ZN(n1295) );
NAND2_X1 U1012 ( .A1(n1289), .A2(G221), .ZN(n1294) );
AND2_X1 U1013 ( .A1(G234), .A2(n1081), .ZN(n1289) );
XNOR2_X1 U1014 ( .A(n1262), .B(n1296), .ZN(n1292) );
XNOR2_X1 U1015 ( .A(n1097), .B(n1160), .ZN(n1262) );
XNOR2_X1 U1016 ( .A(n1297), .B(G146), .ZN(n1160) );
INV_X1 U1017 ( .A(G140), .ZN(n1297) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1238), .ZN(n1076) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1298), .ZN(n1238) );
INV_X1 U1020 ( .A(n1028), .ZN(n1024) );
XOR2_X1 U1021 ( .A(n1299), .B(G472), .Z(n1028) );
NAND2_X1 U1022 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U1023 ( .A(KEYINPUT40), .B(n1302), .Z(n1301) );
INV_X1 U1024 ( .A(n1241), .ZN(n1302) );
XOR2_X1 U1025 ( .A(n1144), .B(n1303), .Z(n1300) );
INV_X1 U1026 ( .A(n1138), .ZN(n1303) );
XOR2_X1 U1027 ( .A(n1304), .B(n1305), .Z(n1138) );
AND3_X1 U1028 ( .A1(G210), .A2(n1081), .A3(n1266), .ZN(n1305) );
INV_X1 U1029 ( .A(G101), .ZN(n1304) );
XOR2_X1 U1030 ( .A(n1306), .B(n1307), .Z(n1144) );
XOR2_X1 U1031 ( .A(n1251), .B(n1308), .Z(n1306) );
XOR2_X1 U1032 ( .A(n1309), .B(n1310), .Z(n1251) );
XOR2_X1 U1033 ( .A(KEYINPUT57), .B(KEYINPUT28), .Z(n1310) );
XOR2_X1 U1034 ( .A(n1099), .B(n1311), .Z(n1309) );
NOR2_X1 U1035 ( .A1(G134), .A2(KEYINPUT55), .ZN(n1311) );
XNOR2_X1 U1036 ( .A(G131), .B(n1296), .ZN(n1099) );
XNOR2_X1 U1037 ( .A(G137), .B(n1287), .ZN(n1296) );
INV_X1 U1038 ( .A(G128), .ZN(n1287) );
NAND2_X1 U1039 ( .A1(n1040), .A2(n1039), .ZN(n1234) );
NAND3_X1 U1040 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1039) );
INV_X1 U1041 ( .A(n1066), .ZN(n1314) );
NOR2_X1 U1042 ( .A1(n1069), .A2(n1068), .ZN(n1066) );
OR2_X1 U1043 ( .A1(n1068), .A2(KEYINPUT4), .ZN(n1313) );
NAND3_X1 U1044 ( .A1(n1068), .A2(n1069), .A3(KEYINPUT4), .ZN(n1312) );
NAND2_X1 U1045 ( .A1(n1315), .A2(n1241), .ZN(n1069) );
XOR2_X1 U1046 ( .A(n1298), .B(KEYINPUT24), .Z(n1241) );
XOR2_X1 U1047 ( .A(n1202), .B(n1316), .Z(n1315) );
XNOR2_X1 U1048 ( .A(n1198), .B(n1201), .ZN(n1316) );
AND2_X1 U1049 ( .A1(G224), .A2(n1081), .ZN(n1201) );
INV_X1 U1050 ( .A(G953), .ZN(n1081) );
XOR2_X1 U1051 ( .A(n1317), .B(n1121), .Z(n1198) );
XOR2_X1 U1052 ( .A(n1318), .B(n1319), .Z(n1121) );
XOR2_X1 U1053 ( .A(n1320), .B(n1252), .Z(n1319) );
XOR2_X1 U1054 ( .A(G101), .B(G107), .Z(n1252) );
NOR2_X1 U1055 ( .A1(G104), .A2(KEYINPUT3), .ZN(n1320) );
NAND2_X1 U1056 ( .A1(n1321), .A2(n1322), .ZN(n1318) );
NAND2_X1 U1057 ( .A1(n1307), .A2(n1323), .ZN(n1322) );
INV_X1 U1058 ( .A(KEYINPUT58), .ZN(n1323) );
XOR2_X1 U1059 ( .A(G113), .B(n1324), .Z(n1307) );
NAND3_X1 U1060 ( .A1(G113), .A2(n1324), .A3(KEYINPUT58), .ZN(n1321) );
XOR2_X1 U1061 ( .A(G116), .B(G119), .Z(n1324) );
NAND2_X1 U1062 ( .A1(n1325), .A2(KEYINPUT6), .ZN(n1317) );
XOR2_X1 U1063 ( .A(n1123), .B(KEYINPUT32), .Z(n1325) );
XOR2_X1 U1064 ( .A(G110), .B(n1225), .Z(n1123) );
INV_X1 U1065 ( .A(G122), .ZN(n1225) );
XOR2_X1 U1066 ( .A(n1326), .B(n1308), .Z(n1202) );
NOR2_X1 U1067 ( .A1(KEYINPUT21), .A2(n1327), .ZN(n1308) );
XOR2_X1 U1068 ( .A(G143), .B(n1328), .Z(n1327) );
NOR2_X1 U1069 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1328) );
XOR2_X1 U1070 ( .A(n1097), .B(G128), .Z(n1326) );
INV_X1 U1071 ( .A(G125), .ZN(n1097) );
INV_X1 U1072 ( .A(n1166), .ZN(n1068) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1329), .ZN(n1166) );
NAND2_X1 U1074 ( .A1(G214), .A2(n1329), .ZN(n1040) );
NAND2_X1 U1075 ( .A1(n1266), .A2(n1298), .ZN(n1329) );
INV_X1 U1076 ( .A(G902), .ZN(n1298) );
INV_X1 U1077 ( .A(G237), .ZN(n1266) );
endmodule


