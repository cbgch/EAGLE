//Key = 1111001101111100000101111110010011111110001110100110010111011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;

XOR2_X1 U750 ( .A(G107), .B(n1035), .Z(G9) );
NOR2_X1 U751 ( .A1(n1036), .A2(n1037), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1037) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR3_X1 U758 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1049) );
NOR2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR3_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1052) );
XOR2_X1 U763 ( .A(KEYINPUT50), .B(n1063), .Z(n1060) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1051) );
XOR2_X1 U765 ( .A(n1061), .B(KEYINPUT51), .Z(n1064) );
NOR3_X1 U766 ( .A1(n1061), .A2(n1066), .A3(n1067), .ZN(n1047) );
NOR3_X1 U767 ( .A1(n1055), .A2(n1068), .A3(n1069), .ZN(n1067) );
NOR2_X1 U768 ( .A1(KEYINPUT52), .A2(n1070), .ZN(n1069) );
NOR2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
AND2_X1 U770 ( .A1(n1073), .A2(KEYINPUT52), .ZN(n1072) );
NOR4_X1 U771 ( .A1(n1074), .A2(n1050), .A3(n1055), .A4(n1061), .ZN(n1043) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR3_X1 U773 ( .A1(n1038), .A2(G953), .A3(G952), .ZN(n1036) );
AND4_X1 U774 ( .A1(n1077), .A2(n1059), .A3(n1078), .A4(n1079), .ZN(n1038) );
NOR4_X1 U775 ( .A1(n1080), .A2(n1081), .A3(n1050), .A4(n1062), .ZN(n1079) );
INV_X1 U776 ( .A(n1082), .ZN(n1050) );
XNOR2_X1 U777 ( .A(n1083), .B(n1084), .ZN(n1081) );
XOR2_X1 U778 ( .A(KEYINPUT35), .B(G478), .Z(n1084) );
XOR2_X1 U779 ( .A(n1085), .B(n1086), .Z(n1080) );
NAND2_X1 U780 ( .A1(KEYINPUT37), .A2(n1087), .ZN(n1085) );
NOR2_X1 U781 ( .A1(n1063), .A2(n1088), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1077) );
XOR2_X1 U783 ( .A(n1091), .B(KEYINPUT34), .Z(n1089) );
XOR2_X1 U784 ( .A(n1092), .B(n1093), .Z(G72) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND3_X1 U787 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1092) );
NAND3_X1 U788 ( .A1(n1101), .A2(n1095), .A3(n1102), .ZN(n1100) );
NAND2_X1 U789 ( .A1(KEYINPUT33), .A2(n1103), .ZN(n1102) );
NAND2_X1 U790 ( .A1(KEYINPUT9), .A2(n1104), .ZN(n1103) );
OR2_X1 U791 ( .A1(n1105), .A2(KEYINPUT33), .ZN(n1099) );
NAND3_X1 U792 ( .A1(n1105), .A2(n1106), .A3(KEYINPUT33), .ZN(n1098) );
NAND3_X1 U793 ( .A1(n1101), .A2(n1095), .A3(KEYINPUT9), .ZN(n1106) );
INV_X1 U794 ( .A(n1104), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
NAND2_X1 U796 ( .A1(G953), .A2(n1097), .ZN(n1108) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1107) );
XOR2_X1 U798 ( .A(n1111), .B(G125), .Z(n1110) );
NAND2_X1 U799 ( .A1(KEYINPUT0), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U800 ( .A(KEYINPUT61), .B(n1113), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(G69) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1095), .ZN(n1115) );
AND2_X1 U803 ( .A1(G224), .A2(G898), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1117), .A2(KEYINPUT24), .ZN(n1114) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR3_X1 U806 ( .A1(n1120), .A2(KEYINPUT20), .A3(G953), .ZN(n1119) );
INV_X1 U807 ( .A(n1121), .ZN(n1120) );
NAND3_X1 U808 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1118) );
XOR2_X1 U809 ( .A(KEYINPUT11), .B(n1125), .Z(n1124) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U811 ( .A1(n1128), .A2(G953), .ZN(n1123) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1126), .ZN(n1122) );
XNOR2_X1 U813 ( .A(n1129), .B(n1130), .ZN(n1127) );
NAND2_X1 U814 ( .A1(KEYINPUT3), .A2(n1131), .ZN(n1129) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U816 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1132), .A2(n1138), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1083), .A2(n1139), .A3(n1140), .ZN(n1138) );
NOR3_X1 U820 ( .A1(n1141), .A2(n1142), .A3(n1137), .ZN(n1140) );
INV_X1 U821 ( .A(n1143), .ZN(n1141) );
NOR2_X1 U822 ( .A1(n1144), .A2(n1143), .ZN(n1139) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1142), .ZN(n1144) );
INV_X1 U824 ( .A(G478), .ZN(n1142) );
NOR2_X1 U825 ( .A1(n1132), .A2(n1146), .ZN(G60) );
NOR3_X1 U826 ( .A1(n1086), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR3_X1 U827 ( .A1(n1149), .A2(n1087), .A3(n1137), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1087), .ZN(n1150) );
INV_X1 U830 ( .A(G475), .ZN(n1087) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(G6) );
NOR2_X1 U832 ( .A1(n1132), .A2(n1154), .ZN(G57) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U834 ( .A1(KEYINPUT54), .A2(n1157), .ZN(n1155) );
XOR2_X1 U835 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U836 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U837 ( .A1(n1162), .A2(n1137), .ZN(n1160) );
INV_X1 U838 ( .A(G472), .ZN(n1162) );
XNOR2_X1 U839 ( .A(n1163), .B(n1164), .ZN(n1158) );
NOR2_X1 U840 ( .A1(n1132), .A2(n1165), .ZN(G54) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U843 ( .A1(KEYINPUT8), .A2(n1113), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1170), .A2(n1137), .ZN(n1168) );
INV_X1 U845 ( .A(G469), .ZN(n1170) );
NOR2_X1 U846 ( .A1(n1132), .A2(n1171), .ZN(G51) );
XOR2_X1 U847 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U848 ( .A1(n1091), .A2(n1137), .ZN(n1173) );
NAND2_X1 U849 ( .A1(G902), .A2(n1040), .ZN(n1137) );
INV_X1 U850 ( .A(n1145), .ZN(n1040) );
NOR2_X1 U851 ( .A1(n1121), .A2(n1101), .ZN(n1145) );
NAND4_X1 U852 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1101) );
NOR4_X1 U853 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR2_X1 U854 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
INV_X1 U855 ( .A(KEYINPUT43), .ZN(n1183) );
NOR2_X1 U856 ( .A1(n1184), .A2(n1185), .ZN(n1180) );
INV_X1 U857 ( .A(KEYINPUT13), .ZN(n1185) );
NOR3_X1 U858 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1179) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR3_X1 U860 ( .A1(n1070), .A2(KEYINPUT43), .A3(n1191), .ZN(n1190) );
NOR3_X1 U861 ( .A1(n1192), .A2(KEYINPUT13), .A3(n1046), .ZN(n1189) );
INV_X1 U862 ( .A(n1193), .ZN(n1046) );
INV_X1 U863 ( .A(n1061), .ZN(n1187) );
NOR3_X1 U864 ( .A1(n1194), .A2(n1191), .A3(n1192), .ZN(n1178) );
NAND3_X1 U865 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
XOR2_X1 U866 ( .A(n1198), .B(KEYINPUT60), .Z(n1197) );
NAND2_X1 U867 ( .A1(KEYINPUT53), .A2(n1186), .ZN(n1196) );
NAND2_X1 U868 ( .A1(n1199), .A2(n1200), .ZN(n1195) );
INV_X1 U869 ( .A(KEYINPUT53), .ZN(n1200) );
OR2_X1 U870 ( .A1(n1201), .A2(n1065), .ZN(n1199) );
AND3_X1 U871 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1176) );
NAND2_X1 U872 ( .A1(n1205), .A2(n1206), .ZN(n1121) );
NOR4_X1 U873 ( .A1(n1035), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1206) );
INV_X1 U874 ( .A(n1210), .ZN(n1208) );
AND3_X1 U875 ( .A1(n1082), .A2(n1075), .A3(n1211), .ZN(n1035) );
AND4_X1 U876 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1153), .ZN(n1205) );
NAND3_X1 U877 ( .A1(n1211), .A2(n1082), .A3(n1076), .ZN(n1153) );
NAND3_X1 U878 ( .A1(n1215), .A2(n1216), .A3(KEYINPUT56), .ZN(n1172) );
NAND2_X1 U879 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
INV_X1 U880 ( .A(KEYINPUT5), .ZN(n1218) );
XOR2_X1 U881 ( .A(n1219), .B(n1220), .Z(n1217) );
NAND2_X1 U882 ( .A1(KEYINPUT12), .A2(n1221), .ZN(n1220) );
NAND3_X1 U883 ( .A1(n1222), .A2(n1221), .A3(KEYINPUT5), .ZN(n1215) );
NAND2_X1 U884 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
NAND2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U886 ( .A(KEYINPUT62), .B(n1227), .Z(n1223) );
NOR2_X1 U887 ( .A1(n1226), .A2(n1225), .ZN(n1227) );
XNOR2_X1 U888 ( .A(n1228), .B(n1164), .ZN(n1225) );
NAND2_X1 U889 ( .A1(KEYINPUT49), .A2(n1229), .ZN(n1228) );
XOR2_X1 U890 ( .A(n1219), .B(KEYINPUT12), .Z(n1222) );
NOR2_X1 U891 ( .A1(n1095), .A2(G952), .ZN(n1132) );
XOR2_X1 U892 ( .A(n1230), .B(n1231), .Z(G48) );
NAND4_X1 U893 ( .A1(KEYINPUT10), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1231) );
NOR2_X1 U894 ( .A1(n1198), .A2(n1191), .ZN(n1233) );
XOR2_X1 U895 ( .A(n1174), .B(n1235), .Z(G45) );
NAND2_X1 U896 ( .A1(KEYINPUT57), .A2(G143), .ZN(n1235) );
NAND4_X1 U897 ( .A1(n1057), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1174) );
NOR2_X1 U898 ( .A1(n1070), .A2(n1186), .ZN(n1238) );
INV_X1 U899 ( .A(n1073), .ZN(n1070) );
XNOR2_X1 U900 ( .A(G140), .B(n1175), .ZN(G42) );
NAND3_X1 U901 ( .A1(n1076), .A2(n1068), .A3(n1239), .ZN(n1175) );
XNOR2_X1 U902 ( .A(G137), .B(n1184), .ZN(G39) );
NAND3_X1 U903 ( .A1(n1234), .A2(n1193), .A3(n1239), .ZN(n1184) );
XOR2_X1 U904 ( .A(n1202), .B(n1240), .Z(G36) );
NAND2_X1 U905 ( .A1(KEYINPUT32), .A2(G134), .ZN(n1240) );
NAND3_X1 U906 ( .A1(n1073), .A2(n1075), .A3(n1239), .ZN(n1202) );
XNOR2_X1 U907 ( .A(n1182), .B(n1241), .ZN(G33) );
NOR2_X1 U908 ( .A1(KEYINPUT63), .A2(n1242), .ZN(n1241) );
NAND3_X1 U909 ( .A1(n1073), .A2(n1076), .A3(n1239), .ZN(n1182) );
NOR2_X1 U910 ( .A1(n1186), .A2(n1061), .ZN(n1239) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1059), .ZN(n1061) );
INV_X1 U912 ( .A(n1058), .ZN(n1243) );
INV_X1 U913 ( .A(n1232), .ZN(n1186) );
NOR2_X1 U914 ( .A1(n1065), .A2(n1244), .ZN(n1232) );
INV_X1 U915 ( .A(n1201), .ZN(n1244) );
XNOR2_X1 U916 ( .A(G128), .B(n1204), .ZN(G30) );
NAND4_X1 U917 ( .A1(n1245), .A2(n1201), .A3(n1057), .A4(n1246), .ZN(n1204) );
NOR2_X1 U918 ( .A1(n1247), .A2(n1192), .ZN(n1246) );
NAND2_X1 U919 ( .A1(n1248), .A2(n1249), .ZN(G3) );
NAND2_X1 U920 ( .A1(G101), .A2(n1214), .ZN(n1249) );
XOR2_X1 U921 ( .A(n1250), .B(KEYINPUT14), .Z(n1248) );
OR2_X1 U922 ( .A1(n1214), .A2(G101), .ZN(n1250) );
NAND3_X1 U923 ( .A1(n1193), .A2(n1211), .A3(n1073), .ZN(n1214) );
XOR2_X1 U924 ( .A(n1229), .B(n1203), .Z(G27) );
NAND4_X1 U925 ( .A1(n1057), .A2(n1201), .A3(n1068), .A4(n1251), .ZN(n1203) );
NOR2_X1 U926 ( .A1(n1055), .A2(n1191), .ZN(n1251) );
INV_X1 U927 ( .A(n1076), .ZN(n1191) );
INV_X1 U928 ( .A(n1071), .ZN(n1055) );
NAND2_X1 U929 ( .A1(n1042), .A2(n1252), .ZN(n1201) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1253), .A4(n1097), .ZN(n1252) );
INV_X1 U931 ( .A(G900), .ZN(n1097) );
INV_X1 U932 ( .A(G125), .ZN(n1229) );
XNOR2_X1 U933 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1254), .A2(n1082), .A3(n1237), .A4(n1236), .ZN(n1213) );
NOR2_X1 U935 ( .A1(n1255), .A2(n1256), .ZN(n1082) );
XNOR2_X1 U936 ( .A(n1212), .B(n1257), .ZN(G21) );
XOR2_X1 U937 ( .A(KEYINPUT30), .B(G119), .Z(n1257) );
NAND3_X1 U938 ( .A1(n1254), .A2(n1193), .A3(n1234), .ZN(n1212) );
INV_X1 U939 ( .A(n1192), .ZN(n1234) );
NAND2_X1 U940 ( .A1(n1256), .A2(n1255), .ZN(n1192) );
INV_X1 U941 ( .A(n1258), .ZN(n1255) );
XOR2_X1 U942 ( .A(G116), .B(n1209), .Z(G18) );
AND3_X1 U943 ( .A1(n1073), .A2(n1075), .A3(n1254), .ZN(n1209) );
INV_X1 U944 ( .A(n1247), .ZN(n1075) );
NAND2_X1 U945 ( .A1(n1237), .A2(n1259), .ZN(n1247) );
XNOR2_X1 U946 ( .A(KEYINPUT59), .B(n1260), .ZN(n1259) );
NAND2_X1 U947 ( .A1(n1261), .A2(n1262), .ZN(G15) );
NAND2_X1 U948 ( .A1(G113), .A2(n1210), .ZN(n1262) );
XOR2_X1 U949 ( .A(KEYINPUT23), .B(n1263), .Z(n1261) );
NOR2_X1 U950 ( .A1(G113), .A2(n1210), .ZN(n1263) );
NAND3_X1 U951 ( .A1(n1073), .A2(n1076), .A3(n1254), .ZN(n1210) );
AND3_X1 U952 ( .A1(n1057), .A2(n1264), .A3(n1071), .ZN(n1254) );
NOR2_X1 U953 ( .A1(n1062), .A2(n1265), .ZN(n1071) );
XOR2_X1 U954 ( .A(KEYINPUT21), .B(n1266), .Z(n1265) );
NOR2_X1 U955 ( .A1(n1260), .A2(n1237), .ZN(n1076) );
INV_X1 U956 ( .A(n1236), .ZN(n1260) );
NOR2_X1 U957 ( .A1(n1256), .A2(n1258), .ZN(n1073) );
XNOR2_X1 U958 ( .A(G110), .B(n1267), .ZN(G12) );
NAND2_X1 U959 ( .A1(KEYINPUT22), .A2(n1207), .ZN(n1267) );
AND3_X1 U960 ( .A1(n1068), .A2(n1211), .A3(n1193), .ZN(n1207) );
NOR2_X1 U961 ( .A1(n1236), .A2(n1237), .ZN(n1193) );
XNOR2_X1 U962 ( .A(G478), .B(n1268), .ZN(n1237) );
NOR2_X1 U963 ( .A1(n1083), .A2(KEYINPUT48), .ZN(n1268) );
NOR2_X1 U964 ( .A1(n1143), .A2(G902), .ZN(n1083) );
XOR2_X1 U965 ( .A(n1269), .B(n1270), .Z(n1143) );
XOR2_X1 U966 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U967 ( .A(G128), .B(G122), .Z(n1272) );
XOR2_X1 U968 ( .A(KEYINPUT18), .B(G134), .Z(n1271) );
XOR2_X1 U969 ( .A(n1273), .B(n1274), .Z(n1269) );
XOR2_X1 U970 ( .A(G116), .B(G107), .Z(n1274) );
XOR2_X1 U971 ( .A(n1275), .B(n1276), .Z(n1273) );
NOR2_X1 U972 ( .A1(KEYINPUT4), .A2(n1277), .ZN(n1276) );
NAND2_X1 U973 ( .A1(n1278), .A2(G217), .ZN(n1275) );
XOR2_X1 U974 ( .A(n1086), .B(G475), .Z(n1236) );
NOR2_X1 U975 ( .A1(n1151), .A2(G902), .ZN(n1086) );
INV_X1 U976 ( .A(n1149), .ZN(n1151) );
XOR2_X1 U977 ( .A(n1279), .B(n1280), .Z(n1149) );
XOR2_X1 U978 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U979 ( .A(n1152), .B(n1283), .Z(n1282) );
NAND3_X1 U980 ( .A1(n1284), .A2(n1285), .A3(KEYINPUT42), .ZN(n1283) );
NAND2_X1 U981 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
INV_X1 U982 ( .A(KEYINPUT45), .ZN(n1287) );
XOR2_X1 U983 ( .A(G143), .B(n1288), .Z(n1286) );
NAND3_X1 U984 ( .A1(n1288), .A2(G143), .A3(KEYINPUT45), .ZN(n1284) );
AND3_X1 U985 ( .A1(G214), .A2(n1289), .A3(n1290), .ZN(n1288) );
XOR2_X1 U986 ( .A(n1095), .B(KEYINPUT39), .Z(n1290) );
INV_X1 U987 ( .A(G104), .ZN(n1152) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1279) );
XOR2_X1 U989 ( .A(G122), .B(G113), .Z(n1292) );
XOR2_X1 U990 ( .A(n1242), .B(G140), .Z(n1291) );
AND3_X1 U991 ( .A1(n1245), .A2(n1264), .A3(n1057), .ZN(n1211) );
INV_X1 U992 ( .A(n1198), .ZN(n1057) );
NAND2_X1 U993 ( .A1(n1059), .A2(n1058), .ZN(n1198) );
NAND3_X1 U994 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1058) );
INV_X1 U995 ( .A(n1088), .ZN(n1295) );
NOR2_X1 U996 ( .A1(n1090), .A2(n1296), .ZN(n1088) );
NAND3_X1 U997 ( .A1(KEYINPUT55), .A2(n1296), .A3(n1090), .ZN(n1294) );
INV_X1 U998 ( .A(n1091), .ZN(n1296) );
NAND2_X1 U999 ( .A1(G210), .A2(n1297), .ZN(n1091) );
OR2_X1 U1000 ( .A1(n1090), .A2(KEYINPUT55), .ZN(n1293) );
NAND2_X1 U1001 ( .A1(n1298), .A2(n1299), .ZN(n1090) );
XOR2_X1 U1002 ( .A(n1300), .B(n1301), .Z(n1298) );
XOR2_X1 U1003 ( .A(n1219), .B(n1164), .Z(n1301) );
NAND2_X1 U1004 ( .A1(n1302), .A2(n1303), .ZN(n1219) );
OR2_X1 U1005 ( .A1(n1304), .A2(n1126), .ZN(n1303) );
XOR2_X1 U1006 ( .A(n1305), .B(KEYINPUT40), .Z(n1302) );
NAND2_X1 U1007 ( .A1(n1126), .A2(n1304), .ZN(n1305) );
XNOR2_X1 U1008 ( .A(n1306), .B(n1130), .ZN(n1304) );
AND2_X1 U1009 ( .A1(n1307), .A2(n1308), .ZN(n1130) );
NAND2_X1 U1010 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U1011 ( .A(n1311), .B(G107), .Z(n1309) );
NAND2_X1 U1012 ( .A1(n1312), .A2(G101), .ZN(n1307) );
XOR2_X1 U1013 ( .A(n1313), .B(n1311), .Z(n1312) );
NAND2_X1 U1014 ( .A1(KEYINPUT6), .A2(G104), .ZN(n1311) );
INV_X1 U1015 ( .A(G107), .ZN(n1313) );
NAND2_X1 U1016 ( .A1(KEYINPUT1), .A2(n1314), .ZN(n1306) );
XOR2_X1 U1017 ( .A(KEYINPUT58), .B(n1131), .Z(n1314) );
XNOR2_X1 U1018 ( .A(n1315), .B(n1316), .ZN(n1131) );
NOR2_X1 U1019 ( .A1(KEYINPUT16), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1020 ( .A(G110), .B(n1318), .ZN(n1126) );
NOR2_X1 U1021 ( .A1(KEYINPUT31), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U1022 ( .A(G122), .B(KEYINPUT7), .ZN(n1319) );
XOR2_X1 U1023 ( .A(G125), .B(n1226), .Z(n1300) );
AND2_X1 U1024 ( .A1(G224), .A2(n1095), .ZN(n1226) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1297), .ZN(n1059) );
NAND2_X1 U1026 ( .A1(n1289), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1027 ( .A1(n1042), .A2(n1320), .ZN(n1264) );
NAND4_X1 U1028 ( .A1(n1128), .A2(G953), .A3(G902), .A4(n1253), .ZN(n1320) );
XNOR2_X1 U1029 ( .A(G898), .B(KEYINPUT27), .ZN(n1128) );
NAND3_X1 U1030 ( .A1(n1253), .A2(n1095), .A3(G952), .ZN(n1042) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1253) );
XOR2_X1 U1032 ( .A(n1065), .B(KEYINPUT2), .Z(n1245) );
NAND2_X1 U1033 ( .A1(n1321), .A2(n1062), .ZN(n1065) );
XNOR2_X1 U1034 ( .A(n1322), .B(G469), .ZN(n1062) );
NAND2_X1 U1035 ( .A1(n1323), .A2(n1299), .ZN(n1322) );
XOR2_X1 U1036 ( .A(n1166), .B(n1113), .Z(n1323) );
XOR2_X1 U1037 ( .A(n1324), .B(n1325), .Z(n1113) );
XOR2_X1 U1038 ( .A(G146), .B(G128), .Z(n1325) );
NAND2_X1 U1039 ( .A1(KEYINPUT46), .A2(G143), .ZN(n1324) );
XOR2_X1 U1040 ( .A(n1326), .B(n1327), .Z(n1166) );
XOR2_X1 U1041 ( .A(G104), .B(n1328), .Z(n1327) );
XOR2_X1 U1042 ( .A(G110), .B(G107), .Z(n1328) );
XOR2_X1 U1043 ( .A(n1329), .B(n1330), .Z(n1326) );
INV_X1 U1044 ( .A(n1109), .ZN(n1330) );
XNOR2_X1 U1045 ( .A(n1331), .B(n1332), .ZN(n1109) );
XOR2_X1 U1046 ( .A(n1310), .B(n1333), .Z(n1329) );
NOR2_X1 U1047 ( .A1(G953), .A2(n1096), .ZN(n1333) );
INV_X1 U1048 ( .A(G227), .ZN(n1096) );
XOR2_X1 U1049 ( .A(KEYINPUT21), .B(n1063), .Z(n1321) );
INV_X1 U1050 ( .A(n1266), .ZN(n1063) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1334), .ZN(n1266) );
AND2_X1 U1052 ( .A1(n1335), .A2(n1256), .ZN(n1068) );
XOR2_X1 U1053 ( .A(n1336), .B(n1136), .Z(n1256) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1334), .ZN(n1136) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1337), .ZN(n1334) );
XOR2_X1 U1056 ( .A(KEYINPUT38), .B(G902), .Z(n1337) );
NAND2_X1 U1057 ( .A1(n1134), .A2(n1299), .ZN(n1336) );
XNOR2_X1 U1058 ( .A(n1338), .B(n1339), .ZN(n1134) );
XNOR2_X1 U1059 ( .A(n1332), .B(n1340), .ZN(n1339) );
XOR2_X1 U1060 ( .A(n1341), .B(n1281), .Z(n1340) );
XOR2_X1 U1061 ( .A(G125), .B(G146), .Z(n1281) );
NAND2_X1 U1062 ( .A1(n1278), .A2(G221), .ZN(n1341) );
AND2_X1 U1063 ( .A1(G234), .A2(n1095), .ZN(n1278) );
XOR2_X1 U1064 ( .A(G137), .B(G140), .Z(n1332) );
XOR2_X1 U1065 ( .A(n1342), .B(n1343), .Z(n1338) );
NOR2_X1 U1066 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1067 ( .A(n1346), .B(KEYINPUT44), .Z(n1345) );
NAND2_X1 U1068 ( .A1(G110), .A2(n1347), .ZN(n1346) );
NOR2_X1 U1069 ( .A1(G110), .A2(n1347), .ZN(n1344) );
XOR2_X1 U1070 ( .A(G128), .B(G119), .Z(n1347) );
XNOR2_X1 U1071 ( .A(KEYINPUT26), .B(KEYINPUT19), .ZN(n1342) );
XOR2_X1 U1072 ( .A(n1258), .B(KEYINPUT28), .Z(n1335) );
XOR2_X1 U1073 ( .A(n1348), .B(G472), .Z(n1258) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1299), .ZN(n1348) );
INV_X1 U1075 ( .A(G902), .ZN(n1299) );
XOR2_X1 U1076 ( .A(n1161), .B(n1350), .Z(n1349) );
XNOR2_X1 U1077 ( .A(n1351), .B(n1156), .ZN(n1350) );
XNOR2_X1 U1078 ( .A(n1310), .B(n1352), .ZN(n1156) );
AND3_X1 U1079 ( .A1(G210), .A2(n1095), .A3(n1289), .ZN(n1352) );
INV_X1 U1080 ( .A(G237), .ZN(n1289) );
INV_X1 U1081 ( .A(G953), .ZN(n1095) );
INV_X1 U1082 ( .A(G101), .ZN(n1310) );
NAND2_X1 U1083 ( .A1(n1353), .A2(KEYINPUT25), .ZN(n1351) );
XOR2_X1 U1084 ( .A(n1163), .B(n1354), .Z(n1353) );
NOR2_X1 U1085 ( .A1(KEYINPUT47), .A2(n1164), .ZN(n1354) );
XOR2_X1 U1086 ( .A(n1355), .B(G128), .Z(n1164) );
NAND2_X1 U1087 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1088 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1089 ( .A(KEYINPUT36), .B(G143), .Z(n1359) );
XOR2_X1 U1090 ( .A(KEYINPUT29), .B(n1230), .Z(n1358) );
INV_X1 U1091 ( .A(G146), .ZN(n1230) );
XOR2_X1 U1092 ( .A(n1360), .B(KEYINPUT17), .Z(n1356) );
NAND2_X1 U1093 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1094 ( .A(KEYINPUT29), .B(G146), .Z(n1362) );
XOR2_X1 U1095 ( .A(KEYINPUT36), .B(n1277), .Z(n1361) );
INV_X1 U1096 ( .A(G143), .ZN(n1277) );
XNOR2_X1 U1097 ( .A(G137), .B(n1331), .ZN(n1163) );
XNOR2_X1 U1098 ( .A(n1242), .B(G134), .ZN(n1331) );
INV_X1 U1099 ( .A(G131), .ZN(n1242) );
XNOR2_X1 U1100 ( .A(n1315), .B(n1363), .ZN(n1161) );
XOR2_X1 U1101 ( .A(KEYINPUT41), .B(n1317), .Z(n1363) );
XOR2_X1 U1102 ( .A(G116), .B(KEYINPUT15), .Z(n1317) );
XNOR2_X1 U1103 ( .A(G113), .B(G119), .ZN(n1315) );
endmodule


