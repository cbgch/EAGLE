//Key = 0111111101011000001010011111011011011100011010100010001110010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;

XOR2_X1 U713 ( .A(n993), .B(n994), .Z(G9) );
NOR2_X1 U714 ( .A1(KEYINPUT16), .A2(n995), .ZN(n994) );
NOR2_X1 U715 ( .A1(n996), .A2(n997), .ZN(G75) );
NOR4_X1 U716 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n997) );
XOR2_X1 U717 ( .A(KEYINPUT61), .B(n1002), .Z(n999) );
AND4_X1 U718 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NAND4_X1 U719 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n998) );
NAND4_X1 U720 ( .A1(n1011), .A2(n1004), .A3(n1012), .A4(n1013), .ZN(n1008) );
NAND3_X1 U721 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND2_X1 U722 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U723 ( .A1(n1019), .A2(n1020), .ZN(n1015) );
NAND2_X1 U724 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U725 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U726 ( .A1(n1025), .A2(n1026), .ZN(n1014) );
XOR2_X1 U727 ( .A(KEYINPUT14), .B(n1018), .Z(n1026) );
NAND2_X1 U728 ( .A1(n1005), .A2(n1027), .ZN(n1007) );
NAND2_X1 U729 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U730 ( .A1(n1012), .A2(n1030), .ZN(n1029) );
OR2_X1 U731 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U732 ( .A1(n1004), .A2(n1033), .ZN(n1028) );
AND3_X1 U733 ( .A1(n1018), .A2(n1019), .A3(n1011), .ZN(n1005) );
INV_X1 U734 ( .A(n1034), .ZN(n1011) );
NOR3_X1 U735 ( .A1(n1035), .A2(G953), .A3(n1036), .ZN(n996) );
INV_X1 U736 ( .A(n1009), .ZN(n1036) );
NAND4_X1 U737 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1009) );
NOR4_X1 U738 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
XNOR2_X1 U739 ( .A(n1045), .B(n1046), .ZN(n1044) );
XNOR2_X1 U740 ( .A(G478), .B(KEYINPUT57), .ZN(n1046) );
XNOR2_X1 U741 ( .A(n1047), .B(KEYINPUT55), .ZN(n1042) );
XNOR2_X1 U742 ( .A(n1048), .B(KEYINPUT18), .ZN(n1041) );
NOR3_X1 U743 ( .A1(n1049), .A2(n1006), .A3(n1023), .ZN(n1039) );
NOR2_X1 U744 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
INV_X1 U745 ( .A(n1052), .ZN(n1050) );
XOR2_X1 U746 ( .A(KEYINPUT41), .B(n1053), .Z(n1038) );
NOR2_X1 U747 ( .A1(n1054), .A2(n1052), .ZN(n1053) );
XOR2_X1 U748 ( .A(n1051), .B(KEYINPUT11), .Z(n1054) );
XNOR2_X1 U749 ( .A(G469), .B(n1055), .ZN(n1037) );
NAND2_X1 U750 ( .A1(KEYINPUT33), .A2(n1056), .ZN(n1055) );
XNOR2_X1 U751 ( .A(KEYINPUT4), .B(n1057), .ZN(n1056) );
XNOR2_X1 U752 ( .A(KEYINPUT22), .B(n1000), .ZN(n1035) );
INV_X1 U753 ( .A(G952), .ZN(n1000) );
XOR2_X1 U754 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U755 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1010), .ZN(n1061) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1060) );
NAND2_X1 U759 ( .A1(G953), .A2(n1064), .ZN(n1066) );
INV_X1 U760 ( .A(G900), .ZN(n1064) );
XOR2_X1 U761 ( .A(n1067), .B(n1068), .Z(n1065) );
XOR2_X1 U762 ( .A(n1069), .B(n1070), .Z(n1067) );
NAND2_X1 U763 ( .A1(KEYINPUT42), .A2(n1071), .ZN(n1069) );
NAND2_X1 U764 ( .A1(n1010), .A2(n1072), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(G69) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
INV_X1 U768 ( .A(n1075), .ZN(n1078) );
NOR2_X1 U769 ( .A1(KEYINPUT51), .A2(n1079), .ZN(n1075) );
XOR2_X1 U770 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U772 ( .A(KEYINPUT62), .B(n1084), .Z(n1083) );
NAND2_X1 U773 ( .A1(n1010), .A2(n1085), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U775 ( .A1(n1088), .A2(n1076), .ZN(n1077) );
NAND2_X1 U776 ( .A1(G953), .A2(n1089), .ZN(n1076) );
INV_X1 U777 ( .A(n1082), .ZN(n1088) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(G66) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U781 ( .A1(n1090), .A2(n1096), .ZN(G63) );
NOR3_X1 U782 ( .A1(n1045), .A2(n1097), .A3(n1098), .ZN(n1096) );
NOR3_X1 U783 ( .A1(n1099), .A2(n1100), .A3(n1095), .ZN(n1098) );
INV_X1 U784 ( .A(G478), .ZN(n1100) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
AND2_X1 U786 ( .A1(n1001), .A2(G478), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1090), .A2(n1103), .ZN(G60) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND3_X1 U789 ( .A1(n1106), .A2(n1001), .A3(G475), .ZN(n1104) );
XNOR2_X1 U790 ( .A(KEYINPUT52), .B(n1107), .ZN(n1106) );
XOR2_X1 U791 ( .A(n1108), .B(n1109), .Z(G6) );
XNOR2_X1 U792 ( .A(G104), .B(KEYINPUT3), .ZN(n1108) );
NOR2_X1 U793 ( .A1(n1090), .A2(n1110), .ZN(G57) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1112) );
XNOR2_X1 U796 ( .A(n1115), .B(n1116), .ZN(n1114) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U798 ( .A1(KEYINPUT35), .A2(n1119), .ZN(n1113) );
AND2_X1 U799 ( .A1(n1118), .A2(n1117), .ZN(n1111) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1117) );
XOR2_X1 U801 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U802 ( .A1(n1124), .A2(n1095), .ZN(n1123) );
INV_X1 U803 ( .A(G472), .ZN(n1124) );
NOR3_X1 U804 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
NOR2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
INV_X1 U807 ( .A(KEYINPUT36), .ZN(n1131) );
XOR2_X1 U808 ( .A(n1132), .B(KEYINPUT12), .Z(n1130) );
AND3_X1 U809 ( .A1(n1129), .A2(n1132), .A3(KEYINPUT36), .ZN(n1126) );
XNOR2_X1 U810 ( .A(n1133), .B(n1134), .ZN(n1129) );
NOR2_X1 U811 ( .A1(KEYINPUT36), .A2(n1132), .ZN(n1125) );
XOR2_X1 U812 ( .A(n1135), .B(KEYINPUT38), .Z(n1132) );
INV_X1 U813 ( .A(KEYINPUT7), .ZN(n1118) );
NOR2_X1 U814 ( .A1(n1090), .A2(n1136), .ZN(G54) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1137) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1095), .ZN(n1142) );
XNOR2_X1 U819 ( .A(n1144), .B(n1145), .ZN(n1141) );
NOR2_X1 U820 ( .A1(G140), .A2(KEYINPUT47), .ZN(n1145) );
NOR2_X1 U821 ( .A1(KEYINPUT17), .A2(n1146), .ZN(n1144) );
XOR2_X1 U822 ( .A(KEYINPUT26), .B(n1147), .Z(n1146) );
NOR2_X1 U823 ( .A1(n1090), .A2(n1148), .ZN(G51) );
XOR2_X1 U824 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1149) );
NOR2_X1 U826 ( .A1(n1052), .A2(n1095), .ZN(n1152) );
NAND2_X1 U827 ( .A1(G902), .A2(n1001), .ZN(n1095) );
NAND3_X1 U828 ( .A1(n1153), .A2(n1086), .A3(n1154), .ZN(n1001) );
XOR2_X1 U829 ( .A(n1087), .B(KEYINPUT21), .Z(n1154) );
AND4_X1 U830 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1086) );
NOR4_X1 U831 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n993), .ZN(n1158) );
AND2_X1 U832 ( .A1(n1032), .A2(n1162), .ZN(n993) );
NOR2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1157) );
NOR3_X1 U834 ( .A1(n1165), .A2(n1021), .A3(n1166), .ZN(n1164) );
NAND3_X1 U835 ( .A1(n1162), .A2(n1167), .A3(n1168), .ZN(n1156) );
INV_X1 U836 ( .A(KEYINPUT2), .ZN(n1168) );
NAND2_X1 U837 ( .A1(n1109), .A2(KEYINPUT2), .ZN(n1155) );
AND2_X1 U838 ( .A1(n1031), .A2(n1162), .ZN(n1109) );
AND4_X1 U839 ( .A1(n1169), .A2(n1033), .A3(n1019), .A4(n1170), .ZN(n1162) );
INV_X1 U840 ( .A(n1072), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1171), .A2(n1172), .ZN(n1072) );
NOR4_X1 U842 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
NOR4_X1 U843 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U845 ( .A(n1025), .B(KEYINPUT39), .ZN(n1181) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1184), .ZN(n1179) );
XNOR2_X1 U847 ( .A(n1185), .B(KEYINPUT37), .ZN(n1183) );
INV_X1 U848 ( .A(n1186), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1010), .A2(G952), .ZN(n1090) );
XOR2_X1 U850 ( .A(G146), .B(n1178), .Z(G48) );
AND3_X1 U851 ( .A1(n1031), .A2(n1169), .A3(n1187), .ZN(n1178) );
XNOR2_X1 U852 ( .A(G143), .B(n1186), .ZN(G45) );
NAND4_X1 U853 ( .A1(n1169), .A2(n1033), .A3(n1017), .A4(n1188), .ZN(n1186) );
NOR3_X1 U854 ( .A1(n1189), .A2(n1185), .A3(n1190), .ZN(n1188) );
XOR2_X1 U855 ( .A(G140), .B(n1191), .Z(G42) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1182), .ZN(n1191) );
XOR2_X1 U857 ( .A(n1176), .B(n1193), .Z(G39) );
NOR2_X1 U858 ( .A1(KEYINPUT40), .A2(n1194), .ZN(n1193) );
AND3_X1 U859 ( .A1(n1018), .A2(n1187), .A3(n1004), .ZN(n1176) );
XNOR2_X1 U860 ( .A(n1071), .B(n1195), .ZN(G36) );
NOR3_X1 U861 ( .A1(n1184), .A2(KEYINPUT43), .A3(n1185), .ZN(n1195) );
INV_X1 U862 ( .A(n1196), .ZN(n1185) );
NAND4_X1 U863 ( .A1(n1017), .A2(n1018), .A3(n1032), .A4(n1033), .ZN(n1184) );
XOR2_X1 U864 ( .A(n1175), .B(n1197), .Z(G33) );
XOR2_X1 U865 ( .A(KEYINPUT60), .B(G131), .Z(n1197) );
NOR2_X1 U866 ( .A1(n1166), .A2(n1182), .ZN(n1175) );
NAND4_X1 U867 ( .A1(n1018), .A2(n1031), .A3(n1033), .A4(n1196), .ZN(n1182) );
NOR2_X1 U868 ( .A1(n1198), .A2(n1023), .ZN(n1018) );
XNOR2_X1 U869 ( .A(G128), .B(n1199), .ZN(G30) );
NOR2_X1 U870 ( .A1(n1174), .A2(KEYINPUT48), .ZN(n1199) );
AND3_X1 U871 ( .A1(n1032), .A2(n1169), .A3(n1187), .ZN(n1174) );
AND4_X1 U872 ( .A1(n1033), .A2(n1047), .A3(n1043), .A4(n1196), .ZN(n1187) );
XOR2_X1 U873 ( .A(G101), .B(n1200), .Z(G3) );
NOR3_X1 U874 ( .A1(n1201), .A2(n1166), .A3(n1165), .ZN(n1200) );
XNOR2_X1 U875 ( .A(KEYINPUT50), .B(n1021), .ZN(n1201) );
XNOR2_X1 U876 ( .A(n1173), .B(n1202), .ZN(G27) );
NOR2_X1 U877 ( .A1(G125), .A2(KEYINPUT49), .ZN(n1202) );
AND4_X1 U878 ( .A1(n1169), .A2(n1196), .A3(n1012), .A4(n1203), .ZN(n1173) );
NOR2_X1 U879 ( .A1(n1167), .A2(n1192), .ZN(n1203) );
INV_X1 U880 ( .A(n1031), .ZN(n1167) );
NAND2_X1 U881 ( .A1(n1034), .A2(n1204), .ZN(n1196) );
NAND4_X1 U882 ( .A1(n1205), .A2(G902), .A3(G953), .A4(n1206), .ZN(n1204) );
XNOR2_X1 U883 ( .A(G900), .B(KEYINPUT15), .ZN(n1205) );
XOR2_X1 U884 ( .A(G122), .B(n1163), .Z(G24) );
AND4_X1 U885 ( .A1(n1207), .A2(n1019), .A3(n1208), .A4(n1048), .ZN(n1163) );
NOR2_X1 U886 ( .A1(n1043), .A2(n1047), .ZN(n1019) );
XOR2_X1 U887 ( .A(G119), .B(n1161), .Z(G21) );
AND4_X1 U888 ( .A1(n1207), .A2(n1004), .A3(n1047), .A4(n1043), .ZN(n1161) );
XOR2_X1 U889 ( .A(G116), .B(n1160), .Z(G18) );
AND3_X1 U890 ( .A1(n1017), .A2(n1032), .A3(n1207), .ZN(n1160) );
NOR2_X1 U891 ( .A1(n1048), .A2(n1189), .ZN(n1032) );
INV_X1 U892 ( .A(n1208), .ZN(n1189) );
XOR2_X1 U893 ( .A(G113), .B(n1209), .Z(G15) );
NOR2_X1 U894 ( .A1(KEYINPUT28), .A2(n1087), .ZN(n1209) );
NAND3_X1 U895 ( .A1(n1017), .A2(n1031), .A3(n1207), .ZN(n1087) );
AND3_X1 U896 ( .A1(n1169), .A2(n1170), .A3(n1012), .ZN(n1207) );
NOR2_X1 U897 ( .A1(n1210), .A2(n1006), .ZN(n1012) );
INV_X1 U898 ( .A(n1003), .ZN(n1210) );
NOR2_X1 U899 ( .A1(n1208), .A2(n1190), .ZN(n1031) );
INV_X1 U900 ( .A(n1048), .ZN(n1190) );
INV_X1 U901 ( .A(n1166), .ZN(n1017) );
NAND2_X1 U902 ( .A1(n1211), .A2(n1047), .ZN(n1166) );
XNOR2_X1 U903 ( .A(n1212), .B(n1159), .ZN(G12) );
NOR3_X1 U904 ( .A1(n1192), .A2(n1021), .A3(n1165), .ZN(n1159) );
NAND3_X1 U905 ( .A1(n1033), .A2(n1170), .A3(n1004), .ZN(n1165) );
NOR2_X1 U906 ( .A1(n1048), .A2(n1208), .ZN(n1004) );
XOR2_X1 U907 ( .A(G478), .B(n1213), .Z(n1208) );
NOR2_X1 U908 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U909 ( .A1(KEYINPUT58), .A2(n1045), .ZN(n1215) );
AND2_X1 U910 ( .A1(KEYINPUT45), .A2(n1045), .ZN(n1214) );
NOR2_X1 U911 ( .A1(n1101), .A2(G902), .ZN(n1045) );
INV_X1 U912 ( .A(n1099), .ZN(n1101) );
NAND2_X1 U913 ( .A1(n1216), .A2(n1217), .ZN(n1099) );
NAND2_X1 U914 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U915 ( .A(KEYINPUT59), .B(n1220), .Z(n1216) );
NOR2_X1 U916 ( .A1(n1218), .A2(n1219), .ZN(n1220) );
XNOR2_X1 U917 ( .A(n1221), .B(n1222), .ZN(n1219) );
XNOR2_X1 U918 ( .A(G116), .B(n995), .ZN(n1222) );
XOR2_X1 U919 ( .A(n1223), .B(n1224), .Z(n1221) );
NAND2_X1 U920 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NAND2_X1 U921 ( .A1(G134), .A2(n1227), .ZN(n1226) );
XOR2_X1 U922 ( .A(KEYINPUT63), .B(n1228), .Z(n1225) );
NOR2_X1 U923 ( .A1(G134), .A2(n1227), .ZN(n1228) );
XNOR2_X1 U924 ( .A(n1229), .B(G128), .ZN(n1227) );
INV_X1 U925 ( .A(G143), .ZN(n1229) );
NOR3_X1 U926 ( .A1(n1094), .A2(G953), .A3(n1230), .ZN(n1218) );
XNOR2_X1 U927 ( .A(n1231), .B(G475), .ZN(n1048) );
NAND2_X1 U928 ( .A1(n1105), .A2(n1107), .ZN(n1231) );
XNOR2_X1 U929 ( .A(n1232), .B(n1233), .ZN(n1105) );
XOR2_X1 U930 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U931 ( .A(G146), .B(G131), .Z(n1235) );
NOR2_X1 U932 ( .A1(KEYINPUT10), .A2(n1236), .ZN(n1234) );
XOR2_X1 U933 ( .A(n1237), .B(G125), .Z(n1236) );
NAND2_X1 U934 ( .A1(KEYINPUT54), .A2(G140), .ZN(n1237) );
XNOR2_X1 U935 ( .A(n1238), .B(n1239), .ZN(n1232) );
XOR2_X1 U936 ( .A(n1240), .B(n1241), .Z(n1239) );
NAND2_X1 U937 ( .A1(KEYINPUT1), .A2(n1242), .ZN(n1241) );
INV_X1 U938 ( .A(G104), .ZN(n1242) );
NAND2_X1 U939 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
NAND4_X1 U940 ( .A1(G214), .A2(n1245), .A3(n1246), .A4(n1010), .ZN(n1244) );
XOR2_X1 U941 ( .A(n1247), .B(KEYINPUT53), .Z(n1243) );
NAND2_X1 U942 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND3_X1 U943 ( .A1(n1246), .A2(n1010), .A3(G214), .ZN(n1249) );
INV_X1 U944 ( .A(n1245), .ZN(n1248) );
XOR2_X1 U945 ( .A(G143), .B(KEYINPUT19), .Z(n1245) );
NAND2_X1 U946 ( .A1(n1034), .A2(n1250), .ZN(n1170) );
NAND3_X1 U947 ( .A1(n1082), .A2(n1206), .A3(G902), .ZN(n1250) );
NOR2_X1 U948 ( .A1(G898), .A2(n1010), .ZN(n1082) );
NAND3_X1 U949 ( .A1(n1206), .A2(n1010), .A3(G952), .ZN(n1034) );
NAND2_X1 U950 ( .A1(G237), .A2(G234), .ZN(n1206) );
NOR2_X1 U951 ( .A1(n1003), .A2(n1006), .ZN(n1033) );
NOR2_X1 U952 ( .A1(n1251), .A2(n1252), .ZN(n1006) );
NAND3_X1 U953 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1003) );
NAND2_X1 U954 ( .A1(KEYINPUT13), .A2(G469), .ZN(n1255) );
NAND3_X1 U955 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1254) );
INV_X1 U956 ( .A(KEYINPUT13), .ZN(n1257) );
OR2_X1 U957 ( .A1(n1258), .A2(n1256), .ZN(n1253) );
AND2_X1 U958 ( .A1(KEYINPUT20), .A2(n1143), .ZN(n1256) );
INV_X1 U959 ( .A(G469), .ZN(n1143) );
XNOR2_X1 U960 ( .A(n1057), .B(KEYINPUT56), .ZN(n1258) );
NAND2_X1 U961 ( .A1(n1259), .A2(n1107), .ZN(n1057) );
XNOR2_X1 U962 ( .A(n1140), .B(n1260), .ZN(n1259) );
XOR2_X1 U963 ( .A(n1261), .B(G140), .Z(n1260) );
NAND2_X1 U964 ( .A1(KEYINPUT5), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U965 ( .A(n1147), .B(n1139), .ZN(n1262) );
XOR2_X1 U966 ( .A(n1263), .B(KEYINPUT30), .Z(n1139) );
XNOR2_X1 U967 ( .A(n1264), .B(n995), .ZN(n1147) );
XOR2_X1 U968 ( .A(G110), .B(n1265), .Z(n1140) );
NOR2_X1 U969 ( .A1(G953), .A2(n1063), .ZN(n1265) );
INV_X1 U970 ( .A(G227), .ZN(n1063) );
INV_X1 U971 ( .A(n1169), .ZN(n1021) );
NOR2_X1 U972 ( .A1(n1024), .A2(n1023), .ZN(n1169) );
AND2_X1 U973 ( .A1(G214), .A2(n1266), .ZN(n1023) );
INV_X1 U974 ( .A(n1198), .ZN(n1024) );
XOR2_X1 U975 ( .A(n1051), .B(n1052), .Z(n1198) );
NAND2_X1 U976 ( .A1(G210), .A2(n1266), .ZN(n1052) );
NAND2_X1 U977 ( .A1(n1246), .A2(n1107), .ZN(n1266) );
NAND2_X1 U978 ( .A1(n1267), .A2(n1107), .ZN(n1051) );
XOR2_X1 U979 ( .A(n1151), .B(n1268), .Z(n1267) );
XNOR2_X1 U980 ( .A(n1269), .B(KEYINPUT9), .ZN(n1268) );
NAND2_X1 U981 ( .A1(KEYINPUT24), .A2(n1150), .ZN(n1269) );
XOR2_X1 U982 ( .A(n1084), .B(KEYINPUT0), .Z(n1150) );
XNOR2_X1 U983 ( .A(n1270), .B(n1271), .ZN(n1084) );
XOR2_X1 U984 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U985 ( .A(KEYINPUT27), .B(G116), .Z(n1273) );
XOR2_X1 U986 ( .A(n1274), .B(n1238), .Z(n1270) );
XOR2_X1 U987 ( .A(G113), .B(n1224), .Z(n1238) );
XOR2_X1 U988 ( .A(G122), .B(KEYINPUT32), .Z(n1224) );
NAND2_X1 U989 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U990 ( .A1(n1277), .A2(G107), .ZN(n1276) );
NAND2_X1 U991 ( .A1(n1278), .A2(n995), .ZN(n1275) );
INV_X1 U992 ( .A(G107), .ZN(n995) );
XNOR2_X1 U993 ( .A(KEYINPUT8), .B(n1277), .ZN(n1278) );
INV_X1 U994 ( .A(n1264), .ZN(n1277) );
XOR2_X1 U995 ( .A(G104), .B(n1119), .Z(n1264) );
XOR2_X1 U996 ( .A(n1135), .B(n1279), .Z(n1151) );
XOR2_X1 U997 ( .A(G125), .B(n1280), .Z(n1279) );
NOR2_X1 U998 ( .A1(G953), .A2(n1089), .ZN(n1280) );
INV_X1 U999 ( .A(G224), .ZN(n1089) );
INV_X1 U1000 ( .A(n1025), .ZN(n1192) );
NOR2_X1 U1001 ( .A1(n1047), .A2(n1211), .ZN(n1025) );
INV_X1 U1002 ( .A(n1043), .ZN(n1211) );
XNOR2_X1 U1003 ( .A(n1281), .B(n1282), .ZN(n1043) );
NOR2_X1 U1004 ( .A1(n1252), .A2(n1094), .ZN(n1282) );
INV_X1 U1005 ( .A(G217), .ZN(n1094) );
AND2_X1 U1006 ( .A1(n1283), .A2(n1107), .ZN(n1252) );
XNOR2_X1 U1007 ( .A(KEYINPUT31), .B(n1230), .ZN(n1283) );
NAND2_X1 U1008 ( .A1(n1284), .A2(n1107), .ZN(n1281) );
INV_X1 U1009 ( .A(G902), .ZN(n1107) );
XNOR2_X1 U1010 ( .A(n1093), .B(KEYINPUT34), .ZN(n1284) );
XNOR2_X1 U1011 ( .A(n1285), .B(n1286), .ZN(n1093) );
XOR2_X1 U1012 ( .A(n1272), .B(n1068), .Z(n1286) );
XOR2_X1 U1013 ( .A(G125), .B(G140), .Z(n1068) );
XNOR2_X1 U1014 ( .A(n1212), .B(G119), .ZN(n1272) );
XNOR2_X1 U1015 ( .A(n1287), .B(n1288), .ZN(n1285) );
XOR2_X1 U1016 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR3_X1 U1017 ( .A1(n1251), .A2(G953), .A3(n1230), .ZN(n1289) );
INV_X1 U1018 ( .A(G234), .ZN(n1230) );
INV_X1 U1019 ( .A(G221), .ZN(n1251) );
XOR2_X1 U1020 ( .A(G472), .B(n1291), .Z(n1047) );
NOR2_X1 U1021 ( .A1(n1292), .A2(G902), .ZN(n1291) );
NOR2_X1 U1022 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U1023 ( .A(n1295), .B(KEYINPUT44), .Z(n1294) );
NAND2_X1 U1024 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XNOR2_X1 U1025 ( .A(n1298), .B(KEYINPUT6), .ZN(n1296) );
NOR2_X1 U1026 ( .A1(n1297), .A2(n1298), .ZN(n1293) );
XNOR2_X1 U1027 ( .A(n1115), .B(n1119), .ZN(n1298) );
XOR2_X1 U1028 ( .A(G101), .B(KEYINPUT25), .Z(n1119) );
NAND3_X1 U1029 ( .A1(n1246), .A2(n1010), .A3(G210), .ZN(n1115) );
INV_X1 U1030 ( .A(G953), .ZN(n1010) );
INV_X1 U1031 ( .A(G237), .ZN(n1246) );
XNOR2_X1 U1032 ( .A(n1263), .B(n1299), .ZN(n1297) );
INV_X1 U1033 ( .A(n1120), .ZN(n1299) );
XNOR2_X1 U1034 ( .A(n1300), .B(G113), .ZN(n1120) );
NAND2_X1 U1035 ( .A1(n1301), .A2(KEYINPUT46), .ZN(n1300) );
XNOR2_X1 U1036 ( .A(G119), .B(G116), .ZN(n1301) );
XNOR2_X1 U1037 ( .A(n1070), .B(n1134), .ZN(n1263) );
XNOR2_X1 U1038 ( .A(n1071), .B(KEYINPUT29), .ZN(n1134) );
INV_X1 U1039 ( .A(G134), .ZN(n1071) );
XOR2_X1 U1040 ( .A(n1135), .B(n1302), .Z(n1070) );
INV_X1 U1041 ( .A(n1133), .ZN(n1302) );
XOR2_X1 U1042 ( .A(G131), .B(n1290), .Z(n1133) );
XNOR2_X1 U1043 ( .A(n1194), .B(KEYINPUT23), .ZN(n1290) );
INV_X1 U1044 ( .A(G137), .ZN(n1194) );
XNOR2_X1 U1045 ( .A(G143), .B(n1287), .ZN(n1135) );
XOR2_X1 U1046 ( .A(G146), .B(G128), .Z(n1287) );
INV_X1 U1047 ( .A(G110), .ZN(n1212) );
endmodule


