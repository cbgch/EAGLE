//Key = 1001011100110100001011010111000101111000101100001000010110001111


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
n2243, n2244, n2245, n2246, n2247, n2248, n2249;

OR2_X1 U1265 ( .A1(n2248), .A2(STATO_REG_0__SCAN_IN), .ZN(n1693) );
INV_X2 U1266 ( .A(n1693), .ZN(n1694) );
INV_X2 U1267 ( .A(U280), .ZN(n1843) );
NAND2_X1 U1268 ( .A1(n1695), .A2(n1696), .ZN(U344) );
NAND2_X1 U1269 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1697), .ZN(n1696) );
NAND2_X1 U1270 ( .A1(n1698), .A2(DATA_IN_7_), .ZN(n1695) );
NAND2_X1 U1271 ( .A1(n1699), .A2(n1700), .ZN(U343) );
NAND2_X1 U1272 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1697), .ZN(n1700) );
NAND2_X1 U1273 ( .A1(n1698), .A2(DATA_IN_6_), .ZN(n1699) );
NAND2_X1 U1274 ( .A1(n1701), .A2(n1702), .ZN(U342) );
NAND2_X1 U1275 ( .A1(n1698), .A2(DATA_IN_5_), .ZN(n1702) );
XOR2_X1 U1276 ( .A(KEYINPUT53), .B(n1703), .Z(n1701) );
NOR2_X1 U1277 ( .A1(n1698), .A2(n1704), .ZN(n1703) );
NAND2_X1 U1278 ( .A1(n1705), .A2(n1706), .ZN(U341) );
NAND2_X1 U1279 ( .A1(n1698), .A2(DATA_IN_4_), .ZN(n1706) );
XOR2_X1 U1280 ( .A(KEYINPUT13), .B(n1707), .Z(n1705) );
NOR2_X1 U1281 ( .A1(n1698), .A2(n1708), .ZN(n1707) );
NAND2_X1 U1282 ( .A1(n1709), .A2(n1710), .ZN(U340) );
NAND2_X1 U1283 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1697), .ZN(n1710) );
NAND2_X1 U1284 ( .A1(n1698), .A2(DATA_IN_3_), .ZN(n1709) );
NAND2_X1 U1285 ( .A1(n1711), .A2(n1712), .ZN(U339) );
NAND2_X1 U1286 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1697), .ZN(n1712) );
NAND2_X1 U1287 ( .A1(n1713), .A2(n1698), .ZN(n1711) );
XNOR2_X1 U1288 ( .A(KEYINPUT24), .B(n1714), .ZN(n1713) );
NAND2_X1 U1289 ( .A1(n1715), .A2(n1716), .ZN(U338) );
NAND2_X1 U1290 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1697), .ZN(n1716) );
NAND2_X1 U1291 ( .A1(n1698), .A2(DATA_IN_1_), .ZN(n1715) );
NAND2_X1 U1292 ( .A1(n1717), .A2(n1718), .ZN(U337) );
NAND2_X1 U1293 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1697), .ZN(n1718) );
NAND2_X1 U1294 ( .A1(n1698), .A2(DATA_IN_0_), .ZN(n1717) );
INV_X1 U1295 ( .A(n1697), .ZN(n1698) );
NAND2_X1 U1296 ( .A1(n1719), .A2(n1720), .ZN(n1697) );
OR2_X1 U1297 ( .A1(n1721), .A2(STATO_REG_0__SCAN_IN), .ZN(n1720) );
NAND2_X1 U1298 ( .A1(n1722), .A2(n1723), .ZN(U336) );
NAND2_X1 U1299 ( .A1(n1724), .A2(DATA_IN_7_), .ZN(n1723) );
NAND2_X1 U1300 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1725), .ZN(n1722) );
NAND2_X1 U1301 ( .A1(n1726), .A2(n1727), .ZN(U335) );
NAND2_X1 U1302 ( .A1(n1724), .A2(DATA_IN_6_), .ZN(n1727) );
NAND2_X1 U1303 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1725), .ZN(n1726) );
NAND2_X1 U1304 ( .A1(n1728), .A2(n1729), .ZN(U334) );
NAND2_X1 U1305 ( .A1(n1724), .A2(DATA_IN_5_), .ZN(n1729) );
NAND2_X1 U1306 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1725), .ZN(n1728) );
NAND2_X1 U1307 ( .A1(n1730), .A2(n1731), .ZN(U333) );
NAND2_X1 U1308 ( .A1(n1724), .A2(DATA_IN_4_), .ZN(n1731) );
NAND2_X1 U1309 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1725), .ZN(n1730) );
NAND2_X1 U1310 ( .A1(n1732), .A2(n1733), .ZN(U332) );
NAND2_X1 U1311 ( .A1(n1724), .A2(DATA_IN_3_), .ZN(n1733) );
NAND2_X1 U1312 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1725), .ZN(n1732) );
NAND2_X1 U1313 ( .A1(n1734), .A2(n1735), .ZN(U331) );
NAND2_X1 U1314 ( .A1(n1736), .A2(n1725), .ZN(n1735) );
XNOR2_X1 U1315 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT35), .ZN(n1736) );
NAND2_X1 U1316 ( .A1(n1724), .A2(DATA_IN_2_), .ZN(n1734) );
NAND2_X1 U1317 ( .A1(n1737), .A2(n1738), .ZN(U330) );
NAND2_X1 U1318 ( .A1(n1739), .A2(n1724), .ZN(n1738) );
XNOR2_X1 U1319 ( .A(DATA_IN_1_), .B(KEYINPUT26), .ZN(n1739) );
NAND2_X1 U1320 ( .A1(n1740), .A2(n1725), .ZN(n1737) );
XNOR2_X1 U1321 ( .A(n1741), .B(KEYINPUT51), .ZN(n1740) );
NAND2_X1 U1322 ( .A1(n1742), .A2(n1743), .ZN(U329) );
NAND2_X1 U1323 ( .A1(n1724), .A2(DATA_IN_0_), .ZN(n1743) );
AND2_X1 U1324 ( .A1(n1744), .A2(n1719), .ZN(n1724) );
NAND2_X1 U1325 ( .A1(n1745), .A2(n1746), .ZN(n1744) );
NAND2_X1 U1326 ( .A1(n1747), .A2(n1748), .ZN(n1746) );
XNOR2_X1 U1327 ( .A(KEYINPUT27), .B(n1749), .ZN(n1747) );
XOR2_X1 U1328 ( .A(n1750), .B(KEYINPUT19), .Z(n1742) );
NAND2_X1 U1329 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1725), .ZN(n1750) );
NAND2_X1 U1330 ( .A1(n1719), .A2(n1751), .ZN(n1725) );
NAND2_X1 U1331 ( .A1(n1752), .A2(n1745), .ZN(n1751) );
NAND2_X1 U1332 ( .A1(n1748), .A2(n1749), .ZN(n1752) );
NAND2_X1 U1333 ( .A1(n1753), .A2(n1754), .ZN(n1749) );
NAND2_X1 U1334 ( .A1(n1755), .A2(n1756), .ZN(n1754) );
XNOR2_X1 U1335 ( .A(KEYINPUT16), .B(n1757), .ZN(n1755) );
NAND3_X1 U1336 ( .A1(n1758), .A2(n1759), .A3(n1760), .ZN(n1753) );
NAND2_X1 U1337 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1757), .ZN(n1760) );
NAND3_X1 U1338 ( .A1(n1761), .A2(n1762), .A3(n1763), .ZN(n1759) );
NAND2_X1 U1339 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1764), .ZN(n1763) );
NAND3_X1 U1340 ( .A1(n1765), .A2(n1766), .A3(n1767), .ZN(n1762) );
XOR2_X1 U1341 ( .A(n1768), .B(KEYINPUT9), .Z(n1767) );
NAND2_X1 U1342 ( .A1(DATA_IN_5_), .A2(n1769), .ZN(n1768) );
NAND3_X1 U1343 ( .A1(n1770), .A2(n1771), .A3(n1772), .ZN(n1766) );
NAND2_X1 U1344 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1773), .ZN(n1772) );
NAND3_X1 U1345 ( .A1(n1774), .A2(n1775), .A3(n1776), .ZN(n1771) );
NAND2_X1 U1346 ( .A1(DATA_IN_3_), .A2(n1777), .ZN(n1776) );
NAND3_X1 U1347 ( .A1(n1778), .A2(n1779), .A3(n1780), .ZN(n1775) );
NAND2_X1 U1348 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1714), .ZN(n1780) );
NAND3_X1 U1349 ( .A1(n1781), .A2(n1782), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1779) );
INV_X1 U1350 ( .A(DATA_IN_0_), .ZN(n1782) );
NAND2_X1 U1351 ( .A1(DATA_IN_1_), .A2(n1741), .ZN(n1781) );
NAND2_X1 U1352 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1783), .ZN(n1778) );
NAND2_X1 U1353 ( .A1(DATA_IN_2_), .A2(n1784), .ZN(n1774) );
NAND2_X1 U1354 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1785), .ZN(n1770) );
NAND2_X1 U1355 ( .A1(DATA_IN_4_), .A2(n1786), .ZN(n1765) );
NAND2_X1 U1356 ( .A1(n1787), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1761) );
XNOR2_X1 U1357 ( .A(DATA_IN_5_), .B(KEYINPUT45), .ZN(n1787) );
NAND2_X1 U1358 ( .A1(DATA_IN_6_), .A2(n1788), .ZN(n1758) );
XNOR2_X1 U1359 ( .A(n1721), .B(KEYINPUT44), .ZN(n1748) );
NAND2_X1 U1360 ( .A1(n1789), .A2(n1790), .ZN(n1721) );
NAND3_X1 U1361 ( .A1(n1791), .A2(n1792), .A3(n1793), .ZN(n1790) );
NAND2_X1 U1362 ( .A1(DATA_IN_7_), .A2(n1794), .ZN(n1793) );
NAND3_X1 U1363 ( .A1(n1795), .A2(n1796), .A3(n1797), .ZN(n1792) );
OR2_X1 U1364 ( .A1(n1764), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1797) );
NAND3_X1 U1365 ( .A1(n1798), .A2(n1799), .A3(n1800), .ZN(n1796) );
NAND2_X1 U1366 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1801), .ZN(n1800) );
NAND3_X1 U1367 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(n1799) );
NAND2_X1 U1368 ( .A1(DATA_IN_4_), .A2(n1708), .ZN(n1804) );
NAND3_X1 U1369 ( .A1(n1805), .A2(n1806), .A3(n1807), .ZN(n1803) );
XOR2_X1 U1370 ( .A(n1808), .B(KEYINPUT58), .Z(n1807) );
NAND2_X1 U1371 ( .A1(n1809), .A2(RMAX_REG_2__SCAN_IN), .ZN(n1808) );
XNOR2_X1 U1372 ( .A(DATA_IN_2_), .B(KEYINPUT30), .ZN(n1809) );
NAND3_X1 U1373 ( .A1(n1810), .A2(n1811), .A3(n1812), .ZN(n1806) );
NAND2_X1 U1374 ( .A1(DATA_IN_2_), .A2(n1813), .ZN(n1812) );
NAND3_X1 U1375 ( .A1(n1814), .A2(n1815), .A3(DATA_IN_0_), .ZN(n1811) );
INV_X1 U1376 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1815) );
NAND2_X1 U1377 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1783), .ZN(n1814) );
NAND2_X1 U1378 ( .A1(DATA_IN_1_), .A2(n1816), .ZN(n1810) );
NAND2_X1 U1379 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1785), .ZN(n1805) );
NAND2_X1 U1380 ( .A1(n1817), .A2(n1818), .ZN(n1802) );
XNOR2_X1 U1381 ( .A(DATA_IN_3_), .B(KEYINPUT55), .ZN(n1817) );
NAND2_X1 U1382 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1773), .ZN(n1798) );
NAND2_X1 U1383 ( .A1(DATA_IN_5_), .A2(n1704), .ZN(n1795) );
NAND2_X1 U1384 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1764), .ZN(n1791) );
XOR2_X1 U1385 ( .A(KEYINPUT42), .B(n1819), .Z(n1789) );
NOR2_X1 U1386 ( .A1(DATA_IN_7_), .A2(n1794), .ZN(n1819) );
NAND2_X1 U1387 ( .A1(n1820), .A2(n1821), .ZN(U328) );
NAND2_X1 U1388 ( .A1(n1822), .A2(DATA_IN_7_), .ZN(n1821) );
NAND2_X1 U1389 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1823), .ZN(n1820) );
NAND2_X1 U1390 ( .A1(n1824), .A2(n1825), .ZN(U327) );
NAND2_X1 U1391 ( .A1(n1822), .A2(DATA_IN_6_), .ZN(n1825) );
NAND2_X1 U1392 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1823), .ZN(n1824) );
NAND2_X1 U1393 ( .A1(n1826), .A2(n1827), .ZN(U326) );
NAND2_X1 U1394 ( .A1(n1822), .A2(DATA_IN_5_), .ZN(n1827) );
NAND2_X1 U1395 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1823), .ZN(n1826) );
NAND2_X1 U1396 ( .A1(n1828), .A2(n1829), .ZN(U325) );
NAND2_X1 U1397 ( .A1(n1822), .A2(DATA_IN_4_), .ZN(n1829) );
NAND2_X1 U1398 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1823), .ZN(n1828) );
NAND2_X1 U1399 ( .A1(n1830), .A2(n1831), .ZN(U324) );
NAND2_X1 U1400 ( .A1(n1822), .A2(DATA_IN_3_), .ZN(n1831) );
NAND2_X1 U1401 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1823), .ZN(n1830) );
NAND2_X1 U1402 ( .A1(n1832), .A2(n1833), .ZN(U323) );
NAND2_X1 U1403 ( .A1(n1822), .A2(DATA_IN_2_), .ZN(n1833) );
XOR2_X1 U1404 ( .A(n1834), .B(KEYINPUT22), .Z(n1832) );
NAND2_X1 U1405 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1823), .ZN(n1834) );
NAND2_X1 U1406 ( .A1(n1835), .A2(n1836), .ZN(U322) );
NAND2_X1 U1407 ( .A1(n1822), .A2(DATA_IN_1_), .ZN(n1836) );
NAND2_X1 U1408 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1823), .ZN(n1835) );
NAND2_X1 U1409 ( .A1(n1837), .A2(n1838), .ZN(U321) );
NAND2_X1 U1410 ( .A1(n1822), .A2(DATA_IN_0_), .ZN(n1838) );
AND2_X1 U1411 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1839), .ZN(n1822) );
NAND2_X1 U1412 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1823), .ZN(n1837) );
NAND2_X1 U1413 ( .A1(n1719), .A2(n1839), .ZN(n1823) );
NAND2_X1 U1414 ( .A1(n1745), .A2(n1840), .ZN(n1839) );
INV_X1 U1415 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1745) );
INV_X1 U1416 ( .A(U375), .ZN(n1719) );
NOR2_X1 U1417 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1418 ( .A1(n1841), .A2(n1842), .ZN(U320) );
NAND2_X1 U1419 ( .A1(n1694), .A2(DATA_IN_7_), .ZN(n1842) );
NAND2_X1 U1420 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1843), .ZN(n1841) );
NAND2_X1 U1421 ( .A1(n1844), .A2(n1845), .ZN(U319) );
NAND2_X1 U1422 ( .A1(n1694), .A2(DATA_IN_6_), .ZN(n1845) );
NAND2_X1 U1423 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1843), .ZN(n1844) );
NAND2_X1 U1424 ( .A1(n1846), .A2(n1847), .ZN(U318) );
NAND2_X1 U1425 ( .A1(n1694), .A2(DATA_IN_5_), .ZN(n1847) );
NAND2_X1 U1426 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1843), .ZN(n1846) );
NAND2_X1 U1427 ( .A1(n1848), .A2(n1849), .ZN(U317) );
NAND2_X1 U1428 ( .A1(n1694), .A2(DATA_IN_4_), .ZN(n1849) );
NAND2_X1 U1429 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1843), .ZN(n1848) );
NAND2_X1 U1430 ( .A1(n1850), .A2(n1851), .ZN(U316) );
NAND2_X1 U1431 ( .A1(n1694), .A2(DATA_IN_3_), .ZN(n1851) );
XOR2_X1 U1432 ( .A(n1852), .B(KEYINPUT15), .Z(n1850) );
NAND2_X1 U1433 ( .A1(n1853), .A2(n1843), .ZN(n1852) );
XOR2_X1 U1434 ( .A(REG1_REG_3__SCAN_IN), .B(KEYINPUT49), .Z(n1853) );
NAND2_X1 U1435 ( .A1(n1854), .A2(n1855), .ZN(U315) );
NAND2_X1 U1436 ( .A1(n1856), .A2(DATA_IN_2_), .ZN(n1855) );
XNOR2_X1 U1437 ( .A(n1694), .B(KEYINPUT0), .ZN(n1856) );
NAND2_X1 U1438 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1843), .ZN(n1854) );
NAND2_X1 U1439 ( .A1(n1857), .A2(n1858), .ZN(U314) );
NAND2_X1 U1440 ( .A1(n1694), .A2(DATA_IN_1_), .ZN(n1858) );
NAND2_X1 U1441 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1843), .ZN(n1857) );
NAND2_X1 U1442 ( .A1(n1859), .A2(n1860), .ZN(U313) );
NAND2_X1 U1443 ( .A1(n1694), .A2(DATA_IN_0_), .ZN(n1860) );
NAND2_X1 U1444 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1843), .ZN(n1859) );
NAND2_X1 U1445 ( .A1(n1861), .A2(n1862), .ZN(U312) );
NAND2_X1 U1446 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1694), .ZN(n1862) );
NAND2_X1 U1447 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1843), .ZN(n1861) );
NAND2_X1 U1448 ( .A1(n1863), .A2(n1864), .ZN(U311) );
NAND2_X1 U1449 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1694), .ZN(n1864) );
NAND2_X1 U1450 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1843), .ZN(n1863) );
NAND2_X1 U1451 ( .A1(n1865), .A2(n1866), .ZN(U310) );
NAND2_X1 U1452 ( .A1(n1867), .A2(n1694), .ZN(n1866) );
XNOR2_X1 U1453 ( .A(REG1_REG_5__SCAN_IN), .B(KEYINPUT18), .ZN(n1867) );
NAND2_X1 U1454 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1843), .ZN(n1865) );
NAND2_X1 U1455 ( .A1(n1868), .A2(n1869), .ZN(U309) );
NAND2_X1 U1456 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1694), .ZN(n1869) );
NAND2_X1 U1457 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1843), .ZN(n1868) );
NAND2_X1 U1458 ( .A1(n1870), .A2(n1871), .ZN(U308) );
NAND2_X1 U1459 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1694), .ZN(n1871) );
NAND2_X1 U1460 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1843), .ZN(n1870) );
NAND2_X1 U1461 ( .A1(n1872), .A2(n1873), .ZN(U307) );
NAND2_X1 U1462 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1694), .ZN(n1873) );
NAND2_X1 U1463 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1843), .ZN(n1872) );
NAND2_X1 U1464 ( .A1(n1874), .A2(n1875), .ZN(U306) );
NAND2_X1 U1465 ( .A1(n1876), .A2(REG1_REG_1__SCAN_IN), .ZN(n1875) );
XNOR2_X1 U1466 ( .A(n1694), .B(KEYINPUT48), .ZN(n1876) );
NAND2_X1 U1467 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1843), .ZN(n1874) );
NAND2_X1 U1468 ( .A1(n1877), .A2(n1878), .ZN(U305) );
NAND2_X1 U1469 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1694), .ZN(n1878) );
NAND2_X1 U1470 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1843), .ZN(n1877) );
NAND2_X1 U1471 ( .A1(n1879), .A2(n1880), .ZN(U304) );
NAND2_X1 U1472 ( .A1(n1881), .A2(REG2_REG_7__SCAN_IN), .ZN(n1880) );
XNOR2_X1 U1473 ( .A(n1694), .B(KEYINPUT36), .ZN(n1881) );
NAND2_X1 U1474 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1843), .ZN(n1879) );
NAND2_X1 U1475 ( .A1(n1882), .A2(n1883), .ZN(U303) );
NAND2_X1 U1476 ( .A1(n1694), .A2(n1884), .ZN(n1883) );
XOR2_X1 U1477 ( .A(REG2_REG_6__SCAN_IN), .B(KEYINPUT1), .Z(n1884) );
NAND2_X1 U1478 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1843), .ZN(n1882) );
NAND2_X1 U1479 ( .A1(n1885), .A2(n1886), .ZN(U302) );
NAND2_X1 U1480 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1843), .ZN(n1886) );
XOR2_X1 U1481 ( .A(n1887), .B(KEYINPUT2), .Z(n1885) );
NAND2_X1 U1482 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1694), .ZN(n1887) );
NAND2_X1 U1483 ( .A1(n1888), .A2(n1889), .ZN(U301) );
NAND2_X1 U1484 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1694), .ZN(n1889) );
NAND2_X1 U1485 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1843), .ZN(n1888) );
NAND2_X1 U1486 ( .A1(n1890), .A2(n1891), .ZN(U300) );
NAND2_X1 U1487 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1694), .ZN(n1891) );
NAND2_X1 U1488 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1843), .ZN(n1890) );
NAND2_X1 U1489 ( .A1(n1892), .A2(n1893), .ZN(U299) );
NAND2_X1 U1490 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1694), .ZN(n1893) );
NAND2_X1 U1491 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1843), .ZN(n1892) );
NAND2_X1 U1492 ( .A1(n1894), .A2(n1895), .ZN(U298) );
NAND2_X1 U1493 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1694), .ZN(n1895) );
NAND2_X1 U1494 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1843), .ZN(n1894) );
NAND2_X1 U1495 ( .A1(n1896), .A2(n1897), .ZN(U297) );
NAND2_X1 U1496 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1843), .ZN(n1897) );
XOR2_X1 U1497 ( .A(KEYINPUT3), .B(n1898), .Z(n1896) );
AND2_X1 U1498 ( .A1(n1694), .A2(REG2_REG_0__SCAN_IN), .ZN(n1898) );
NAND2_X1 U1499 ( .A1(n1899), .A2(n1900), .ZN(U296) );
NAND2_X1 U1500 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1694), .ZN(n1900) );
NAND2_X1 U1501 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1843), .ZN(n1899) );
NAND2_X1 U1502 ( .A1(n1901), .A2(n1902), .ZN(U295) );
NAND2_X1 U1503 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1694), .ZN(n1902) );
NAND2_X1 U1504 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1843), .ZN(n1901) );
NAND2_X1 U1505 ( .A1(n1903), .A2(n1904), .ZN(U294) );
NAND2_X1 U1506 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1694), .ZN(n1904) );
NAND2_X1 U1507 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1843), .ZN(n1903) );
NAND2_X1 U1508 ( .A1(n1905), .A2(n1906), .ZN(U293) );
NAND2_X1 U1509 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1694), .ZN(n1906) );
NAND2_X1 U1510 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1843), .ZN(n1905) );
NAND2_X1 U1511 ( .A1(n1907), .A2(n1908), .ZN(U292) );
NAND2_X1 U1512 ( .A1(n1909), .A2(n1843), .ZN(n1908) );
XNOR2_X1 U1513 ( .A(n1910), .B(KEYINPUT8), .ZN(n1909) );
NAND2_X1 U1514 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1694), .ZN(n1907) );
NAND2_X1 U1515 ( .A1(n1911), .A2(n1912), .ZN(U291) );
NAND2_X1 U1516 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1694), .ZN(n1912) );
NAND2_X1 U1517 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1843), .ZN(n1911) );
NAND2_X1 U1518 ( .A1(n1913), .A2(n1914), .ZN(U290) );
NAND2_X1 U1519 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1694), .ZN(n1914) );
NAND2_X1 U1520 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1843), .ZN(n1913) );
NAND2_X1 U1521 ( .A1(n1915), .A2(n1916), .ZN(U289) );
NAND2_X1 U1522 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1694), .ZN(n1916) );
NAND2_X1 U1523 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1843), .ZN(n1915) );
NAND3_X1 U1524 ( .A1(n1917), .A2(n1918), .A3(n1919), .ZN(U288) );
NOR3_X1 U1525 ( .A1(n1920), .A2(n1921), .A3(n1922), .ZN(n1919) );
NOR3_X1 U1526 ( .A1(n1923), .A2(n1924), .A3(n1925), .ZN(n1922) );
XNOR2_X1 U1527 ( .A(KEYINPUT60), .B(n1926), .ZN(n1923) );
AND2_X1 U1528 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1927), .ZN(n1920) );
NAND2_X1 U1529 ( .A1(n1928), .A2(REG4_REG_7__SCAN_IN), .ZN(n1918) );
NAND2_X1 U1530 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1843), .ZN(n1917) );
NAND4_X1 U1531 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(U287));
NOR3_X1 U1532 ( .A1(n1933), .A2(n1921), .A3(n1934), .ZN(n1932) );
NOR3_X1 U1533 ( .A1(n1935), .A2(n1936), .A3(n1937), .ZN(n1934) );
NOR3_X1 U1534 ( .A1(n1938), .A2(n1939), .A3(n1937), .ZN(n1921) );
NOR2_X1 U1535 ( .A1(n1940), .A2(n1925), .ZN(n1933) );
XOR2_X1 U1536 ( .A(n1941), .B(n1942), .Z(n1940) );
XNOR2_X1 U1537 ( .A(KEYINPUT25), .B(n1926), .ZN(n1942) );
NAND2_X1 U1538 ( .A1(KEYINPUT60), .A2(n1943), .ZN(n1941) );
NAND2_X1 U1539 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1843), .ZN(n1931) );
NAND2_X1 U1540 ( .A1(n1927), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1930) );
NAND2_X1 U1541 ( .A1(n1928), .A2(REG4_REG_6__SCAN_IN), .ZN(n1929) );
NAND4_X1 U1542 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .ZN(U286));
NOR3_X1 U1543 ( .A1(n1948), .A2(n1949), .A3(n1950), .ZN(n1947) );
NOR3_X1 U1544 ( .A1(n1937), .A2(n1939), .A3(n1951), .ZN(n1950) );
NOR3_X1 U1545 ( .A1(n1952), .A2(n1953), .A3(n1936), .ZN(n1951) );
NOR2_X1 U1546 ( .A1(n1954), .A2(n1955), .ZN(n1952) );
INV_X1 U1547 ( .A(n1935), .ZN(n1939) );
NAND2_X1 U1548 ( .A1(n1953), .A2(n1956), .ZN(n1935) );
NAND2_X1 U1549 ( .A1(n1957), .A2(n1938), .ZN(n1956) );
INV_X1 U1550 ( .A(n1936), .ZN(n1938) );
NOR2_X1 U1551 ( .A1(n1958), .A2(n1959), .ZN(n1936) );
NAND2_X1 U1552 ( .A1(n1959), .A2(n1958), .ZN(n1957) );
NOR3_X1 U1553 ( .A1(n1925), .A2(n1924), .A3(n1960), .ZN(n1949) );
NOR2_X1 U1554 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
INV_X1 U1555 ( .A(n1943), .ZN(n1924) );
NAND2_X1 U1556 ( .A1(n1963), .A2(n1964), .ZN(n1943) );
XNOR2_X1 U1557 ( .A(n1961), .B(KEYINPUT5), .ZN(n1964) );
XOR2_X1 U1558 ( .A(n1962), .B(KEYINPUT38), .Z(n1963) );
NAND2_X1 U1559 ( .A1(n1926), .A2(n1965), .ZN(n1962) );
NAND2_X1 U1560 ( .A1(n1959), .A2(n1966), .ZN(n1965) );
OR2_X1 U1561 ( .A1(n1966), .A2(n1959), .ZN(n1926) );
INV_X1 U1562 ( .A(n1955), .ZN(n1959) );
NOR2_X1 U1563 ( .A1(n1955), .A2(n1967), .ZN(n1948) );
NAND2_X1 U1564 ( .A1(n1968), .A2(n1969), .ZN(n1955) );
NAND3_X1 U1565 ( .A1(n1970), .A2(n1971), .A3(n1972), .ZN(n1969) );
XOR2_X1 U1566 ( .A(n1973), .B(n1974), .Z(n1972) );
NAND2_X1 U1567 ( .A1(n1975), .A2(n1976), .ZN(n1971) );
XNOR2_X1 U1568 ( .A(n1977), .B(KEYINPUT11), .ZN(n1976) );
NAND2_X1 U1569 ( .A1(n1978), .A2(n1979), .ZN(n1970) );
NAND2_X1 U1570 ( .A1(n1980), .A2(n1981), .ZN(n1979) );
XNOR2_X1 U1571 ( .A(KEYINPUT31), .B(n1982), .ZN(n1980) );
NAND3_X1 U1572 ( .A1(n1983), .A2(n1984), .A3(n1985), .ZN(n1968) );
XOR2_X1 U1573 ( .A(n1986), .B(n1973), .Z(n1985) );
NAND2_X1 U1574 ( .A1(n1987), .A2(n1988), .ZN(n1973) );
NAND2_X1 U1575 ( .A1(DATA_IN_6_), .A2(n1989), .ZN(n1988) );
NAND2_X1 U1576 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1987) );
NAND2_X1 U1577 ( .A1(KEYINPUT33), .A2(n1974), .ZN(n1986) );
NAND2_X1 U1578 ( .A1(n1990), .A2(n1991), .ZN(n1974) );
NAND2_X1 U1579 ( .A1(RESTART), .A2(n1788), .ZN(n1991) );
INV_X1 U1580 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1788) );
NAND2_X1 U1581 ( .A1(n1992), .A2(n1989), .ZN(n1990) );
NAND2_X1 U1582 ( .A1(n1993), .A2(n1994), .ZN(n1984) );
NAND2_X1 U1583 ( .A1(n1975), .A2(n1977), .ZN(n1993) );
INV_X1 U1584 ( .A(n1982), .ZN(n1975) );
NAND2_X1 U1585 ( .A1(n1981), .A2(n1982), .ZN(n1983) );
NAND2_X1 U1586 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1843), .ZN(n1946) );
NAND2_X1 U1587 ( .A1(n1927), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1945) );
NAND2_X1 U1588 ( .A1(n1928), .A2(REG4_REG_5__SCAN_IN), .ZN(n1944) );
NAND4_X1 U1589 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .ZN(U285));
NOR3_X1 U1590 ( .A1(n1999), .A2(n2000), .A3(n2001), .ZN(n1998) );
NOR3_X1 U1591 ( .A1(n1925), .A2(n1961), .A3(n2002), .ZN(n2001) );
NOR2_X1 U1592 ( .A1(n2003), .A2(n2004), .ZN(n2002) );
XOR2_X1 U1593 ( .A(KEYINPUT50), .B(n2005), .Z(n2004) );
AND2_X1 U1594 ( .A1(n2005), .A2(n2003), .ZN(n1961) );
NAND2_X1 U1595 ( .A1(n1966), .A2(n2006), .ZN(n2003) );
NAND2_X1 U1596 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
OR2_X1 U1597 ( .A1(n2008), .A2(n2007), .ZN(n1966) );
NOR3_X1 U1598 ( .A1(n1937), .A2(n1953), .A3(n2009), .ZN(n2000) );
NOR2_X1 U1599 ( .A1(n2010), .A2(n2011), .ZN(n2009) );
AND2_X1 U1600 ( .A1(n2012), .A2(n2013), .ZN(n2010) );
AND3_X1 U1601 ( .A1(n2014), .A2(n2012), .A3(n2013), .ZN(n1953) );
XNOR2_X1 U1602 ( .A(KEYINPUT40), .B(n2011), .ZN(n2014) );
NAND2_X1 U1603 ( .A1(n1958), .A2(n2015), .ZN(n2011) );
NAND2_X1 U1604 ( .A1(n2007), .A2(n2016), .ZN(n2015) );
INV_X1 U1605 ( .A(n1954), .ZN(n1958) );
NOR2_X1 U1606 ( .A1(n2016), .A2(n2007), .ZN(n1954) );
AND2_X1 U1607 ( .A1(n2007), .A2(n2017), .ZN(n1999) );
XOR2_X1 U1608 ( .A(n2018), .B(n1982), .Z(n2007) );
NAND2_X1 U1609 ( .A1(n2019), .A2(n2020), .ZN(n1982) );
NAND2_X1 U1610 ( .A1(RESTART), .A2(n1769), .ZN(n2020) );
NAND2_X1 U1611 ( .A1(n2021), .A2(n1989), .ZN(n2019) );
XNOR2_X1 U1612 ( .A(n1978), .B(n1977), .ZN(n2018) );
INV_X1 U1613 ( .A(n1981), .ZN(n1977) );
NAND2_X1 U1614 ( .A1(n2022), .A2(n2023), .ZN(n1981) );
NAND2_X1 U1615 ( .A1(RESTART), .A2(n1704), .ZN(n2023) );
NAND2_X1 U1616 ( .A1(n1801), .A2(n1989), .ZN(n2022) );
INV_X1 U1617 ( .A(DATA_IN_5_), .ZN(n1801) );
INV_X1 U1618 ( .A(n1994), .ZN(n1978) );
NAND2_X1 U1619 ( .A1(n2024), .A2(n2025), .ZN(n1994) );
NAND2_X1 U1620 ( .A1(n2026), .A2(n2027), .ZN(n2025) );
OR2_X1 U1621 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
NAND2_X1 U1622 ( .A1(n2029), .A2(n2028), .ZN(n2024) );
NAND2_X1 U1623 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1843), .ZN(n1997) );
NAND2_X1 U1624 ( .A1(n1927), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1996) );
NAND2_X1 U1625 ( .A1(n1928), .A2(REG4_REG_4__SCAN_IN), .ZN(n1995) );
NAND4_X1 U1626 ( .A1(n2030), .A2(n2031), .A3(n2032), .A4(n2033), .ZN(U284));
NOR3_X1 U1627 ( .A1(n2034), .A2(n2035), .A3(n2036), .ZN(n2033) );
NOR2_X1 U1628 ( .A1(n1910), .A2(n2037), .ZN(n2036) );
AND2_X1 U1629 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1927), .ZN(n2035) );
XOR2_X1 U1630 ( .A(n2038), .B(KEYINPUT34), .Z(n2034) );
NAND2_X1 U1631 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1843), .ZN(n2038) );
NAND2_X1 U1632 ( .A1(n2017), .A2(n2039), .ZN(n2032) );
NAND3_X1 U1633 ( .A1(n2040), .A2(n2041), .A3(n2042), .ZN(n2031) );
XNOR2_X1 U1634 ( .A(KEYINPUT57), .B(n1925), .ZN(n2042) );
NAND2_X1 U1635 ( .A1(n2043), .A2(n2044), .ZN(n2041) );
NAND2_X1 U1636 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
NAND2_X1 U1637 ( .A1(KEYINPUT41), .A2(n2047), .ZN(n2046) );
INV_X1 U1638 ( .A(n2048), .ZN(n2043) );
NAND2_X1 U1639 ( .A1(n2005), .A2(n2049), .ZN(n2040) );
INV_X1 U1640 ( .A(KEYINPUT41), .ZN(n2049) );
AND2_X1 U1641 ( .A1(n2047), .A2(n2048), .ZN(n2005) );
NAND2_X1 U1642 ( .A1(n2008), .A2(n2050), .ZN(n2048) );
OR2_X1 U1643 ( .A1(n2051), .A2(n2039), .ZN(n2008) );
XOR2_X1 U1644 ( .A(n2045), .B(KEYINPUT12), .Z(n2047) );
NAND2_X1 U1645 ( .A1(n2052), .A2(n2053), .ZN(n2030) );
XOR2_X1 U1646 ( .A(n2012), .B(n2013), .Z(n2052) );
NAND2_X1 U1647 ( .A1(n2016), .A2(n2050), .ZN(n2012) );
NAND2_X1 U1648 ( .A1(n2039), .A2(n2051), .ZN(n2050) );
INV_X1 U1649 ( .A(n2054), .ZN(n2051) );
NAND2_X1 U1650 ( .A1(n2054), .A2(n2055), .ZN(n2016) );
XNOR2_X1 U1651 ( .A(n2039), .B(KEYINPUT47), .ZN(n2055) );
XOR2_X1 U1652 ( .A(n2056), .B(n2028), .Z(n2039) );
NAND2_X1 U1653 ( .A1(n2057), .A2(n2058), .ZN(n2028) );
NAND2_X1 U1654 ( .A1(RESTART), .A2(n1708), .ZN(n2058) );
NAND2_X1 U1655 ( .A1(n1773), .A2(n1989), .ZN(n2057) );
XNOR2_X1 U1656 ( .A(n2029), .B(n2026), .ZN(n2056) );
AND2_X1 U1657 ( .A1(n2059), .A2(n2060), .ZN(n2026) );
NAND2_X1 U1658 ( .A1(n2061), .A2(n2062), .ZN(n2060) );
NAND2_X1 U1659 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
OR2_X1 U1660 ( .A1(n2063), .A2(n2064), .ZN(n2059) );
AND3_X1 U1661 ( .A1(n2065), .A2(n2066), .A3(n2067), .ZN(n2029) );
NAND2_X1 U1662 ( .A1(KEYINPUT54), .A2(n1786), .ZN(n2067) );
NAND3_X1 U1663 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n2068), .A3(RESTART), .ZN(n2066) );
NAND2_X1 U1664 ( .A1(n2069), .A2(n1989), .ZN(n2065) );
NAND2_X1 U1665 ( .A1(n2070), .A2(n2068), .ZN(n2069) );
INV_X1 U1666 ( .A(KEYINPUT54), .ZN(n2068) );
NAND4_X1 U1667 ( .A1(n2071), .A2(n2072), .A3(n2073), .A4(n2074), .ZN(U283));
NOR3_X1 U1668 ( .A1(n2075), .A2(n2076), .A3(n2077), .ZN(n2074) );
NOR3_X1 U1669 ( .A1(n1925), .A2(n2045), .A3(n2078), .ZN(n2077) );
NOR2_X1 U1670 ( .A1(n2079), .A2(n2080), .ZN(n2078) );
NOR2_X1 U1671 ( .A1(n2081), .A2(n2082), .ZN(n2079) );
AND3_X1 U1672 ( .A1(n2080), .A2(n2083), .A3(n2084), .ZN(n2045) );
XNOR2_X1 U1673 ( .A(n2082), .B(KEYINPUT37), .ZN(n2084) );
AND3_X1 U1674 ( .A1(n2085), .A2(n2086), .A3(n2087), .ZN(n2080) );
OR2_X1 U1675 ( .A1(n2088), .A2(KEYINPUT21), .ZN(n2087) );
NAND4_X1 U1676 ( .A1(KEYINPUT10), .A2(n2088), .A3(KEYINPUT21), .A4(n2089),
.ZN(n2086) );
NAND2_X1 U1677 ( .A1(n2090), .A2(n2091), .ZN(n2085) );
NAND2_X1 U1678 ( .A1(KEYINPUT10), .A2(n2088), .ZN(n2090) );
NOR3_X1 U1679 ( .A1(n2092), .A2(n2013), .A3(n2093), .ZN(n2076) );
NOR2_X1 U1680 ( .A1(n2094), .A2(n2095), .ZN(n2093) );
AND2_X1 U1681 ( .A1(n2094), .A2(n2096), .ZN(n2013) );
OR2_X1 U1682 ( .A1(n2054), .A2(n2095), .ZN(n2096) );
NOR2_X1 U1683 ( .A1(n2097), .A2(n2089), .ZN(n2095) );
NOR2_X1 U1684 ( .A1(n2091), .A2(n2088), .ZN(n2054) );
NOR2_X1 U1685 ( .A1(n2098), .A2(n2081), .ZN(n2094) );
XNOR2_X1 U1686 ( .A(n2053), .B(KEYINPUT32), .ZN(n2092) );
NOR2_X1 U1687 ( .A1(n2097), .A2(n1967), .ZN(n2075) );
INV_X1 U1688 ( .A(n2088), .ZN(n2097) );
XOR2_X1 U1689 ( .A(n2099), .B(n2064), .Z(n2088) );
NAND2_X1 U1690 ( .A1(n2100), .A2(n2101), .ZN(n2064) );
NAND2_X1 U1691 ( .A1(RESTART), .A2(n1777), .ZN(n2101) );
NAND2_X1 U1692 ( .A1(n1910), .A2(n1989), .ZN(n2100) );
NAND2_X1 U1693 ( .A1(n2102), .A2(n2103), .ZN(n2099) );
NAND2_X1 U1694 ( .A1(n2061), .A2(n2104), .ZN(n2103) );
NAND2_X1 U1695 ( .A1(KEYINPUT62), .A2(n2063), .ZN(n2104) );
INV_X1 U1696 ( .A(n2105), .ZN(n2061) );
NAND2_X1 U1697 ( .A1(n2063), .A2(n2105), .ZN(n2102) );
NAND2_X1 U1698 ( .A1(n2106), .A2(n2107), .ZN(n2105) );
NAND2_X1 U1699 ( .A1(n2108), .A2(n2109), .ZN(n2107) );
NAND2_X1 U1700 ( .A1(n2110), .A2(n2111), .ZN(n2108) );
XOR2_X1 U1701 ( .A(n2112), .B(KEYINPUT43), .Z(n2111) );
INV_X1 U1702 ( .A(n2113), .ZN(n2110) );
NAND2_X1 U1703 ( .A1(n2113), .A2(n2112), .ZN(n2106) );
NAND2_X1 U1704 ( .A1(n2114), .A2(n2115), .ZN(n2063) );
NAND2_X1 U1705 ( .A1(RESTART), .A2(n1818), .ZN(n2115) );
NAND2_X1 U1706 ( .A1(n1785), .A2(n1989), .ZN(n2114) );
NAND2_X1 U1707 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1843), .ZN(n2073) );
NAND2_X1 U1708 ( .A1(n1927), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2072) );
NAND2_X1 U1709 ( .A1(n1928), .A2(REG4_REG_2__SCAN_IN), .ZN(n2071) );
NAND4_X1 U1710 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(U282));
NOR4_X1 U1711 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2119));
AND2_X1 U1712 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1843), .ZN(n2123) );
AND2_X1 U1713 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1927), .ZN(n2122) );
NOR3_X1 U1714 ( .A1(n2083), .A2(n2098), .A3(n1937), .ZN(n2121) );
INV_X1 U1715 ( .A(n2053), .ZN(n1937) );
NOR2_X1 U1716 ( .A1(n2081), .A2(n2124), .ZN(n2120) );
NAND2_X1 U1717 ( .A1(n2017), .A2(n2125), .ZN(n2118) );
INV_X1 U1718 ( .A(n1967), .ZN(n2017) );
NAND2_X1 U1719 ( .A1(n2126), .A2(n1928), .ZN(n2117) );
XNOR2_X1 U1720 ( .A(REG4_REG_1__SCAN_IN), .B(KEYINPUT56), .ZN(n2126) );
NAND3_X1 U1721 ( .A1(n2127), .A2(n2128), .A3(n2129), .ZN(n2116) );
OR2_X1 U1722 ( .A1(n2082), .A2(KEYINPUT61), .ZN(n2128) );
NAND2_X1 U1723 ( .A1(KEYINPUT61), .A2(n2130), .ZN(n2127) );
NAND2_X1 U1724 ( .A1(n2081), .A2(n2131), .ZN(n2130) );
INV_X1 U1725 ( .A(n2083), .ZN(n2081) );
NAND2_X1 U1726 ( .A1(n2091), .A2(n2132), .ZN(n2083) );
NAND2_X1 U1727 ( .A1(n2125), .A2(n2133), .ZN(n2132) );
INV_X1 U1728 ( .A(n2089), .ZN(n2091) );
NOR2_X1 U1729 ( .A1(n2133), .A2(n2125), .ZN(n2089) );
XOR2_X1 U1730 ( .A(n2134), .B(n2113), .Z(n2125) );
NAND2_X1 U1731 ( .A1(n2135), .A2(n2136), .ZN(n2113) );
NAND2_X1 U1732 ( .A1(RESTART), .A2(n1813), .ZN(n2136) );
NAND2_X1 U1733 ( .A1(n1714), .A2(n1989), .ZN(n2135) );
XNOR2_X1 U1734 ( .A(n2109), .B(n2112), .ZN(n2134) );
NAND2_X1 U1735 ( .A1(n2137), .A2(n2138), .ZN(n2112) );
NAND2_X1 U1736 ( .A1(RESTART), .A2(n1784), .ZN(n2138) );
NAND2_X1 U1737 ( .A1(n2139), .A2(n1989), .ZN(n2137) );
NAND2_X1 U1738 ( .A1(n2140), .A2(n2141), .ZN(n2109) );
NAND2_X1 U1739 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
NAND2_X1 U1740 ( .A1(n2144), .A2(n2145), .ZN(n2142) );
OR2_X1 U1741 ( .A1(n2144), .A2(n2145), .ZN(n2140) );
NAND4_X1 U1742 ( .A1(n2124), .A2(n2146), .A3(n2147), .A4(n2148), .ZN(U281));
NAND2_X1 U1743 ( .A1(n1928), .A2(REG4_REG_0__SCAN_IN), .ZN(n2148) );
INV_X1 U1744 ( .A(n2037), .ZN(n1928) );
NAND2_X1 U1745 ( .A1(n2149), .A2(AVERAGE), .ZN(n2037) );
NOR2_X1 U1746 ( .A1(n2150), .A2(n2151), .ZN(n2147) );
NOR2_X1 U1747 ( .A1(n2152), .A2(n1967), .ZN(n2151) );
NAND3_X1 U1748 ( .A1(n2153), .A2(n2154), .A3(n2155), .ZN(n1967) );
NAND2_X1 U1749 ( .A1(n2156), .A2(n1989), .ZN(n2153) );
NAND4_X1 U1750 ( .A1(ENABLE), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(n2156));
INV_X1 U1751 ( .A(AVERAGE), .ZN(n2159) );
NAND2_X1 U1752 ( .A1(REG4_REG_7__SCAN_IN), .A2(n2160), .ZN(n2157) );
AND2_X1 U1753 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1927), .ZN(n2150) );
NOR3_X1 U1754 ( .A1(ENABLE), .A2(RESTART), .A3(n2161), .ZN(n1927) );
NAND2_X1 U1755 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1843), .ZN(n2146) );
AND2_X1 U1756 ( .A1(n2162), .A2(n2163), .ZN(n2124) );
NAND2_X1 U1757 ( .A1(n2098), .A2(n2053), .ZN(n2163) );
NOR2_X1 U1758 ( .A1(n2154), .A2(n2161), .ZN(n2053) );
NAND2_X1 U1759 ( .A1(RESTART), .A2(n2164), .ZN(n2154) );
NAND2_X1 U1760 ( .A1(n2165), .A2(n2166), .ZN(n2164) );
NAND3_X1 U1761 ( .A1(n2167), .A2(n2168), .A3(n2169), .ZN(n2166) );
NAND2_X1 U1762 ( .A1(n1794), .A2(n1756), .ZN(n2169) );
INV_X1 U1763 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1756) );
INV_X1 U1764 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1794) );
NAND2_X1 U1765 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2170), .ZN(n2168) );
NAND2_X1 U1766 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
INV_X1 U1767 ( .A(n2173), .ZN(n2172) );
XNOR2_X1 U1768 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT28), .ZN(n2171) );
NAND2_X1 U1769 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2173), .ZN(n2167) );
NAND2_X1 U1770 ( .A1(n2174), .A2(n2175), .ZN(n2173) );
NAND2_X1 U1771 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2175) );
NAND2_X1 U1772 ( .A1(n2176), .A2(n2177), .ZN(n2174) );
NAND2_X1 U1773 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
NAND3_X1 U1774 ( .A1(n2180), .A2(n2181), .A3(n2182), .ZN(n2179) );
NAND2_X1 U1775 ( .A1(n1708), .A2(n1786), .ZN(n2182) );
INV_X1 U1776 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1786) );
INV_X1 U1777 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1708) );
NAND3_X1 U1778 ( .A1(n2183), .A2(n2184), .A3(n2185), .ZN(n2181) );
NAND2_X1 U1779 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2185) );
NAND3_X1 U1780 ( .A1(n2186), .A2(n2187), .A3(n2188), .ZN(n2184) );
XOR2_X1 U1781 ( .A(n2189), .B(KEYINPUT17), .Z(n2188) );
NAND2_X1 U1782 ( .A1(n2190), .A2(n2191), .ZN(n2189) );
NAND2_X1 U1783 ( .A1(n2192), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2191) );
XNOR2_X1 U1784 ( .A(RMIN_REG_0__SCAN_IN), .B(KEYINPUT20), .ZN(n2192) );
XOR2_X1 U1785 ( .A(KEYINPUT23), .B(n2193), .Z(n2190) );
NOR2_X1 U1786 ( .A1(n1816), .A2(n1741), .ZN(n2193) );
NAND2_X1 U1787 ( .A1(n1816), .A2(n1741), .ZN(n2187) );
INV_X1 U1788 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1741) );
INV_X1 U1789 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1816) );
NAND2_X1 U1790 ( .A1(n1813), .A2(n1784), .ZN(n2186) );
INV_X1 U1791 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1784) );
INV_X1 U1792 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1813) );
NAND2_X1 U1793 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2183) );
NAND2_X1 U1794 ( .A1(n1818), .A2(n1777), .ZN(n2180) );
INV_X1 U1795 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1777) );
INV_X1 U1796 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1818) );
NAND2_X1 U1797 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2178) );
XOR2_X1 U1798 ( .A(n2194), .B(KEYINPUT52), .Z(n2176) );
NAND2_X1 U1799 ( .A1(n1769), .A2(n1704), .ZN(n2194) );
INV_X1 U1800 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1704) );
INV_X1 U1801 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1769) );
XOR2_X1 U1802 ( .A(n2195), .B(KEYINPUT14), .Z(n2165) );
NAND2_X1 U1803 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2195) );
AND3_X1 U1804 ( .A1(n2196), .A2(n2197), .A3(n2133), .ZN(n2098) );
OR3_X1 U1805 ( .A1(n2152), .A2(KEYINPUT29), .A3(n2198), .ZN(n2197) );
NAND2_X1 U1806 ( .A1(KEYINPUT29), .A2(n2198), .ZN(n2196) );
NAND2_X1 U1807 ( .A1(n2129), .A2(n2082), .ZN(n2162) );
INV_X1 U1808 ( .A(n2131), .ZN(n2082) );
NAND3_X1 U1809 ( .A1(n2199), .A2(n2200), .A3(n2133), .ZN(n2131) );
NAND2_X1 U1810 ( .A1(n2198), .A2(n2152), .ZN(n2133) );
OR3_X1 U1811 ( .A1(n2198), .A2(KEYINPUT4), .A3(n2152), .ZN(n2200) );
XNOR2_X1 U1812 ( .A(n2201), .B(n2202), .ZN(n2198) );
NOR2_X1 U1813 ( .A1(KEYINPUT46), .A2(n2203), .ZN(n2202) );
NAND2_X1 U1814 ( .A1(KEYINPUT4), .A2(n2152), .ZN(n2199) );
XNOR2_X1 U1815 ( .A(n2204), .B(n2144), .ZN(n2152) );
NAND2_X1 U1816 ( .A1(n2205), .A2(n2206), .ZN(n2144) );
NAND2_X1 U1817 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1989), .ZN(n2206) );
NAND2_X1 U1818 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2205) );
XNOR2_X1 U1819 ( .A(n2143), .B(n2145), .ZN(n2204) );
NAND3_X1 U1820 ( .A1(n2207), .A2(n2208), .A3(n2209), .ZN(n2145) );
OR2_X1 U1821 ( .A1(KEYINPUT7), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2209) );
NAND3_X1 U1822 ( .A1(KEYINPUT7), .A2(RMAX_REG_1__SCAN_IN), .A3(RESTART),
.ZN(n2208) );
NAND2_X1 U1823 ( .A1(n2210), .A2(n1989), .ZN(n2207) );
NAND2_X1 U1824 ( .A1(KEYINPUT7), .A2(n1783), .ZN(n2210) );
NAND2_X1 U1825 ( .A1(n2211), .A2(n2201), .ZN(n2143) );
NAND2_X1 U1826 ( .A1(n2212), .A2(n2213), .ZN(n2201) );
NAND2_X1 U1827 ( .A1(DATA_IN_0_), .A2(n1989), .ZN(n2213) );
NAND2_X1 U1828 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2212) );
XOR2_X1 U1829 ( .A(n2203), .B(KEYINPUT63), .Z(n2211) );
NAND2_X1 U1830 ( .A1(n2214), .A2(n2215), .ZN(n2203) );
NAND2_X1 U1831 ( .A1(n2216), .A2(n1989), .ZN(n2215) );
INV_X1 U1832 ( .A(RESTART), .ZN(n1989) );
NAND2_X1 U1833 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2217), .ZN(n2216) );
NAND2_X1 U1834 ( .A1(n2218), .A2(n2219), .ZN(n2214) );
INV_X1 U1835 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2219) );
NAND2_X1 U1836 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2220), .ZN(n2218) );
NAND2_X1 U1837 ( .A1(RESTART), .A2(n2217), .ZN(n2220) );
INV_X1 U1838 ( .A(KEYINPUT39), .ZN(n2217) );
INV_X1 U1839 ( .A(n1925), .ZN(n2129) );
NAND4_X1 U1840 ( .A1(n2221), .A2(n2149), .A3(n2222), .A4(n2160), .ZN(n1925));
NAND3_X1 U1841 ( .A1(n2223), .A2(n1757), .A3(n2224), .ZN(n2160) );
NAND2_X1 U1842 ( .A1(n2225), .A2(n1992), .ZN(n2224) );
INV_X1 U1843 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1992) );
INV_X1 U1844 ( .A(DATA_IN_7_), .ZN(n1757) );
NAND2_X1 U1845 ( .A1(n2158), .A2(n2226), .ZN(n2222) );
INV_X1 U1846 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2226) );
NAND3_X1 U1847 ( .A1(n2225), .A2(n2227), .A3(DATA_IN_7_), .ZN(n2158) );
NAND2_X1 U1848 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2223), .ZN(n2227) );
NAND2_X1 U1849 ( .A1(n2228), .A2(n1764), .ZN(n2223) );
INV_X1 U1850 ( .A(DATA_IN_6_), .ZN(n1764) );
XOR2_X1 U1851 ( .A(KEYINPUT6), .B(n2229), .Z(n2228) );
NAND2_X1 U1852 ( .A1(n2229), .A2(DATA_IN_6_), .ZN(n2225) );
AND2_X1 U1853 ( .A1(n2230), .A2(n2231), .ZN(n2229) );
NAND2_X1 U1854 ( .A1(n2021), .A2(n2232), .ZN(n2231) );
NAND2_X1 U1855 ( .A1(DATA_IN_5_), .A2(n2233), .ZN(n2232) );
INV_X1 U1856 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2021) );
OR2_X1 U1857 ( .A1(n2233), .A2(DATA_IN_5_), .ZN(n2230) );
NAND2_X1 U1858 ( .A1(n2234), .A2(n2235), .ZN(n2233) );
NAND2_X1 U1859 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2235) );
NAND3_X1 U1860 ( .A1(n2236), .A2(n2237), .A3(n2238), .ZN(n2234) );
NAND2_X1 U1861 ( .A1(n1773), .A2(n2070), .ZN(n2238) );
INV_X1 U1862 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2070) );
INV_X1 U1863 ( .A(DATA_IN_4_), .ZN(n1773) );
NAND3_X1 U1864 ( .A1(n2239), .A2(n2240), .A3(n2241), .ZN(n2237) );
NAND2_X1 U1865 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2241) );
NAND3_X1 U1866 ( .A1(n2242), .A2(n2243), .A3(n2244), .ZN(n2240) );
NAND2_X1 U1867 ( .A1(n1714), .A2(n2139), .ZN(n2244) );
INV_X1 U1868 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2139) );
INV_X1 U1869 ( .A(DATA_IN_2_), .ZN(n1714) );
NAND2_X1 U1870 ( .A1(n2245), .A2(n2246), .ZN(n2243) );
INV_X1 U1871 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2246) );
OR2_X1 U1872 ( .A1(n2247), .A2(n1783), .ZN(n2245) );
NAND2_X1 U1873 ( .A1(n2247), .A2(n1783), .ZN(n2242) );
INV_X1 U1874 ( .A(DATA_IN_1_), .ZN(n1783) );
NAND2_X1 U1875 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2247) );
NAND2_X1 U1876 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2239) );
NAND2_X1 U1877 ( .A1(n1785), .A2(n1910), .ZN(n2236) );
INV_X1 U1878 ( .A(REG4_REG_3__SCAN_IN), .ZN(n1910) );
INV_X1 U1879 ( .A(DATA_IN_3_), .ZN(n1785) );
NOR3_X1 U1880 ( .A1(n2161), .A2(RESTART), .A3(n1840), .ZN(n2149) );
INV_X1 U1881 ( .A(ENABLE), .ZN(n1840) );
INV_X1 U1882 ( .A(n2155), .ZN(n2161) );
NOR2_X1 U1883 ( .A1(n2248), .A2(n1843), .ZN(n2155) );
XNOR2_X1 U1884 ( .A(AVERAGE), .B(KEYINPUT59), .ZN(n2221) );
NAND2_X1 U1885 ( .A1(n1693), .A2(n2249), .ZN(U280) );
NAND2_X1 U1886 ( .A1(STATO_REG_0__SCAN_IN), .A2(n2248), .ZN(n2249) );
INV_X1 U1887 ( .A(STATO_REG_1__SCAN_IN), .ZN(n2248) );
endmodule


