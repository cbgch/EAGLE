//Key = 0010110111101111011001000110101110101100000001110010111001011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359;

XNOR2_X1 U743 ( .A(G107), .B(n1028), .ZN(G9) );
OR3_X1 U744 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1034) );
NAND2_X1 U748 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND4_X1 U750 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NOR3_X1 U752 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1048) );
XOR2_X1 U754 ( .A(n1055), .B(KEYINPUT6), .Z(n1042) );
NAND4_X1 U755 ( .A1(n1056), .A2(n1045), .A3(n1047), .A4(n1057), .ZN(n1055) );
INV_X1 U756 ( .A(n1058), .ZN(n1045) );
XNOR2_X1 U757 ( .A(n1053), .B(KEYINPUT13), .ZN(n1056) );
NAND4_X1 U758 ( .A1(n1059), .A2(n1054), .A3(n1046), .A4(n1060), .ZN(n1037) );
NOR2_X1 U759 ( .A1(n1061), .A2(n1058), .ZN(n1060) );
NAND2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1040), .A2(n1064), .ZN(n1063) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1047), .A2(n1069), .ZN(n1062) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U767 ( .A1(n1035), .A2(G952), .A3(n1074), .ZN(n1032) );
INV_X1 U768 ( .A(n1038), .ZN(n1074) );
NAND4_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1038) );
NOR4_X1 U770 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1068), .ZN(n1078) );
XOR2_X1 U771 ( .A(n1082), .B(KEYINPUT25), .Z(n1079) );
NAND2_X1 U772 ( .A1(G469), .A2(n1083), .ZN(n1082) );
NOR3_X1 U773 ( .A1(n1084), .A2(n1050), .A3(n1072), .ZN(n1077) );
NOR2_X1 U774 ( .A1(G469), .A2(n1083), .ZN(n1084) );
XNOR2_X1 U775 ( .A(n1085), .B(n1086), .ZN(n1076) );
NOR2_X1 U776 ( .A1(n1087), .A2(KEYINPUT3), .ZN(n1086) );
INV_X1 U777 ( .A(n1088), .ZN(n1087) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1075) );
NOR2_X1 U779 ( .A1(n1091), .A2(KEYINPUT58), .ZN(n1090) );
INV_X1 U780 ( .A(n1092), .ZN(n1035) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(G72) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U783 ( .A1(n1097), .A2(KEYINPUT22), .A3(G953), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U785 ( .A(KEYINPUT55), .B(n1100), .ZN(n1099) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1095) );
NAND2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U788 ( .A(G953), .B(KEYINPUT7), .ZN(n1103) );
XOR2_X1 U789 ( .A(n1105), .B(n1106), .Z(n1101) );
XOR2_X1 U790 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U791 ( .A(n1109), .B(G131), .Z(n1108) );
NAND2_X1 U792 ( .A1(KEYINPUT18), .A2(n1110), .ZN(n1109) );
XOR2_X1 U793 ( .A(G134), .B(n1111), .Z(n1105) );
XOR2_X1 U794 ( .A(KEYINPUT39), .B(G137), .Z(n1111) );
NAND2_X1 U795 ( .A1(G953), .A2(n1112), .ZN(n1093) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(G69) );
XOR2_X1 U798 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U799 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U802 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U803 ( .A(KEYINPUT38), .B(n1121), .Z(n1118) );
AND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1130), .ZN(G63) );
NOR3_X1 U809 ( .A1(n1091), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR3_X1 U810 ( .A1(n1133), .A2(n1089), .A3(n1129), .ZN(n1132) );
INV_X1 U811 ( .A(n1134), .ZN(n1133) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1134), .ZN(n1131) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1089), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1137), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1129), .ZN(n1139) );
XNOR2_X1 U817 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1124), .A2(n1142), .ZN(G57) );
NOR2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U820 ( .A(KEYINPUT43), .B(n1145), .Z(n1144) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U822 ( .A(n1148), .B(KEYINPUT29), .Z(n1147) );
AND2_X1 U823 ( .A1(n1148), .A2(n1146), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1149) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1129), .ZN(n1154) );
OR2_X1 U828 ( .A1(n1152), .A2(n1151), .ZN(n1153) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U831 ( .A1(KEYINPUT52), .A2(n1160), .ZN(n1158) );
NAND2_X1 U832 ( .A1(KEYINPUT15), .A2(n1161), .ZN(n1160) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1156) );
NAND2_X1 U834 ( .A1(KEYINPUT15), .A2(n1164), .ZN(n1163) );
NAND2_X1 U835 ( .A1(n1165), .A2(KEYINPUT52), .ZN(n1164) );
INV_X1 U836 ( .A(n1159), .ZN(n1165) );
NAND3_X1 U837 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1159) );
OR2_X1 U838 ( .A1(n1169), .A2(KEYINPUT54), .ZN(n1168) );
NAND3_X1 U839 ( .A1(KEYINPUT54), .A2(n1169), .A3(n1170), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1166) );
NAND2_X1 U841 ( .A1(KEYINPUT54), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U842 ( .A(KEYINPUT36), .B(n1169), .ZN(n1173) );
INV_X1 U843 ( .A(KEYINPUT12), .ZN(n1152) );
NOR2_X1 U844 ( .A1(n1124), .A2(n1174), .ZN(G54) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1177), .B(n1107), .ZN(n1176) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1175) );
XNOR2_X1 U848 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1182), .A2(n1129), .ZN(n1181) );
NOR2_X1 U850 ( .A1(n1183), .A2(n1184), .ZN(G51) );
XOR2_X1 U851 ( .A(n1121), .B(n1185), .Z(n1184) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U853 ( .A1(n1088), .A2(n1129), .ZN(n1187) );
NAND2_X1 U854 ( .A1(G902), .A2(n1036), .ZN(n1129) );
INV_X1 U855 ( .A(n1136), .ZN(n1036) );
NOR3_X1 U856 ( .A1(n1098), .A2(n1188), .A3(n1122), .ZN(n1136) );
NAND2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1122) );
AND4_X1 U858 ( .A1(n1191), .A2(n1141), .A3(n1192), .A4(n1193), .ZN(n1190) );
OR3_X1 U859 ( .A1(n1029), .A2(n1030), .A3(n1194), .ZN(n1141) );
NOR4_X1 U860 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1189) );
NOR3_X1 U861 ( .A1(n1031), .A2(n1199), .A3(n1029), .ZN(n1198) );
XNOR2_X1 U862 ( .A(n1047), .B(KEYINPUT33), .ZN(n1199) );
INV_X1 U863 ( .A(n1051), .ZN(n1031) );
NAND4_X1 U864 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1098) );
NOR4_X1 U865 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
INV_X1 U866 ( .A(n1208), .ZN(n1204) );
NAND4_X1 U867 ( .A1(n1209), .A2(n1040), .A3(n1067), .A4(n1052), .ZN(n1202) );
NOR2_X1 U868 ( .A1(KEYINPUT44), .A2(n1210), .ZN(n1186) );
XOR2_X1 U869 ( .A(n1211), .B(n1212), .Z(n1210) );
XNOR2_X1 U870 ( .A(n1213), .B(n1169), .ZN(n1212) );
NAND2_X1 U871 ( .A1(KEYINPUT47), .A2(G125), .ZN(n1211) );
XNOR2_X1 U872 ( .A(n1124), .B(KEYINPUT50), .ZN(n1183) );
NOR2_X1 U873 ( .A1(n1123), .A2(G952), .ZN(n1124) );
XOR2_X1 U874 ( .A(n1200), .B(n1214), .Z(G48) );
NOR2_X1 U875 ( .A1(G146), .A2(KEYINPUT63), .ZN(n1214) );
NAND4_X1 U876 ( .A1(n1209), .A2(n1052), .A3(n1215), .A4(n1081), .ZN(n1200) );
XNOR2_X1 U877 ( .A(G143), .B(n1201), .ZN(G45) );
NAND4_X1 U878 ( .A1(n1215), .A2(n1057), .A3(n1216), .A4(n1217), .ZN(n1201) );
AND3_X1 U879 ( .A1(n1218), .A2(n1219), .A3(n1080), .ZN(n1217) );
XOR2_X1 U880 ( .A(G140), .B(n1220), .Z(G42) );
NOR4_X1 U881 ( .A1(n1221), .A2(n1222), .A3(n1194), .A4(n1223), .ZN(n1220) );
XNOR2_X1 U882 ( .A(n1040), .B(KEYINPUT49), .ZN(n1221) );
INV_X1 U883 ( .A(n1224), .ZN(n1040) );
XOR2_X1 U884 ( .A(G137), .B(n1207), .Z(G39) );
NOR4_X1 U885 ( .A1(n1223), .A2(n1224), .A3(n1061), .A4(n1225), .ZN(n1207) );
INV_X1 U886 ( .A(n1209), .ZN(n1223) );
XOR2_X1 U887 ( .A(G134), .B(n1206), .Z(G36) );
AND2_X1 U888 ( .A1(n1226), .A2(n1051), .ZN(n1206) );
XOR2_X1 U889 ( .A(G131), .B(n1205), .Z(G33) );
AND2_X1 U890 ( .A1(n1226), .A2(n1052), .ZN(n1205) );
NOR4_X1 U891 ( .A1(n1224), .A2(n1065), .A3(n1227), .A4(n1228), .ZN(n1226) );
NAND2_X1 U892 ( .A1(n1073), .A2(n1229), .ZN(n1224) );
XNOR2_X1 U893 ( .A(G128), .B(n1208), .ZN(G30) );
NAND4_X1 U894 ( .A1(n1230), .A2(n1231), .A3(n1051), .A4(n1232), .ZN(n1208) );
NOR2_X1 U895 ( .A1(n1225), .A2(n1070), .ZN(n1232) );
OR2_X1 U896 ( .A1(n1209), .A2(KEYINPUT0), .ZN(n1231) );
NOR3_X1 U897 ( .A1(n1233), .A2(n1228), .A3(n1227), .ZN(n1209) );
NAND2_X1 U898 ( .A1(KEYINPUT0), .A2(n1234), .ZN(n1230) );
NAND3_X1 U899 ( .A1(n1219), .A2(n1227), .A3(n1068), .ZN(n1234) );
XNOR2_X1 U900 ( .A(G101), .B(n1191), .ZN(G3) );
OR3_X1 U901 ( .A1(n1065), .A2(n1029), .A3(n1061), .ZN(n1191) );
INV_X1 U902 ( .A(n1216), .ZN(n1065) );
NAND3_X1 U903 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(G27) );
NAND2_X1 U904 ( .A1(KEYINPUT40), .A2(n1100), .ZN(n1237) );
OR3_X1 U905 ( .A1(n1100), .A2(KEYINPUT40), .A3(G125), .ZN(n1236) );
NAND2_X1 U906 ( .A1(G125), .A2(n1238), .ZN(n1235) );
NAND2_X1 U907 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
INV_X1 U908 ( .A(KEYINPUT40), .ZN(n1240) );
XNOR2_X1 U909 ( .A(n1188), .B(KEYINPUT14), .ZN(n1239) );
INV_X1 U910 ( .A(n1100), .ZN(n1188) );
NAND4_X1 U911 ( .A1(n1067), .A2(n1052), .A3(n1046), .A4(n1241), .ZN(n1100) );
NOR4_X1 U912 ( .A1(n1050), .A2(n1228), .A3(n1233), .A4(n1070), .ZN(n1241) );
INV_X1 U913 ( .A(n1215), .ZN(n1070) );
INV_X1 U914 ( .A(n1219), .ZN(n1228) );
NAND2_X1 U915 ( .A1(n1058), .A2(n1242), .ZN(n1219) );
NAND4_X1 U916 ( .A1(n1104), .A2(G902), .A3(G953), .A4(n1243), .ZN(n1242) );
XNOR2_X1 U917 ( .A(G900), .B(KEYINPUT16), .ZN(n1104) );
INV_X1 U918 ( .A(n1222), .ZN(n1067) );
XOR2_X1 U919 ( .A(G122), .B(n1197), .Z(G24) );
AND4_X1 U920 ( .A1(n1244), .A2(n1047), .A3(n1218), .A4(n1080), .ZN(n1197) );
INV_X1 U921 ( .A(n1030), .ZN(n1047) );
NAND2_X1 U922 ( .A1(n1233), .A2(n1245), .ZN(n1030) );
XNOR2_X1 U923 ( .A(KEYINPUT46), .B(n1225), .ZN(n1245) );
XOR2_X1 U924 ( .A(G119), .B(n1196), .Z(G21) );
AND4_X1 U925 ( .A1(n1244), .A2(n1053), .A3(n1081), .A4(n1068), .ZN(n1196) );
XOR2_X1 U926 ( .A(G116), .B(n1195), .Z(G18) );
AND3_X1 U927 ( .A1(n1216), .A2(n1051), .A3(n1244), .ZN(n1195) );
NOR2_X1 U928 ( .A1(n1080), .A2(n1246), .ZN(n1051) );
INV_X1 U929 ( .A(n1218), .ZN(n1246) );
XOR2_X1 U930 ( .A(n1193), .B(n1247), .Z(G15) );
NAND2_X1 U931 ( .A1(KEYINPUT28), .A2(G113), .ZN(n1247) );
NAND3_X1 U932 ( .A1(n1216), .A2(n1052), .A3(n1244), .ZN(n1193) );
AND4_X1 U933 ( .A1(n1046), .A2(n1215), .A3(n1248), .A4(n1054), .ZN(n1244) );
INV_X1 U934 ( .A(n1194), .ZN(n1052) );
NAND2_X1 U935 ( .A1(n1249), .A2(n1080), .ZN(n1194) );
XNOR2_X1 U936 ( .A(n1218), .B(KEYINPUT56), .ZN(n1249) );
NOR2_X1 U937 ( .A1(n1068), .A2(n1225), .ZN(n1216) );
INV_X1 U938 ( .A(n1081), .ZN(n1225) );
XNOR2_X1 U939 ( .A(G110), .B(n1192), .ZN(G12) );
OR4_X1 U940 ( .A1(n1222), .A2(n1061), .A3(n1029), .A4(n1233), .ZN(n1192) );
INV_X1 U941 ( .A(n1068), .ZN(n1233) );
XOR2_X1 U942 ( .A(n1250), .B(n1128), .Z(n1068) );
NAND2_X1 U943 ( .A1(G217), .A2(n1251), .ZN(n1128) );
OR2_X1 U944 ( .A1(n1127), .A2(G902), .ZN(n1250) );
XNOR2_X1 U945 ( .A(n1252), .B(n1253), .ZN(n1127) );
XNOR2_X1 U946 ( .A(n1254), .B(n1255), .ZN(n1253) );
XOR2_X1 U947 ( .A(KEYINPUT10), .B(G137), .Z(n1255) );
XOR2_X1 U948 ( .A(n1256), .B(n1257), .Z(n1252) );
XOR2_X1 U949 ( .A(n1258), .B(n1259), .Z(n1256) );
NOR2_X1 U950 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U951 ( .A(KEYINPUT34), .B(G221), .Z(n1261) );
NAND3_X1 U952 ( .A1(n1262), .A2(n1248), .A3(n1215), .ZN(n1029) );
NOR2_X1 U953 ( .A1(n1073), .A2(n1072), .ZN(n1215) );
INV_X1 U954 ( .A(n1229), .ZN(n1072) );
NAND2_X1 U955 ( .A1(G214), .A2(n1263), .ZN(n1229) );
XOR2_X1 U956 ( .A(n1264), .B(n1088), .Z(n1073) );
NAND2_X1 U957 ( .A1(G210), .A2(n1263), .ZN(n1088) );
NAND2_X1 U958 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
INV_X1 U959 ( .A(G237), .ZN(n1265) );
NAND2_X1 U960 ( .A1(KEYINPUT59), .A2(n1085), .ZN(n1264) );
NAND2_X1 U961 ( .A1(n1267), .A2(n1266), .ZN(n1085) );
XOR2_X1 U962 ( .A(n1268), .B(n1121), .Z(n1267) );
XNOR2_X1 U963 ( .A(n1269), .B(n1270), .ZN(n1121) );
XOR2_X1 U964 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U965 ( .A(n1273), .B(n1257), .Z(n1269) );
XOR2_X1 U966 ( .A(G110), .B(G119), .Z(n1257) );
XNOR2_X1 U967 ( .A(n1274), .B(n1275), .ZN(n1273) );
NAND2_X1 U968 ( .A1(KEYINPUT60), .A2(G122), .ZN(n1275) );
NAND2_X1 U969 ( .A1(KEYINPUT8), .A2(n1276), .ZN(n1274) );
NAND2_X1 U970 ( .A1(n1277), .A2(n1278), .ZN(n1268) );
NAND2_X1 U971 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U972 ( .A1(KEYINPUT53), .A2(n1281), .ZN(n1280) );
NAND2_X1 U973 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U974 ( .A1(n1213), .A2(n1284), .ZN(n1277) );
NAND2_X1 U975 ( .A1(n1283), .A2(n1285), .ZN(n1284) );
NAND2_X1 U976 ( .A1(n1286), .A2(KEYINPUT53), .ZN(n1285) );
INV_X1 U977 ( .A(n1279), .ZN(n1286) );
XOR2_X1 U978 ( .A(G125), .B(n1287), .Z(n1279) );
NOR2_X1 U979 ( .A1(n1288), .A2(KEYINPUT35), .ZN(n1287) );
INV_X1 U980 ( .A(KEYINPUT11), .ZN(n1283) );
INV_X1 U981 ( .A(n1282), .ZN(n1213) );
NAND2_X1 U982 ( .A1(G224), .A2(n1289), .ZN(n1282) );
XNOR2_X1 U983 ( .A(KEYINPUT9), .B(n1123), .ZN(n1289) );
NAND2_X1 U984 ( .A1(n1058), .A2(n1290), .ZN(n1248) );
NAND4_X1 U985 ( .A1(G902), .A2(G953), .A3(n1243), .A4(n1120), .ZN(n1290) );
INV_X1 U986 ( .A(G898), .ZN(n1120) );
NAND3_X1 U987 ( .A1(n1092), .A2(n1243), .A3(n1291), .ZN(n1058) );
XNOR2_X1 U988 ( .A(G952), .B(KEYINPUT57), .ZN(n1291) );
NAND2_X1 U989 ( .A1(n1292), .A2(G234), .ZN(n1243) );
XNOR2_X1 U990 ( .A(G237), .B(KEYINPUT30), .ZN(n1292) );
XOR2_X1 U991 ( .A(G953), .B(KEYINPUT21), .Z(n1092) );
XNOR2_X1 U992 ( .A(KEYINPUT0), .B(n1227), .ZN(n1262) );
INV_X1 U993 ( .A(n1057), .ZN(n1227) );
NOR2_X1 U994 ( .A1(n1050), .A2(n1046), .ZN(n1057) );
AND3_X1 U995 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1046) );
NAND2_X1 U996 ( .A1(n1296), .A2(n1182), .ZN(n1295) );
NAND2_X1 U997 ( .A1(n1297), .A2(n1298), .ZN(n1294) );
INV_X1 U998 ( .A(KEYINPUT62), .ZN(n1298) );
NAND2_X1 U999 ( .A1(n1299), .A2(n1083), .ZN(n1297) );
XNOR2_X1 U1000 ( .A(KEYINPUT23), .B(n1182), .ZN(n1299) );
NAND2_X1 U1001 ( .A1(KEYINPUT62), .A2(n1300), .ZN(n1293) );
NAND2_X1 U1002 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1003 ( .A1(KEYINPUT23), .A2(n1182), .ZN(n1302) );
OR3_X1 U1004 ( .A1(n1296), .A2(KEYINPUT23), .A3(n1182), .ZN(n1301) );
INV_X1 U1005 ( .A(G469), .ZN(n1182) );
INV_X1 U1006 ( .A(n1083), .ZN(n1296) );
NAND2_X1 U1007 ( .A1(n1303), .A2(n1266), .ZN(n1083) );
XNOR2_X1 U1008 ( .A(n1178), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1009 ( .A(n1305), .B(n1306), .ZN(n1304) );
NOR2_X1 U1010 ( .A1(KEYINPUT1), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1011 ( .A(n1180), .B(n1308), .Z(n1307) );
NAND2_X1 U1012 ( .A1(n1309), .A2(n1177), .ZN(n1308) );
XOR2_X1 U1013 ( .A(G110), .B(G140), .Z(n1177) );
XNOR2_X1 U1014 ( .A(KEYINPUT37), .B(KEYINPUT26), .ZN(n1309) );
NAND2_X1 U1015 ( .A1(G227), .A2(n1123), .ZN(n1180) );
NOR2_X1 U1016 ( .A1(KEYINPUT24), .A2(n1107), .ZN(n1305) );
XNOR2_X1 U1017 ( .A(G128), .B(n1310), .ZN(n1107) );
NOR2_X1 U1018 ( .A1(KEYINPUT41), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1019 ( .A(n1312), .B(n1171), .Z(n1178) );
INV_X1 U1020 ( .A(n1170), .ZN(n1171) );
NAND2_X1 U1021 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
OR2_X1 U1022 ( .A1(n1315), .A2(G101), .ZN(n1314) );
XOR2_X1 U1023 ( .A(n1316), .B(KEYINPUT61), .Z(n1313) );
NAND2_X1 U1024 ( .A1(G101), .A2(n1315), .ZN(n1316) );
XNOR2_X1 U1025 ( .A(G104), .B(n1317), .ZN(n1315) );
INV_X1 U1026 ( .A(n1054), .ZN(n1050) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1251), .ZN(n1054) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1266), .ZN(n1251) );
INV_X1 U1029 ( .A(n1053), .ZN(n1061) );
NOR2_X1 U1030 ( .A1(n1218), .A2(n1080), .ZN(n1053) );
XOR2_X1 U1031 ( .A(n1318), .B(n1140), .Z(n1080) );
INV_X1 U1032 ( .A(G475), .ZN(n1140) );
NAND2_X1 U1033 ( .A1(n1138), .A2(n1266), .ZN(n1318) );
INV_X1 U1034 ( .A(G902), .ZN(n1266) );
XNOR2_X1 U1035 ( .A(n1319), .B(n1320), .ZN(n1138) );
XOR2_X1 U1036 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1037 ( .A(G122), .B(KEYINPUT20), .ZN(n1322) );
NAND2_X1 U1038 ( .A1(KEYINPUT4), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1039 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1040 ( .A(G131), .B(n1326), .ZN(n1325) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1327), .ZN(n1326) );
NOR2_X1 U1042 ( .A1(KEYINPUT19), .A2(n1328), .ZN(n1324) );
XOR2_X1 U1043 ( .A(n1258), .B(n1271), .Z(n1319) );
XNOR2_X1 U1044 ( .A(n1329), .B(G113), .ZN(n1271) );
INV_X1 U1045 ( .A(G104), .ZN(n1329) );
XOR2_X1 U1046 ( .A(G146), .B(n1110), .Z(n1258) );
XNOR2_X1 U1047 ( .A(G140), .B(G125), .ZN(n1110) );
XOR2_X1 U1048 ( .A(n1330), .B(n1089), .Z(n1218) );
INV_X1 U1049 ( .A(G478), .ZN(n1089) );
NAND2_X1 U1050 ( .A1(KEYINPUT5), .A2(n1091), .ZN(n1330) );
NOR2_X1 U1051 ( .A1(n1134), .A2(G902), .ZN(n1091) );
XNOR2_X1 U1052 ( .A(n1331), .B(n1332), .ZN(n1134) );
NOR2_X1 U1053 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XOR2_X1 U1054 ( .A(n1335), .B(KEYINPUT2), .Z(n1334) );
NAND2_X1 U1055 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
NOR2_X1 U1056 ( .A1(n1336), .A2(n1337), .ZN(n1333) );
XNOR2_X1 U1057 ( .A(n1254), .B(n1338), .ZN(n1337) );
XNOR2_X1 U1058 ( .A(n1328), .B(G134), .ZN(n1338) );
INV_X1 U1059 ( .A(G143), .ZN(n1328) );
XNOR2_X1 U1060 ( .A(G122), .B(n1272), .ZN(n1336) );
XNOR2_X1 U1061 ( .A(n1317), .B(G116), .ZN(n1272) );
INV_X1 U1062 ( .A(G107), .ZN(n1317) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1339), .ZN(n1331) );
INV_X1 U1064 ( .A(n1260), .ZN(n1339) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1123), .ZN(n1260) );
INV_X1 U1066 ( .A(G953), .ZN(n1123) );
XOR2_X1 U1067 ( .A(n1081), .B(KEYINPUT51), .Z(n1222) );
XOR2_X1 U1068 ( .A(n1340), .B(n1155), .Z(n1081) );
INV_X1 U1069 ( .A(G472), .ZN(n1155) );
NAND2_X1 U1070 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1071 ( .A(n1343), .B(n1146), .ZN(n1342) );
AND2_X1 U1072 ( .A1(n1344), .A2(n1345), .ZN(n1146) );
NAND2_X1 U1073 ( .A1(n1346), .A2(n1276), .ZN(n1345) );
INV_X1 U1074 ( .A(G101), .ZN(n1276) );
NAND2_X1 U1075 ( .A1(G210), .A2(n1327), .ZN(n1346) );
NAND3_X1 U1076 ( .A1(G210), .A2(n1327), .A3(G101), .ZN(n1344) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1327) );
NAND2_X1 U1078 ( .A1(n1347), .A2(n1348), .ZN(n1343) );
NAND2_X1 U1079 ( .A1(n1349), .A2(n1161), .ZN(n1348) );
XOR2_X1 U1080 ( .A(KEYINPUT31), .B(n1350), .Z(n1347) );
NOR2_X1 U1081 ( .A1(n1161), .A2(n1349), .ZN(n1350) );
XNOR2_X1 U1082 ( .A(n1288), .B(n1170), .ZN(n1349) );
XNOR2_X1 U1083 ( .A(n1351), .B(n1352), .ZN(n1170) );
NOR2_X1 U1084 ( .A1(G137), .A2(KEYINPUT27), .ZN(n1352) );
XNOR2_X1 U1085 ( .A(G131), .B(G134), .ZN(n1351) );
INV_X1 U1086 ( .A(n1169), .ZN(n1288) );
NAND2_X1 U1087 ( .A1(n1353), .A2(n1354), .ZN(n1169) );
NAND2_X1 U1088 ( .A1(n1311), .A2(n1355), .ZN(n1354) );
XOR2_X1 U1089 ( .A(KEYINPUT17), .B(n1356), .Z(n1353) );
NOR2_X1 U1090 ( .A1(n1311), .A2(n1355), .ZN(n1356) );
XNOR2_X1 U1091 ( .A(KEYINPUT45), .B(n1254), .ZN(n1355) );
INV_X1 U1092 ( .A(G128), .ZN(n1254) );
XNOR2_X1 U1093 ( .A(G146), .B(G143), .ZN(n1311) );
INV_X1 U1094 ( .A(n1162), .ZN(n1161) );
XNOR2_X1 U1095 ( .A(n1357), .B(n1358), .ZN(n1162) );
NOR2_X1 U1096 ( .A1(KEYINPUT42), .A2(n1359), .ZN(n1358) );
XNOR2_X1 U1097 ( .A(G119), .B(KEYINPUT32), .ZN(n1359) );
XNOR2_X1 U1098 ( .A(G113), .B(G116), .ZN(n1357) );
XNOR2_X1 U1099 ( .A(G902), .B(KEYINPUT48), .ZN(n1341) );
endmodule


