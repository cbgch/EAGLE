//Key = 0010111101111010101110010000010110010100100000110100111100000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;

XNOR2_X1 U716 ( .A(G107), .B(n990), .ZN(G9) );
NOR2_X1 U717 ( .A1(n991), .A2(n992), .ZN(G75) );
NOR4_X1 U718 ( .A1(G953), .A2(n993), .A3(n994), .A4(n995), .ZN(n992) );
NOR2_X1 U719 ( .A1(n996), .A2(n997), .ZN(n994) );
NOR2_X1 U720 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR3_X1 U721 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n999) );
NOR4_X1 U722 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NOR3_X1 U723 ( .A1(n1007), .A2(KEYINPUT26), .A3(n1008), .ZN(n1006) );
NOR2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1004) );
NOR2_X1 U725 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U726 ( .A1(n1013), .A2(n1014), .ZN(n1001) );
NOR3_X1 U727 ( .A1(n1015), .A2(n1008), .A3(n1007), .ZN(n1014) );
XOR2_X1 U728 ( .A(n1016), .B(KEYINPUT5), .Z(n1007) );
INV_X1 U729 ( .A(KEYINPUT26), .ZN(n1015) );
NOR3_X1 U730 ( .A1(n1008), .A2(n1017), .A3(n1010), .ZN(n998) );
INV_X1 U731 ( .A(n1018), .ZN(n1010) );
NOR2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U733 ( .A1(n1021), .A2(n1000), .ZN(n1020) );
INV_X1 U734 ( .A(n1022), .ZN(n1000) );
NOR2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U737 ( .A1(n1027), .A2(n1003), .ZN(n1019) );
NOR2_X1 U738 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
INV_X1 U740 ( .A(n1032), .ZN(n1008) );
NOR3_X1 U741 ( .A1(n993), .A2(G953), .A3(G952), .ZN(n991) );
AND4_X1 U742 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n993) );
NOR4_X1 U743 ( .A1(n1037), .A2(n1025), .A3(n1038), .A4(n1039), .ZN(n1036) );
XOR2_X1 U744 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U745 ( .A1(G475), .A2(KEYINPUT41), .ZN(n1041) );
XNOR2_X1 U746 ( .A(n1042), .B(KEYINPUT9), .ZN(n1038) );
NAND3_X1 U747 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1037) );
XOR2_X1 U748 ( .A(n1046), .B(KEYINPUT21), .Z(n1045) );
NAND2_X1 U749 ( .A1(G478), .A2(n1047), .ZN(n1046) );
NAND2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NAND2_X1 U751 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U752 ( .A1(KEYINPUT57), .A2(n1052), .ZN(n1051) );
NAND2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
INV_X1 U754 ( .A(KEYINPUT57), .ZN(n1054) );
OR2_X1 U755 ( .A1(n1053), .A2(n1049), .ZN(n1043) );
NAND2_X1 U756 ( .A1(KEYINPUT37), .A2(n1052), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1035) );
NOR2_X1 U758 ( .A1(G478), .A2(n1047), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1033) );
XOR2_X1 U760 ( .A(n1060), .B(n1061), .Z(G72) );
NOR2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND3_X1 U763 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1060) );
NAND3_X1 U764 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
INV_X1 U765 ( .A(n1072), .ZN(n1071) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1063), .ZN(n1070) );
NAND2_X1 U767 ( .A1(G953), .A2(n1065), .ZN(n1069) );
NAND3_X1 U768 ( .A1(KEYINPUT12), .A2(n1072), .A3(n1074), .ZN(n1067) );
XNOR2_X1 U769 ( .A(n1075), .B(n1076), .ZN(n1072) );
XNOR2_X1 U770 ( .A(KEYINPUT35), .B(n1077), .ZN(n1075) );
NOR2_X1 U771 ( .A1(KEYINPUT1), .A2(n1078), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(n1078) );
XOR2_X1 U773 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U774 ( .A1(G134), .A2(KEYINPUT34), .ZN(n1081) );
OR2_X1 U775 ( .A1(n1074), .A2(KEYINPUT12), .ZN(n1066) );
AND2_X1 U776 ( .A1(n1063), .A2(n1073), .ZN(n1074) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(G69) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U779 ( .A1(G953), .A2(n1087), .ZN(n1086) );
NAND3_X1 U780 ( .A1(G953), .A2(n1088), .A3(n1089), .ZN(n1083) );
INV_X1 U781 ( .A(n1085), .ZN(n1089) );
XNOR2_X1 U782 ( .A(n1090), .B(n1091), .ZN(n1085) );
NOR2_X1 U783 ( .A1(n1092), .A2(G953), .ZN(n1091) );
NOR2_X1 U784 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U786 ( .A1(G953), .A2(n1097), .ZN(n1096) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1095) );
NAND2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U790 ( .A(n1104), .B(KEYINPUT15), .Z(n1102) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
XOR2_X1 U792 ( .A(n1104), .B(KEYINPUT47), .Z(n1106) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1088) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U795 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U796 ( .A(n1111), .B(KEYINPUT24), .Z(n1110) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1107), .A2(n1114), .ZN(G63) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U800 ( .A1(n1112), .A2(G478), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1117), .A2(KEYINPUT62), .ZN(n1115) );
XOR2_X1 U802 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(G60) );
AND2_X1 U804 ( .A1(KEYINPUT6), .A2(n1107), .ZN(n1122) );
NOR3_X1 U805 ( .A1(KEYINPUT6), .A2(G953), .A3(G952), .ZN(n1121) );
XOR2_X1 U806 ( .A(n1123), .B(n1124), .Z(n1120) );
NAND2_X1 U807 ( .A1(n1112), .A2(G475), .ZN(n1123) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(G6) );
NAND2_X1 U809 ( .A1(n1127), .A2(KEYINPUT52), .ZN(n1126) );
XNOR2_X1 U810 ( .A(G104), .B(KEYINPUT61), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1024), .A2(n1128), .ZN(n1125) );
XNOR2_X1 U812 ( .A(KEYINPUT48), .B(n1129), .ZN(n1128) );
NOR2_X1 U813 ( .A1(n1107), .A2(n1130), .ZN(G57) );
XOR2_X1 U814 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U815 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U816 ( .A1(n1112), .A2(G472), .ZN(n1134) );
NAND2_X1 U817 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
OR2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U819 ( .A(n1139), .B(KEYINPUT17), .Z(n1135) );
NAND2_X1 U820 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
XOR2_X1 U821 ( .A(G101), .B(KEYINPUT46), .Z(n1138) );
XNOR2_X1 U822 ( .A(n1140), .B(n1141), .ZN(n1131) );
NOR2_X1 U823 ( .A1(n1107), .A2(n1142), .ZN(G54) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U825 ( .A(n1145), .B(n1079), .Z(n1144) );
XOR2_X1 U826 ( .A(n1146), .B(n1147), .Z(n1143) );
NOR3_X1 U827 ( .A1(n1064), .A2(KEYINPUT0), .A3(G953), .ZN(n1147) );
NAND2_X1 U828 ( .A1(n1112), .A2(G469), .ZN(n1146) );
NOR2_X1 U829 ( .A1(n1107), .A2(n1148), .ZN(G51) );
XOR2_X1 U830 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U831 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U832 ( .A1(n1112), .A2(n1153), .ZN(n1151) );
XOR2_X1 U833 ( .A(KEYINPUT13), .B(n1154), .Z(n1153) );
AND2_X1 U834 ( .A1(G902), .A2(n995), .ZN(n1112) );
OR3_X1 U835 ( .A1(n1094), .A2(n1155), .A3(n1073), .ZN(n995) );
NAND2_X1 U836 ( .A1(n1156), .A2(n1157), .ZN(n1073) );
NOR4_X1 U837 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1157) );
NOR4_X1 U838 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1156) );
INV_X1 U839 ( .A(n1166), .ZN(n1164) );
XOR2_X1 U840 ( .A(KEYINPUT3), .B(n1093), .Z(n1155) );
NAND4_X1 U841 ( .A1(n1167), .A2(n1168), .A3(n990), .A4(n1169), .ZN(n1093) );
NAND4_X1 U842 ( .A1(n1170), .A2(n1029), .A3(n1011), .A4(n1018), .ZN(n990) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1024), .ZN(n1167) );
XOR2_X1 U844 ( .A(n1129), .B(KEYINPUT14), .Z(n1171) );
NAND4_X1 U845 ( .A1(n1012), .A2(n1029), .A3(n1018), .A4(n1172), .ZN(n1129) );
NAND4_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1094) );
NAND4_X1 U847 ( .A1(n1177), .A2(n1016), .A3(n1012), .A4(n1170), .ZN(n1173) );
XNOR2_X1 U848 ( .A(n1022), .B(KEYINPUT16), .ZN(n1177) );
XOR2_X1 U849 ( .A(G125), .B(n1178), .Z(n1149) );
NOR2_X1 U850 ( .A1(n1063), .A2(G952), .ZN(n1107) );
NAND2_X1 U851 ( .A1(n1179), .A2(n1180), .ZN(G48) );
NAND2_X1 U852 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U853 ( .A1(n1165), .A2(n1183), .ZN(n1182) );
OR2_X1 U854 ( .A1(KEYINPUT2), .A2(KEYINPUT25), .ZN(n1183) );
NAND3_X1 U855 ( .A1(KEYINPUT2), .A2(n1184), .A3(n1185), .ZN(n1179) );
INV_X1 U856 ( .A(n1181), .ZN(n1185) );
XOR2_X1 U857 ( .A(G146), .B(KEYINPUT51), .Z(n1181) );
XOR2_X1 U858 ( .A(KEYINPUT25), .B(n1165), .Z(n1184) );
AND3_X1 U859 ( .A1(n1186), .A2(n1024), .A3(n1012), .ZN(n1165) );
XNOR2_X1 U860 ( .A(G143), .B(n1166), .ZN(G45) );
NAND3_X1 U861 ( .A1(n1187), .A2(n1024), .A3(n1188), .ZN(n1166) );
XOR2_X1 U862 ( .A(G140), .B(n1163), .Z(G42) );
AND3_X1 U863 ( .A1(n1013), .A2(n1029), .A3(n1189), .ZN(n1163) );
XOR2_X1 U864 ( .A(G137), .B(n1158), .Z(G39) );
AND3_X1 U865 ( .A1(n1186), .A2(n1013), .A3(n1032), .ZN(n1158) );
XOR2_X1 U866 ( .A(G134), .B(n1162), .Z(G36) );
AND3_X1 U867 ( .A1(n1013), .A2(n1011), .A3(n1187), .ZN(n1162) );
XNOR2_X1 U868 ( .A(n1161), .B(n1190), .ZN(G33) );
XNOR2_X1 U869 ( .A(KEYINPUT40), .B(n1191), .ZN(n1190) );
AND3_X1 U870 ( .A1(n1012), .A2(n1013), .A3(n1187), .ZN(n1161) );
AND3_X1 U871 ( .A1(n1029), .A2(n1192), .A3(n1016), .ZN(n1187) );
INV_X1 U872 ( .A(n1003), .ZN(n1013) );
NAND2_X1 U873 ( .A1(n1193), .A2(n1194), .ZN(n1003) );
XNOR2_X1 U874 ( .A(KEYINPUT4), .B(n1026), .ZN(n1194) );
XOR2_X1 U875 ( .A(G128), .B(n1160), .Z(G30) );
AND3_X1 U876 ( .A1(n1011), .A2(n1024), .A3(n1186), .ZN(n1160) );
AND4_X1 U877 ( .A1(n1029), .A2(n1042), .A3(n1192), .A4(n1195), .ZN(n1186) );
XNOR2_X1 U878 ( .A(n1168), .B(n1196), .ZN(G3) );
NOR2_X1 U879 ( .A1(KEYINPUT33), .A2(n1197), .ZN(n1196) );
NAND4_X1 U880 ( .A1(n1016), .A2(n1032), .A3(n1170), .A4(n1029), .ZN(n1168) );
XOR2_X1 U881 ( .A(G125), .B(n1159), .Z(G27) );
AND3_X1 U882 ( .A1(n1189), .A2(n1024), .A3(n1022), .ZN(n1159) );
AND4_X1 U883 ( .A1(n1198), .A2(n1012), .A3(n1192), .A4(n1195), .ZN(n1189) );
NAND2_X1 U884 ( .A1(n997), .A2(n1199), .ZN(n1192) );
NAND4_X1 U885 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1065), .ZN(n1199) );
INV_X1 U886 ( .A(G900), .ZN(n1065) );
XNOR2_X1 U887 ( .A(G122), .B(n1174), .ZN(G24) );
NAND3_X1 U888 ( .A1(n1188), .A2(n1018), .A3(n1201), .ZN(n1174) );
NOR2_X1 U889 ( .A1(n1195), .A2(n1042), .ZN(n1018) );
AND2_X1 U890 ( .A1(n1202), .A2(n1203), .ZN(n1188) );
XNOR2_X1 U891 ( .A(KEYINPUT58), .B(n1204), .ZN(n1202) );
XOR2_X1 U892 ( .A(n1175), .B(n1205), .Z(G21) );
NAND2_X1 U893 ( .A1(KEYINPUT29), .A2(G119), .ZN(n1205) );
NAND4_X1 U894 ( .A1(n1201), .A2(n1032), .A3(n1042), .A4(n1195), .ZN(n1175) );
XNOR2_X1 U895 ( .A(G116), .B(n1176), .ZN(G18) );
NAND2_X1 U896 ( .A1(n1206), .A2(n1011), .ZN(n1176) );
NOR2_X1 U897 ( .A1(n1203), .A2(n1204), .ZN(n1011) );
XNOR2_X1 U898 ( .A(G113), .B(n1207), .ZN(G15) );
NAND2_X1 U899 ( .A1(n1206), .A2(n1012), .ZN(n1207) );
AND2_X1 U900 ( .A1(n1204), .A2(n1203), .ZN(n1012) );
INV_X1 U901 ( .A(n1208), .ZN(n1204) );
AND2_X1 U902 ( .A1(n1201), .A2(n1016), .ZN(n1206) );
NOR2_X1 U903 ( .A1(n1195), .A2(n1198), .ZN(n1016) );
AND2_X1 U904 ( .A1(n1022), .A2(n1170), .ZN(n1201) );
NOR2_X1 U905 ( .A1(n1030), .A2(n1055), .ZN(n1022) );
XOR2_X1 U906 ( .A(G110), .B(n1209), .Z(G12) );
NOR2_X1 U907 ( .A1(n1210), .A2(n1169), .ZN(n1209) );
NAND3_X1 U908 ( .A1(n1170), .A2(n1029), .A3(n1005), .ZN(n1169) );
AND3_X1 U909 ( .A1(n1198), .A2(n1195), .A3(n1032), .ZN(n1005) );
NOR2_X1 U910 ( .A1(n1208), .A2(n1203), .ZN(n1032) );
XNOR2_X1 U911 ( .A(n1040), .B(G475), .ZN(n1203) );
NAND2_X1 U912 ( .A1(n1124), .A2(n1211), .ZN(n1040) );
XOR2_X1 U913 ( .A(n1212), .B(n1213), .Z(n1124) );
XNOR2_X1 U914 ( .A(n1076), .B(n1214), .ZN(n1213) );
XOR2_X1 U915 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U916 ( .A1(KEYINPUT8), .A2(n1217), .ZN(n1216) );
XOR2_X1 U917 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U918 ( .A(G113), .B(G104), .Z(n1219) );
XNOR2_X1 U919 ( .A(KEYINPUT43), .B(n1220), .ZN(n1218) );
INV_X1 U920 ( .A(G122), .ZN(n1220) );
NAND2_X1 U921 ( .A1(n1221), .A2(G214), .ZN(n1215) );
XOR2_X1 U922 ( .A(G125), .B(G140), .Z(n1076) );
XOR2_X1 U923 ( .A(n1222), .B(n1223), .Z(n1212) );
XNOR2_X1 U924 ( .A(KEYINPUT22), .B(n1224), .ZN(n1223) );
INV_X1 U925 ( .A(G146), .ZN(n1224) );
XNOR2_X1 U926 ( .A(G131), .B(G143), .ZN(n1222) );
XOR2_X1 U927 ( .A(G478), .B(n1225), .Z(n1208) );
NOR2_X1 U928 ( .A1(KEYINPUT39), .A2(n1047), .ZN(n1225) );
NAND2_X1 U929 ( .A1(n1226), .A2(n1211), .ZN(n1047) );
XNOR2_X1 U930 ( .A(n1119), .B(n1118), .ZN(n1226) );
XOR2_X1 U931 ( .A(n1227), .B(n1228), .Z(n1118) );
XNOR2_X1 U932 ( .A(n1229), .B(G107), .ZN(n1228) );
NAND2_X1 U933 ( .A1(G217), .A2(n1230), .ZN(n1227) );
XNOR2_X1 U934 ( .A(n1231), .B(n1232), .ZN(n1119) );
XNOR2_X1 U935 ( .A(n1233), .B(G134), .ZN(n1232) );
XNOR2_X1 U936 ( .A(G128), .B(G122), .ZN(n1231) );
NAND3_X1 U937 ( .A1(n1234), .A2(n1235), .A3(n1034), .ZN(n1195) );
NAND2_X1 U938 ( .A1(n1113), .A2(n1236), .ZN(n1034) );
INV_X1 U939 ( .A(n1059), .ZN(n1113) );
OR2_X1 U940 ( .A1(n1058), .A2(KEYINPUT31), .ZN(n1235) );
NAND3_X1 U941 ( .A1(n1058), .A2(n1059), .A3(KEYINPUT31), .ZN(n1234) );
NAND2_X1 U942 ( .A1(G217), .A2(n1237), .ZN(n1059) );
INV_X1 U943 ( .A(n1236), .ZN(n1058) );
NAND2_X1 U944 ( .A1(n1109), .A2(n1211), .ZN(n1236) );
XOR2_X1 U945 ( .A(n1238), .B(n1239), .Z(n1109) );
XOR2_X1 U946 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U947 ( .A(G119), .B(G110), .Z(n1241) );
XOR2_X1 U948 ( .A(KEYINPUT60), .B(G137), .Z(n1240) );
XOR2_X1 U949 ( .A(n1242), .B(n1243), .Z(n1238) );
XOR2_X1 U950 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U951 ( .A1(n1230), .A2(G221), .ZN(n1245) );
AND2_X1 U952 ( .A1(G234), .A2(n1063), .ZN(n1230) );
NAND2_X1 U953 ( .A1(n1246), .A2(KEYINPUT18), .ZN(n1244) );
XOR2_X1 U954 ( .A(n1247), .B(G140), .Z(n1246) );
NAND2_X1 U955 ( .A1(KEYINPUT49), .A2(G125), .ZN(n1247) );
INV_X1 U956 ( .A(n1042), .ZN(n1198) );
XNOR2_X1 U957 ( .A(n1248), .B(G472), .ZN(n1042) );
NAND2_X1 U958 ( .A1(n1249), .A2(n1211), .ZN(n1248) );
XOR2_X1 U959 ( .A(n1250), .B(n1251), .Z(n1249) );
XNOR2_X1 U960 ( .A(n1197), .B(n1252), .ZN(n1251) );
NOR2_X1 U961 ( .A1(KEYINPUT36), .A2(n1253), .ZN(n1252) );
INV_X1 U962 ( .A(n1137), .ZN(n1253) );
NAND2_X1 U963 ( .A1(n1221), .A2(G210), .ZN(n1137) );
NOR2_X1 U964 ( .A1(G953), .A2(G237), .ZN(n1221) );
NAND2_X1 U965 ( .A1(n1254), .A2(n1255), .ZN(n1250) );
OR2_X1 U966 ( .A1(n1141), .A2(n1140), .ZN(n1255) );
XOR2_X1 U967 ( .A(n1256), .B(KEYINPUT56), .Z(n1254) );
NAND2_X1 U968 ( .A1(n1140), .A2(n1141), .ZN(n1256) );
XNOR2_X1 U969 ( .A(n1257), .B(n1258), .ZN(n1141) );
XOR2_X1 U970 ( .A(G119), .B(n1259), .Z(n1258) );
NOR2_X1 U971 ( .A1(KEYINPUT38), .A2(n1260), .ZN(n1259) );
NAND2_X1 U972 ( .A1(KEYINPUT23), .A2(n1229), .ZN(n1257) );
XOR2_X1 U973 ( .A(n1261), .B(n1262), .Z(n1140) );
NOR2_X1 U974 ( .A1(n1263), .A2(n1055), .ZN(n1029) );
INV_X1 U975 ( .A(n1031), .ZN(n1055) );
NAND2_X1 U976 ( .A1(G221), .A2(n1237), .ZN(n1031) );
NAND2_X1 U977 ( .A1(G234), .A2(n1211), .ZN(n1237) );
INV_X1 U978 ( .A(n1030), .ZN(n1263) );
XOR2_X1 U979 ( .A(n1052), .B(n1049), .Z(n1030) );
INV_X1 U980 ( .A(G469), .ZN(n1049) );
NAND2_X1 U981 ( .A1(n1264), .A2(n1211), .ZN(n1052) );
XOR2_X1 U982 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U983 ( .A(KEYINPUT20), .B(n1064), .ZN(n1266) );
INV_X1 U984 ( .A(G227), .ZN(n1064) );
XOR2_X1 U985 ( .A(n1145), .B(n1267), .Z(n1265) );
NOR2_X1 U986 ( .A1(KEYINPUT42), .A2(n1079), .ZN(n1267) );
NAND2_X1 U987 ( .A1(n1268), .A2(n1269), .ZN(n1079) );
NAND2_X1 U988 ( .A1(n1270), .A2(n1233), .ZN(n1269) );
INV_X1 U989 ( .A(G143), .ZN(n1233) );
XOR2_X1 U990 ( .A(KEYINPUT32), .B(n1271), .Z(n1270) );
NAND2_X1 U991 ( .A1(G143), .A2(n1272), .ZN(n1268) );
XNOR2_X1 U992 ( .A(n1271), .B(KEYINPUT55), .ZN(n1272) );
XOR2_X1 U993 ( .A(n1273), .B(n1274), .Z(n1145) );
XOR2_X1 U994 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U995 ( .A(G140), .B(G110), .Z(n1276) );
XOR2_X1 U996 ( .A(KEYINPUT59), .B(KEYINPUT45), .Z(n1275) );
XOR2_X1 U997 ( .A(n1277), .B(n1278), .Z(n1273) );
XNOR2_X1 U998 ( .A(n1262), .B(G107), .ZN(n1277) );
XOR2_X1 U999 ( .A(G134), .B(n1082), .Z(n1262) );
XNOR2_X1 U1000 ( .A(n1191), .B(G137), .ZN(n1082) );
INV_X1 U1001 ( .A(G131), .ZN(n1191) );
AND2_X1 U1002 ( .A1(n1024), .A2(n1172), .ZN(n1170) );
NAND2_X1 U1003 ( .A1(n997), .A2(n1279), .ZN(n1172) );
NAND4_X1 U1004 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1097), .ZN(n1279) );
INV_X1 U1005 ( .A(G898), .ZN(n1097) );
NAND3_X1 U1006 ( .A1(n1200), .A2(n1063), .A3(G952), .ZN(n997) );
INV_X1 U1007 ( .A(G953), .ZN(n1063) );
NAND2_X1 U1008 ( .A1(G237), .A2(G234), .ZN(n1200) );
NOR2_X1 U1009 ( .A1(n1193), .A2(n1056), .ZN(n1024) );
INV_X1 U1010 ( .A(n1026), .ZN(n1056) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1280), .ZN(n1026) );
INV_X1 U1012 ( .A(n1025), .ZN(n1193) );
XNOR2_X1 U1013 ( .A(n1281), .B(n1154), .ZN(n1025) );
AND2_X1 U1014 ( .A1(G210), .A2(n1280), .ZN(n1154) );
NAND2_X1 U1015 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
INV_X1 U1016 ( .A(G237), .ZN(n1283) );
XNOR2_X1 U1017 ( .A(KEYINPUT7), .B(n1211), .ZN(n1282) );
NAND2_X1 U1018 ( .A1(n1284), .A2(n1211), .ZN(n1281) );
INV_X1 U1019 ( .A(G902), .ZN(n1211) );
XOR2_X1 U1020 ( .A(n1152), .B(n1285), .Z(n1284) );
XOR2_X1 U1021 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U1022 ( .A1(KEYINPUT27), .A2(G125), .ZN(n1287) );
NAND2_X1 U1023 ( .A1(KEYINPUT63), .A2(n1178), .ZN(n1286) );
NOR2_X1 U1024 ( .A1(n1087), .A2(G953), .ZN(n1178) );
INV_X1 U1025 ( .A(G224), .ZN(n1087) );
XOR2_X1 U1026 ( .A(n1288), .B(n1289), .Z(n1152) );
XOR2_X1 U1027 ( .A(n1290), .B(n1104), .Z(n1289) );
NAND2_X1 U1028 ( .A1(n1291), .A2(n1292), .ZN(n1104) );
OR2_X1 U1029 ( .A1(n1293), .A2(n1260), .ZN(n1292) );
XOR2_X1 U1030 ( .A(n1294), .B(KEYINPUT50), .Z(n1291) );
NAND2_X1 U1031 ( .A1(n1260), .A2(n1293), .ZN(n1294) );
NAND2_X1 U1032 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
NAND2_X1 U1033 ( .A1(G119), .A2(n1229), .ZN(n1296) );
XOR2_X1 U1034 ( .A(n1297), .B(KEYINPUT30), .Z(n1295) );
OR2_X1 U1035 ( .A1(n1229), .A2(G119), .ZN(n1297) );
INV_X1 U1036 ( .A(G116), .ZN(n1229) );
XNOR2_X1 U1037 ( .A(G113), .B(KEYINPUT10), .ZN(n1260) );
NAND2_X1 U1038 ( .A1(KEYINPUT53), .A2(n1103), .ZN(n1290) );
INV_X1 U1039 ( .A(n1105), .ZN(n1103) );
XNOR2_X1 U1040 ( .A(n1298), .B(n1278), .ZN(n1105) );
XNOR2_X1 U1041 ( .A(G104), .B(n1197), .ZN(n1278) );
INV_X1 U1042 ( .A(G101), .ZN(n1197) );
NAND2_X1 U1043 ( .A1(KEYINPUT19), .A2(n1299), .ZN(n1298) );
INV_X1 U1044 ( .A(G107), .ZN(n1299) );
XOR2_X1 U1045 ( .A(n1300), .B(n1261), .Z(n1288) );
XOR2_X1 U1046 ( .A(G143), .B(n1271), .Z(n1261) );
XNOR2_X1 U1047 ( .A(n1242), .B(KEYINPUT28), .ZN(n1271) );
XNOR2_X1 U1048 ( .A(G128), .B(G146), .ZN(n1242) );
NAND2_X1 U1049 ( .A1(KEYINPUT11), .A2(n1099), .ZN(n1300) );
XNOR2_X1 U1050 ( .A(G110), .B(G122), .ZN(n1099) );
XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(KEYINPUT44), .ZN(n1210) );
endmodule


