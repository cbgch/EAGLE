//Key = 1110100101100010111000000110011000101110010111101001100100110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339;

XNOR2_X1 U739 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U740 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U741 ( .A1(G953), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
NOR2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U746 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR3_X1 U753 ( .A1(n1043), .A2(n1046), .A3(n1037), .ZN(n1030) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR4_X1 U756 ( .A1(n1051), .A2(n1037), .A3(n1033), .A4(n1043), .ZN(n1026) );
NOR2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR3_X1 U758 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U759 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1021) );
NOR4_X1 U760 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
XNOR2_X1 U761 ( .A(KEYINPUT4), .B(n1062), .ZN(n1061) );
NOR3_X1 U762 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1056) );
NAND2_X1 U763 ( .A1(G469), .A2(n1066), .ZN(n1055) );
XOR2_X1 U764 ( .A(n1067), .B(n1068), .Z(G72) );
NOR2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U768 ( .A1(G227), .A2(n1075), .ZN(n1073) );
XNOR2_X1 U769 ( .A(n1076), .B(n1077), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1069) );
XNOR2_X1 U771 ( .A(n1077), .B(n1080), .ZN(n1079) );
INV_X1 U772 ( .A(n1076), .ZN(n1080) );
XNOR2_X1 U773 ( .A(n1081), .B(n1082), .ZN(n1076) );
NAND2_X1 U774 ( .A1(KEYINPUT7), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U775 ( .A(n1084), .B(n1085), .ZN(n1077) );
NOR2_X1 U776 ( .A1(n1086), .A2(KEYINPUT24), .ZN(n1085) );
XNOR2_X1 U777 ( .A(G134), .B(G137), .ZN(n1084) );
NOR2_X1 U778 ( .A1(G227), .A2(n1072), .ZN(n1078) );
NAND2_X1 U779 ( .A1(n1072), .A2(n1087), .ZN(n1067) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U781 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(G69) );
INV_X1 U782 ( .A(n1093), .ZN(n1092) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1072), .ZN(n1091) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1100), .B(KEYINPUT50), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1101), .A2(G953), .ZN(n1090) );
XOR2_X1 U788 ( .A(n1095), .B(G224), .Z(n1101) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U791 ( .A(n1106), .B(KEYINPUT9), .ZN(n1104) );
INV_X1 U792 ( .A(n1107), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XNOR2_X1 U794 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1114), .ZN(G63) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U798 ( .A1(KEYINPUT42), .A2(n1117), .ZN(n1116) );
INV_X1 U799 ( .A(n1118), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1119), .A2(G478), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1108), .A2(n1120), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1121), .B(n1122), .ZN(n1120) );
AND2_X1 U803 ( .A1(G475), .A2(n1119), .ZN(n1121) );
XNOR2_X1 U804 ( .A(G104), .B(n1123), .ZN(G6) );
NOR2_X1 U805 ( .A1(n1108), .A2(n1124), .ZN(G57) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U807 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U808 ( .A1(n1119), .A2(G472), .ZN(n1128) );
NAND2_X1 U809 ( .A1(n1129), .A2(KEYINPUT10), .ZN(n1127) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U811 ( .A1(KEYINPUT5), .A2(n1132), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1108), .A2(n1133), .ZN(G54) );
XOR2_X1 U813 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U814 ( .A(n1086), .B(n1136), .ZN(n1135) );
XNOR2_X1 U815 ( .A(G110), .B(G140), .ZN(n1136) );
INV_X1 U816 ( .A(n1137), .ZN(n1086) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1134) );
XOR2_X1 U818 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U819 ( .A1(G469), .A2(n1119), .ZN(n1140) );
INV_X1 U820 ( .A(n1113), .ZN(n1119) );
NOR2_X1 U821 ( .A1(n1108), .A2(n1142), .ZN(G51) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U823 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U824 ( .A1(KEYINPUT31), .A2(n1147), .ZN(n1146) );
NAND2_X1 U825 ( .A1(KEYINPUT62), .A2(n1148), .ZN(n1145) );
XNOR2_X1 U826 ( .A(n1149), .B(n1150), .ZN(n1148) );
XNOR2_X1 U827 ( .A(n1151), .B(n1152), .ZN(n1143) );
NAND3_X1 U828 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1151) );
NAND2_X1 U829 ( .A1(KEYINPUT55), .A2(n1113), .ZN(n1154) );
NAND2_X1 U830 ( .A1(G902), .A2(n1023), .ZN(n1113) );
NAND2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
INV_X1 U832 ( .A(KEYINPUT55), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1023), .A2(n1158), .ZN(n1156) );
NAND4_X1 U834 ( .A1(n1159), .A2(n1160), .A3(n1088), .A4(n1161), .ZN(n1023) );
NOR2_X1 U835 ( .A1(n1100), .A2(n1162), .ZN(n1161) );
XNOR2_X1 U836 ( .A(KEYINPUT21), .B(n1089), .ZN(n1162) );
NAND3_X1 U837 ( .A1(n1053), .A2(n1163), .A3(n1164), .ZN(n1089) );
NAND3_X1 U838 ( .A1(n1123), .A2(n1018), .A3(n1165), .ZN(n1100) );
NAND2_X1 U839 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
OR4_X1 U841 ( .A1(n1170), .A2(n1171), .A3(n1048), .A4(KEYINPUT37), .ZN(n1169) );
NAND2_X1 U842 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
NAND2_X1 U843 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U844 ( .A1(KEYINPUT37), .A2(n1044), .ZN(n1175) );
NAND3_X1 U845 ( .A1(n1172), .A2(n1176), .A3(n1052), .ZN(n1018) );
NAND3_X1 U846 ( .A1(n1172), .A2(n1176), .A3(n1053), .ZN(n1123) );
AND4_X1 U847 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1088) );
AND3_X1 U848 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
OR2_X1 U849 ( .A1(n1184), .A2(KEYINPUT39), .ZN(n1179) );
NAND4_X1 U850 ( .A1(n1048), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1177) );
NAND2_X1 U851 ( .A1(n1188), .A2(n1043), .ZN(n1187) );
NAND3_X1 U852 ( .A1(n1045), .A2(n1053), .A3(KEYINPUT39), .ZN(n1188) );
NAND3_X1 U853 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1186) );
NAND2_X1 U854 ( .A1(n1192), .A2(n1044), .ZN(n1190) );
XNOR2_X1 U855 ( .A(n1053), .B(KEYINPUT43), .ZN(n1192) );
NAND2_X1 U856 ( .A1(n1166), .A2(n1163), .ZN(n1189) );
XOR2_X1 U857 ( .A(KEYINPUT26), .B(n1098), .Z(n1160) );
AND2_X1 U858 ( .A1(n1039), .A2(n1193), .ZN(n1098) );
XNOR2_X1 U859 ( .A(KEYINPUT60), .B(n1194), .ZN(n1193) );
INV_X1 U860 ( .A(n1097), .ZN(n1159) );
NAND3_X1 U861 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1097) );
NAND2_X1 U862 ( .A1(n1039), .A2(n1198), .ZN(n1197) );
XOR2_X1 U863 ( .A(KEYINPUT35), .B(n1199), .Z(n1198) );
NOR2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U865 ( .A(n1202), .B(KEYINPUT2), .Z(n1200) );
NOR2_X1 U866 ( .A1(n1072), .A2(G952), .ZN(n1108) );
XNOR2_X1 U867 ( .A(G146), .B(n1203), .ZN(G48) );
NAND3_X1 U868 ( .A1(n1204), .A2(n1053), .A3(n1164), .ZN(n1203) );
XOR2_X1 U869 ( .A(n1163), .B(KEYINPUT23), .Z(n1204) );
XNOR2_X1 U870 ( .A(G143), .B(n1178), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1164), .A2(n1044), .A3(n1062), .A4(n1205), .ZN(n1178) );
XNOR2_X1 U872 ( .A(G140), .B(n1184), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1206), .A2(n1207), .ZN(n1184) );
XOR2_X1 U874 ( .A(n1208), .B(n1209), .Z(G39) );
XNOR2_X1 U875 ( .A(G137), .B(KEYINPUT6), .ZN(n1209) );
NAND4_X1 U876 ( .A1(n1206), .A2(n1166), .A3(n1210), .A4(n1163), .ZN(n1208) );
XNOR2_X1 U877 ( .A(KEYINPUT63), .B(n1185), .ZN(n1210) );
XNOR2_X1 U878 ( .A(G134), .B(n1181), .ZN(G36) );
NAND4_X1 U879 ( .A1(n1206), .A2(n1044), .A3(n1052), .A4(n1185), .ZN(n1181) );
XNOR2_X1 U880 ( .A(G131), .B(n1211), .ZN(G33) );
NAND3_X1 U881 ( .A1(n1206), .A2(n1044), .A3(n1212), .ZN(n1211) );
NOR3_X1 U882 ( .A1(n1213), .A2(KEYINPUT54), .A3(n1214), .ZN(n1212) );
XNOR2_X1 U883 ( .A(n1215), .B(KEYINPUT30), .ZN(n1214) );
NOR2_X1 U884 ( .A1(n1043), .A2(n1216), .ZN(n1206) );
INV_X1 U885 ( .A(n1191), .ZN(n1043) );
NOR2_X1 U886 ( .A1(n1040), .A2(n1065), .ZN(n1191) );
XOR2_X1 U887 ( .A(n1060), .B(KEYINPUT27), .Z(n1040) );
NAND2_X1 U888 ( .A1(n1217), .A2(n1218), .ZN(G30) );
NAND2_X1 U889 ( .A1(G128), .A2(n1183), .ZN(n1218) );
XOR2_X1 U890 ( .A(n1219), .B(KEYINPUT40), .Z(n1217) );
OR2_X1 U891 ( .A1(n1183), .A2(G128), .ZN(n1219) );
NAND3_X1 U892 ( .A1(n1052), .A2(n1163), .A3(n1164), .ZN(n1183) );
NOR3_X1 U893 ( .A1(n1220), .A2(n1215), .A3(n1216), .ZN(n1164) );
XNOR2_X1 U894 ( .A(G101), .B(n1221), .ZN(G3) );
NOR2_X1 U895 ( .A1(n1222), .A2(KEYINPUT11), .ZN(n1221) );
AND3_X1 U896 ( .A1(n1166), .A2(n1172), .A3(n1044), .ZN(n1222) );
INV_X1 U897 ( .A(n1170), .ZN(n1044) );
XNOR2_X1 U898 ( .A(G125), .B(n1182), .ZN(G27) );
NAND3_X1 U899 ( .A1(n1207), .A2(n1039), .A3(n1223), .ZN(n1182) );
NOR3_X1 U900 ( .A1(n1213), .A2(n1215), .A3(n1174), .ZN(n1207) );
INV_X1 U901 ( .A(n1185), .ZN(n1215) );
NAND2_X1 U902 ( .A1(n1025), .A2(n1224), .ZN(n1185) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1074), .ZN(n1224) );
INV_X1 U904 ( .A(G900), .ZN(n1074) );
INV_X1 U905 ( .A(n1053), .ZN(n1213) );
XOR2_X1 U906 ( .A(n1226), .B(n1227), .Z(G24) );
NOR2_X1 U907 ( .A1(n1171), .A2(n1201), .ZN(n1227) );
NAND4_X1 U908 ( .A1(n1223), .A2(n1176), .A3(n1062), .A4(n1205), .ZN(n1201) );
INV_X1 U909 ( .A(n1037), .ZN(n1176) );
NAND2_X1 U910 ( .A1(n1228), .A2(n1229), .ZN(n1037) );
XNOR2_X1 U911 ( .A(G122), .B(KEYINPUT29), .ZN(n1226) );
XOR2_X1 U912 ( .A(G119), .B(n1230), .Z(G21) );
NOR2_X1 U913 ( .A1(n1220), .A2(n1194), .ZN(n1230) );
NAND4_X1 U914 ( .A1(n1223), .A2(n1166), .A3(n1163), .A4(n1202), .ZN(n1194) );
NAND2_X1 U915 ( .A1(n1231), .A2(n1232), .ZN(n1163) );
NAND3_X1 U916 ( .A1(n1058), .A2(n1233), .A3(n1234), .ZN(n1232) );
INV_X1 U917 ( .A(KEYINPUT33), .ZN(n1234) );
NAND2_X1 U918 ( .A1(KEYINPUT33), .A2(n1045), .ZN(n1231) );
INV_X1 U919 ( .A(n1039), .ZN(n1220) );
XNOR2_X1 U920 ( .A(G116), .B(n1195), .ZN(G18) );
NAND2_X1 U921 ( .A1(n1235), .A2(n1052), .ZN(n1195) );
AND2_X1 U922 ( .A1(n1054), .A2(n1062), .ZN(n1052) );
XNOR2_X1 U923 ( .A(G113), .B(n1196), .ZN(G15) );
NAND2_X1 U924 ( .A1(n1235), .A2(n1053), .ZN(n1196) );
NOR2_X1 U925 ( .A1(n1062), .A2(n1054), .ZN(n1053) );
INV_X1 U926 ( .A(n1205), .ZN(n1054) );
NOR3_X1 U927 ( .A1(n1170), .A2(n1171), .A3(n1033), .ZN(n1235) );
INV_X1 U928 ( .A(n1223), .ZN(n1033) );
NOR2_X1 U929 ( .A1(n1049), .A2(n1063), .ZN(n1223) );
INV_X1 U930 ( .A(n1236), .ZN(n1049) );
NAND2_X1 U931 ( .A1(n1228), .A2(n1237), .ZN(n1170) );
XNOR2_X1 U932 ( .A(KEYINPUT33), .B(n1229), .ZN(n1237) );
XOR2_X1 U933 ( .A(n1233), .B(KEYINPUT48), .Z(n1228) );
XNOR2_X1 U934 ( .A(G110), .B(n1238), .ZN(G12) );
NAND3_X1 U935 ( .A1(n1172), .A2(n1239), .A3(n1045), .ZN(n1238) );
INV_X1 U936 ( .A(n1174), .ZN(n1045) );
NAND2_X1 U937 ( .A1(n1229), .A2(n1233), .ZN(n1174) );
XNOR2_X1 U938 ( .A(n1059), .B(KEYINPUT45), .ZN(n1233) );
XOR2_X1 U939 ( .A(n1240), .B(n1112), .Z(n1059) );
NAND2_X1 U940 ( .A1(G217), .A2(n1241), .ZN(n1112) );
NAND2_X1 U941 ( .A1(n1110), .A2(n1242), .ZN(n1240) );
XNOR2_X1 U942 ( .A(n1243), .B(n1244), .ZN(n1110) );
XOR2_X1 U943 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U944 ( .A(n1247), .B(n1248), .Z(n1246) );
AND3_X1 U945 ( .A1(G221), .A2(n1072), .A3(G234), .ZN(n1248) );
NAND3_X1 U946 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1247) );
OR2_X1 U947 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND3_X1 U948 ( .A1(n1253), .A2(n1252), .A3(KEYINPUT59), .ZN(n1250) );
AND2_X1 U949 ( .A1(KEYINPUT25), .A2(n1082), .ZN(n1253) );
OR2_X1 U950 ( .A1(n1082), .A2(KEYINPUT59), .ZN(n1249) );
NAND2_X1 U951 ( .A1(KEYINPUT34), .A2(n1254), .ZN(n1245) );
XNOR2_X1 U952 ( .A(G110), .B(n1255), .ZN(n1243) );
XOR2_X1 U953 ( .A(G137), .B(G119), .Z(n1255) );
INV_X1 U954 ( .A(n1058), .ZN(n1229) );
XNOR2_X1 U955 ( .A(n1256), .B(G472), .ZN(n1058) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1242), .ZN(n1256) );
XNOR2_X1 U957 ( .A(n1258), .B(n1132), .ZN(n1257) );
XOR2_X1 U958 ( .A(n1259), .B(G101), .Z(n1132) );
NAND2_X1 U959 ( .A1(G210), .A2(n1260), .ZN(n1259) );
NOR2_X1 U960 ( .A1(KEYINPUT20), .A2(n1261), .ZN(n1258) );
XOR2_X1 U961 ( .A(n1262), .B(n1130), .Z(n1261) );
XOR2_X1 U962 ( .A(n1263), .B(n1264), .Z(n1130) );
XNOR2_X1 U963 ( .A(G113), .B(KEYINPUT12), .ZN(n1263) );
NAND2_X1 U964 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
NAND2_X1 U965 ( .A1(n1131), .A2(n1267), .ZN(n1266) );
INV_X1 U966 ( .A(KEYINPUT32), .ZN(n1267) );
XOR2_X1 U967 ( .A(n1268), .B(n1150), .Z(n1131) );
NAND3_X1 U968 ( .A1(n1150), .A2(n1268), .A3(KEYINPUT32), .ZN(n1265) );
XNOR2_X1 U969 ( .A(KEYINPUT8), .B(n1029), .ZN(n1239) );
INV_X1 U970 ( .A(n1166), .ZN(n1029) );
NOR2_X1 U971 ( .A1(n1205), .A2(n1062), .ZN(n1166) );
XOR2_X1 U972 ( .A(n1269), .B(n1270), .Z(n1062) );
XOR2_X1 U973 ( .A(KEYINPUT36), .B(G478), .Z(n1270) );
NAND2_X1 U974 ( .A1(n1118), .A2(n1242), .ZN(n1269) );
NAND2_X1 U975 ( .A1(n1271), .A2(n1272), .ZN(n1118) );
NAND2_X1 U976 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
INV_X1 U977 ( .A(n1275), .ZN(n1274) );
XOR2_X1 U978 ( .A(n1276), .B(KEYINPUT58), .Z(n1273) );
NAND2_X1 U979 ( .A1(n1275), .A2(n1277), .ZN(n1271) );
XOR2_X1 U980 ( .A(n1276), .B(KEYINPUT22), .Z(n1277) );
NAND3_X1 U981 ( .A1(G217), .A2(n1072), .A3(G234), .ZN(n1276) );
XNOR2_X1 U982 ( .A(n1278), .B(n1279), .ZN(n1275) );
XOR2_X1 U983 ( .A(G122), .B(n1280), .Z(n1279) );
XNOR2_X1 U984 ( .A(n1281), .B(G134), .ZN(n1280) );
XOR2_X1 U985 ( .A(n1282), .B(n1283), .Z(n1278) );
XNOR2_X1 U986 ( .A(G107), .B(n1284), .ZN(n1282) );
NOR2_X1 U987 ( .A1(KEYINPUT3), .A2(n1254), .ZN(n1284) );
XNOR2_X1 U988 ( .A(n1285), .B(G475), .ZN(n1205) );
NAND2_X1 U989 ( .A1(n1122), .A2(n1242), .ZN(n1285) );
XOR2_X1 U990 ( .A(n1286), .B(n1287), .Z(n1122) );
XOR2_X1 U991 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U992 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U993 ( .A1(KEYINPUT41), .A2(n1281), .ZN(n1291) );
INV_X1 U994 ( .A(G143), .ZN(n1281) );
NAND2_X1 U995 ( .A1(G214), .A2(n1260), .ZN(n1290) );
NOR2_X1 U996 ( .A1(G953), .A2(G237), .ZN(n1260) );
XNOR2_X1 U997 ( .A(n1083), .B(G122), .ZN(n1288) );
INV_X1 U998 ( .A(G131), .ZN(n1083) );
XNOR2_X1 U999 ( .A(n1292), .B(n1293), .ZN(n1286) );
XNOR2_X1 U1000 ( .A(n1252), .B(n1082), .ZN(n1293) );
XNOR2_X1 U1001 ( .A(G125), .B(n1294), .ZN(n1082) );
INV_X1 U1002 ( .A(G140), .ZN(n1294) );
NOR2_X1 U1003 ( .A1(n1216), .A2(n1171), .ZN(n1172) );
NAND2_X1 U1004 ( .A1(n1039), .A2(n1202), .ZN(n1171) );
NAND2_X1 U1005 ( .A1(n1025), .A2(n1295), .ZN(n1202) );
NAND3_X1 U1006 ( .A1(G902), .A2(n1225), .A3(n1093), .ZN(n1295) );
NOR2_X1 U1007 ( .A1(G898), .A2(n1072), .ZN(n1093) );
NAND3_X1 U1008 ( .A1(n1225), .A2(n1072), .A3(G952), .ZN(n1025) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U1010 ( .A1(n1296), .A2(n1065), .ZN(n1039) );
INV_X1 U1011 ( .A(n1041), .ZN(n1065) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1297), .ZN(n1041) );
INV_X1 U1013 ( .A(n1060), .ZN(n1296) );
XNOR2_X1 U1014 ( .A(n1298), .B(n1155), .ZN(n1060) );
AND2_X1 U1015 ( .A1(G210), .A2(n1297), .ZN(n1155) );
NAND2_X1 U1016 ( .A1(n1299), .A2(n1158), .ZN(n1297) );
INV_X1 U1017 ( .A(G237), .ZN(n1299) );
NAND2_X1 U1018 ( .A1(n1300), .A2(n1242), .ZN(n1298) );
XNOR2_X1 U1019 ( .A(n1301), .B(n1147), .ZN(n1300) );
NAND2_X1 U1020 ( .A1(n1302), .A2(n1303), .ZN(n1147) );
NAND2_X1 U1021 ( .A1(n1106), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1022 ( .A1(KEYINPUT51), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1023 ( .A1(n1107), .A2(KEYINPUT51), .ZN(n1302) );
NOR2_X1 U1024 ( .A1(n1106), .A2(n1105), .ZN(n1107) );
INV_X1 U1025 ( .A(n1305), .ZN(n1105) );
XOR2_X1 U1026 ( .A(G110), .B(n1306), .Z(n1305) );
XOR2_X1 U1027 ( .A(KEYINPUT49), .B(G122), .Z(n1306) );
XNOR2_X1 U1028 ( .A(n1307), .B(n1292), .ZN(n1106) );
XOR2_X1 U1029 ( .A(G104), .B(G113), .Z(n1292) );
XOR2_X1 U1030 ( .A(n1308), .B(n1264), .Z(n1307) );
XNOR2_X1 U1031 ( .A(n1309), .B(n1283), .ZN(n1264) );
XOR2_X1 U1032 ( .A(G116), .B(KEYINPUT57), .Z(n1283) );
XNOR2_X1 U1033 ( .A(G119), .B(KEYINPUT15), .ZN(n1309) );
XOR2_X1 U1034 ( .A(n1152), .B(n1310), .Z(n1301) );
NOR2_X1 U1035 ( .A1(KEYINPUT47), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1036 ( .A(n1312), .B(n1150), .ZN(n1311) );
XOR2_X1 U1037 ( .A(G128), .B(n1313), .Z(n1150) );
NAND2_X1 U1038 ( .A1(KEYINPUT0), .A2(n1149), .ZN(n1312) );
INV_X1 U1039 ( .A(G125), .ZN(n1149) );
NAND2_X1 U1040 ( .A1(n1314), .A2(G224), .ZN(n1152) );
XNOR2_X1 U1041 ( .A(G953), .B(KEYINPUT13), .ZN(n1314) );
INV_X1 U1042 ( .A(n1048), .ZN(n1216) );
NOR2_X1 U1043 ( .A1(n1063), .A2(n1236), .ZN(n1048) );
NOR2_X1 U1044 ( .A1(n1315), .A2(n1064), .ZN(n1236) );
NOR2_X1 U1045 ( .A1(n1066), .A2(G469), .ZN(n1064) );
AND2_X1 U1046 ( .A1(n1316), .A2(n1066), .ZN(n1315) );
NAND2_X1 U1047 ( .A1(n1317), .A2(n1242), .ZN(n1066) );
XNOR2_X1 U1048 ( .A(n1158), .B(KEYINPUT1), .ZN(n1242) );
XOR2_X1 U1049 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1050 ( .A(n1141), .B(n1320), .ZN(n1319) );
NAND2_X1 U1051 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1052 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
INV_X1 U1053 ( .A(n1325), .ZN(n1324) );
XNOR2_X1 U1054 ( .A(KEYINPUT38), .B(n1137), .ZN(n1323) );
NAND2_X1 U1055 ( .A1(n1326), .A2(n1325), .ZN(n1321) );
XNOR2_X1 U1056 ( .A(n1138), .B(KEYINPUT18), .ZN(n1325) );
XOR2_X1 U1057 ( .A(n1308), .B(G104), .Z(n1138) );
XNOR2_X1 U1058 ( .A(G101), .B(n1327), .ZN(n1308) );
XOR2_X1 U1059 ( .A(KEYINPUT53), .B(G107), .Z(n1327) );
XNOR2_X1 U1060 ( .A(KEYINPUT28), .B(n1137), .ZN(n1326) );
NAND2_X1 U1061 ( .A1(n1328), .A2(n1329), .ZN(n1137) );
NAND2_X1 U1062 ( .A1(n1330), .A2(n1254), .ZN(n1329) );
XOR2_X1 U1063 ( .A(KEYINPUT14), .B(n1331), .Z(n1328) );
NOR2_X1 U1064 ( .A1(n1254), .A2(n1330), .ZN(n1331) );
XOR2_X1 U1065 ( .A(n1313), .B(KEYINPUT44), .Z(n1330) );
XNOR2_X1 U1066 ( .A(G143), .B(n1252), .ZN(n1313) );
XNOR2_X1 U1067 ( .A(G146), .B(KEYINPUT56), .ZN(n1252) );
INV_X1 U1068 ( .A(G128), .ZN(n1254) );
XNOR2_X1 U1069 ( .A(n1332), .B(n1268), .ZN(n1141) );
XNOR2_X1 U1070 ( .A(n1333), .B(n1334), .ZN(n1268) );
NOR2_X1 U1071 ( .A1(G131), .A2(KEYINPUT61), .ZN(n1334) );
XOR2_X1 U1072 ( .A(n1335), .B(G137), .Z(n1333) );
NAND2_X1 U1073 ( .A1(KEYINPUT17), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1074 ( .A(KEYINPUT46), .B(G134), .Z(n1336) );
NAND2_X1 U1075 ( .A1(G227), .A2(n1072), .ZN(n1332) );
INV_X1 U1076 ( .A(G953), .ZN(n1072) );
XOR2_X1 U1077 ( .A(n1337), .B(n1338), .Z(n1318) );
XNOR2_X1 U1078 ( .A(G140), .B(KEYINPUT19), .ZN(n1338) );
NAND2_X1 U1079 ( .A1(KEYINPUT52), .A2(n1339), .ZN(n1337) );
INV_X1 U1080 ( .A(G110), .ZN(n1339) );
XNOR2_X1 U1081 ( .A(G469), .B(KEYINPUT16), .ZN(n1316) );
INV_X1 U1082 ( .A(n1050), .ZN(n1063) );
NAND2_X1 U1083 ( .A1(G221), .A2(n1241), .ZN(n1050) );
NAND2_X1 U1084 ( .A1(G234), .A2(n1158), .ZN(n1241) );
INV_X1 U1085 ( .A(G902), .ZN(n1158) );
endmodule


