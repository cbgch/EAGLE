//Key = 0101010011010010111100010111101001011000110101111011111101110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365;

XNOR2_X1 U747 ( .A(G107), .B(n1034), .ZN(G9) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
XOR2_X1 U750 ( .A(KEYINPUT20), .B(n1041), .Z(n1038) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
AND4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(KEYINPUT43), .ZN(n1048) );
NOR3_X1 U757 ( .A1(n1051), .A2(n1055), .A3(n1056), .ZN(n1044) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR3_X1 U759 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR3_X1 U760 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1058) );
XOR2_X1 U761 ( .A(KEYINPUT15), .B(n1066), .Z(n1063) );
NOR2_X1 U762 ( .A1(KEYINPUT43), .A2(n1047), .ZN(n1057) );
INV_X1 U763 ( .A(n1067), .ZN(n1047) );
NAND3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1037) );
NAND2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND3_X1 U767 ( .A1(n1075), .A2(n1076), .A3(n1067), .ZN(n1074) );
NAND2_X1 U768 ( .A1(n1052), .A2(n1077), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1080), .ZN(n1079) );
NAND2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
OR2_X1 U773 ( .A1(n1064), .A2(n1085), .ZN(n1081) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1086), .ZN(n1078) );
NOR2_X1 U775 ( .A1(n1062), .A2(n1064), .ZN(n1067) );
INV_X1 U776 ( .A(n1084), .ZN(n1062) );
INV_X1 U777 ( .A(n1043), .ZN(n1071) );
NOR3_X1 U778 ( .A1(n1087), .A2(G953), .A3(G952), .ZN(n1035) );
INV_X1 U779 ( .A(n1068), .ZN(n1087) );
NAND4_X1 U780 ( .A1(n1088), .A2(n1089), .A3(n1084), .A4(n1090), .ZN(n1068) );
NOR4_X1 U781 ( .A1(n1054), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1090) );
XNOR2_X1 U782 ( .A(n1094), .B(KEYINPUT9), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(n1092) );
XNOR2_X1 U784 ( .A(n1097), .B(KEYINPUT26), .ZN(n1095) );
XOR2_X1 U785 ( .A(n1053), .B(KEYINPUT14), .Z(n1091) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(G72) );
NOR2_X1 U787 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U789 ( .A(KEYINPUT11), .B(n1104), .Z(n1103) );
NOR2_X1 U790 ( .A1(G953), .A2(n1105), .ZN(n1102) );
NOR3_X1 U791 ( .A1(n1105), .A2(G953), .A3(n1104), .ZN(n1100) );
AND3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1104) );
NAND2_X1 U793 ( .A1(G953), .A2(n1109), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
XNOR2_X1 U795 ( .A(n1112), .B(KEYINPUT39), .ZN(n1110) );
NAND2_X1 U796 ( .A1(n1113), .A2(G125), .ZN(n1106) );
XNOR2_X1 U797 ( .A(KEYINPUT44), .B(n1114), .ZN(n1113) );
INV_X1 U798 ( .A(n1112), .ZN(n1114) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1112) );
NOR2_X1 U800 ( .A1(KEYINPUT21), .A2(n1117), .ZN(n1116) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U802 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U803 ( .A1(G131), .A2(KEYINPUT56), .ZN(n1121) );
XNOR2_X1 U804 ( .A(n1122), .B(n1123), .ZN(n1118) );
NAND2_X1 U805 ( .A1(KEYINPUT1), .A2(G134), .ZN(n1122) );
XNOR2_X1 U806 ( .A(n1040), .B(KEYINPUT31), .ZN(n1105) );
NAND2_X1 U807 ( .A1(G953), .A2(n1124), .ZN(n1098) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1124) );
NAND2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1127), .A2(n1069), .ZN(n1126) );
XNOR2_X1 U811 ( .A(n1039), .B(n1128), .ZN(n1127) );
NAND2_X1 U812 ( .A1(n1129), .A2(G953), .ZN(n1125) );
NAND2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U814 ( .A1(n1132), .A2(G224), .ZN(n1131) );
INV_X1 U815 ( .A(n1128), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1133), .A2(n1128), .ZN(n1130) );
NAND2_X1 U817 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
NAND2_X1 U818 ( .A1(G953), .A2(n1136), .ZN(n1135) );
XOR2_X1 U819 ( .A(n1137), .B(KEYINPUT2), .Z(n1134) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1133) );
NOR2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(G66) );
NOR3_X1 U822 ( .A1(n1097), .A2(n1140), .A3(n1141), .ZN(n1139) );
NOR4_X1 U823 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
INV_X1 U824 ( .A(n1146), .ZN(n1142) );
NOR2_X1 U825 ( .A1(n1147), .A2(n1146), .ZN(n1140) );
NOR3_X1 U826 ( .A1(n1143), .A2(n1148), .A3(n1144), .ZN(n1147) );
NOR2_X1 U827 ( .A1(n1039), .A2(n1040), .ZN(n1148) );
INV_X1 U828 ( .A(KEYINPUT40), .ZN(n1143) );
NOR2_X1 U829 ( .A1(n1138), .A2(n1149), .ZN(G63) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U831 ( .A1(n1152), .A2(n1145), .ZN(n1150) );
INV_X1 U832 ( .A(G478), .ZN(n1152) );
NOR2_X1 U833 ( .A1(n1138), .A2(n1153), .ZN(G60) );
XOR2_X1 U834 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U835 ( .A1(n1156), .A2(n1145), .ZN(n1154) );
XNOR2_X1 U836 ( .A(G104), .B(n1157), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1138), .A2(n1158), .ZN(G57) );
XOR2_X1 U838 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U839 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
NOR3_X1 U840 ( .A1(n1145), .A2(n1163), .A3(n1164), .ZN(n1162) );
NOR2_X1 U841 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
AND2_X1 U842 ( .A1(n1167), .A2(KEYINPUT19), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1168), .A2(n1167), .ZN(n1161) );
XNOR2_X1 U844 ( .A(n1169), .B(n1170), .ZN(n1167) );
XNOR2_X1 U845 ( .A(n1171), .B(n1172), .ZN(n1169) );
NAND2_X1 U846 ( .A1(KEYINPUT45), .A2(n1173), .ZN(n1171) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1168) );
INV_X1 U848 ( .A(KEYINPUT19), .ZN(n1175) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1166), .ZN(n1174) );
INV_X1 U850 ( .A(KEYINPUT35), .ZN(n1166) );
NOR2_X1 U851 ( .A1(n1164), .A2(n1145), .ZN(n1176) );
INV_X1 U852 ( .A(G472), .ZN(n1164) );
NOR2_X1 U853 ( .A1(n1138), .A2(n1177), .ZN(G54) );
XNOR2_X1 U854 ( .A(n1178), .B(n1179), .ZN(n1177) );
XOR2_X1 U855 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U856 ( .A1(n1182), .A2(n1145), .ZN(n1181) );
NOR2_X1 U857 ( .A1(KEYINPUT29), .A2(n1183), .ZN(n1180) );
XOR2_X1 U858 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U859 ( .A1(KEYINPUT61), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U860 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U861 ( .A1(G110), .A2(KEYINPUT37), .ZN(n1187) );
XOR2_X1 U862 ( .A(n1189), .B(KEYINPUT27), .Z(n1184) );
NOR2_X1 U863 ( .A1(n1138), .A2(n1190), .ZN(G51) );
XOR2_X1 U864 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U865 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U866 ( .A(n1195), .B(KEYINPUT59), .Z(n1194) );
NOR2_X1 U867 ( .A1(n1196), .A2(n1145), .ZN(n1191) );
NAND2_X1 U868 ( .A1(G902), .A2(n1197), .ZN(n1145) );
OR2_X1 U869 ( .A1(n1040), .A2(n1039), .ZN(n1197) );
NAND4_X1 U870 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1039) );
AND4_X1 U871 ( .A1(n1202), .A2(n1157), .A3(n1203), .A4(n1204), .ZN(n1201) );
OR3_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1157) );
NOR3_X1 U873 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1200) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1034), .ZN(n1210) );
OR3_X1 U875 ( .A1(n1206), .A2(n1050), .A3(n1205), .ZN(n1034) );
INV_X1 U876 ( .A(KEYINPUT47), .ZN(n1211) );
NOR4_X1 U877 ( .A1(KEYINPUT47), .A2(n1205), .A3(n1212), .A4(n1050), .ZN(n1209) );
NAND3_X1 U878 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1205) );
NOR2_X1 U879 ( .A1(n1206), .A2(n1216), .ZN(n1208) );
OR2_X1 U880 ( .A1(n1217), .A2(n1085), .ZN(n1198) );
NAND2_X1 U881 ( .A1(n1218), .A2(n1219), .ZN(n1040) );
AND4_X1 U882 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
NOR4_X1 U883 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1218) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NOR3_X1 U885 ( .A1(n1207), .A2(n1230), .A3(n1231), .ZN(n1226) );
INV_X1 U886 ( .A(n1232), .ZN(n1225) );
NOR2_X1 U887 ( .A1(n1069), .A2(G952), .ZN(n1138) );
XNOR2_X1 U888 ( .A(G146), .B(n1232), .ZN(G48) );
NAND4_X1 U889 ( .A1(n1075), .A2(n1233), .A3(n1061), .A4(n1086), .ZN(n1232) );
XOR2_X1 U890 ( .A(G143), .B(n1234), .Z(G45) );
NOR3_X1 U891 ( .A1(n1229), .A2(KEYINPUT42), .A3(n1228), .ZN(n1234) );
NAND3_X1 U892 ( .A1(n1083), .A2(n1086), .A3(n1235), .ZN(n1229) );
NOR3_X1 U893 ( .A1(n1085), .A2(n1236), .A3(n1237), .ZN(n1235) );
XOR2_X1 U894 ( .A(G140), .B(n1224), .Z(G42) );
NOR4_X1 U895 ( .A1(n1060), .A2(n1207), .A3(n1230), .A4(n1061), .ZN(n1224) );
INV_X1 U896 ( .A(n1075), .ZN(n1207) );
XNOR2_X1 U897 ( .A(G137), .B(n1223), .ZN(G39) );
NAND3_X1 U898 ( .A1(n1061), .A2(n1238), .A3(n1239), .ZN(n1223) );
XNOR2_X1 U899 ( .A(G134), .B(n1220), .ZN(G36) );
NAND3_X1 U900 ( .A1(n1238), .A2(n1240), .A3(n1083), .ZN(n1220) );
XNOR2_X1 U901 ( .A(G131), .B(n1241), .ZN(G33) );
NAND4_X1 U902 ( .A1(KEYINPUT57), .A2(n1075), .A3(n1083), .A4(n1238), .ZN(n1241) );
INV_X1 U903 ( .A(n1230), .ZN(n1238) );
NAND3_X1 U904 ( .A1(n1086), .A2(n1242), .A3(n1084), .ZN(n1230) );
NOR2_X1 U905 ( .A1(n1066), .A2(n1243), .ZN(n1084) );
INV_X1 U906 ( .A(n1065), .ZN(n1243) );
XOR2_X1 U907 ( .A(n1222), .B(n1244), .Z(G30) );
XNOR2_X1 U908 ( .A(G128), .B(KEYINPUT24), .ZN(n1244) );
NAND4_X1 U909 ( .A1(n1061), .A2(n1233), .A3(n1213), .A4(n1240), .ZN(n1222) );
NAND2_X1 U910 ( .A1(n1245), .A2(n1246), .ZN(G3) );
OR2_X1 U911 ( .A1(n1199), .A2(G101), .ZN(n1246) );
XOR2_X1 U912 ( .A(n1247), .B(KEYINPUT13), .Z(n1245) );
NAND2_X1 U913 ( .A1(G101), .A2(n1199), .ZN(n1247) );
NAND3_X1 U914 ( .A1(n1213), .A2(n1052), .A3(n1248), .ZN(n1199) );
XNOR2_X1 U915 ( .A(G125), .B(n1221), .ZN(G27) );
NAND4_X1 U916 ( .A1(n1075), .A2(n1076), .A3(n1233), .A4(n1249), .ZN(n1221) );
NOR3_X1 U917 ( .A1(n1085), .A2(n1236), .A3(n1060), .ZN(n1233) );
INV_X1 U918 ( .A(n1242), .ZN(n1236) );
NAND2_X1 U919 ( .A1(n1043), .A2(n1250), .ZN(n1242) );
NAND4_X1 U920 ( .A1(G953), .A2(G902), .A3(n1109), .A4(n1251), .ZN(n1250) );
XOR2_X1 U921 ( .A(KEYINPUT18), .B(G900), .Z(n1109) );
XNOR2_X1 U922 ( .A(G122), .B(n1204), .ZN(G24) );
NAND4_X1 U923 ( .A1(n1252), .A2(n1215), .A3(n1076), .A4(n1253), .ZN(n1204) );
NOR3_X1 U924 ( .A1(n1085), .A2(n1254), .A3(n1237), .ZN(n1253) );
INV_X1 U925 ( .A(n1064), .ZN(n1215) );
NAND2_X1 U926 ( .A1(n1249), .A2(n1060), .ZN(n1064) );
XNOR2_X1 U927 ( .A(n1255), .B(n1256), .ZN(G21) );
NOR2_X1 U928 ( .A1(n1085), .A2(n1257), .ZN(n1256) );
XOR2_X1 U929 ( .A(n1217), .B(KEYINPUT38), .Z(n1257) );
NAND4_X1 U930 ( .A1(n1239), .A2(n1076), .A3(n1061), .A4(n1214), .ZN(n1217) );
XNOR2_X1 U931 ( .A(G116), .B(n1202), .ZN(G18) );
NAND4_X1 U932 ( .A1(n1076), .A2(n1083), .A3(n1258), .A4(n1240), .ZN(n1202) );
INV_X1 U933 ( .A(n1050), .ZN(n1240) );
NAND2_X1 U934 ( .A1(n1259), .A2(n1252), .ZN(n1050) );
XNOR2_X1 U935 ( .A(KEYINPUT49), .B(n1094), .ZN(n1259) );
NOR2_X1 U936 ( .A1(n1254), .A2(n1085), .ZN(n1258) );
XNOR2_X1 U937 ( .A(n1212), .B(KEYINPUT60), .ZN(n1085) );
INV_X1 U938 ( .A(n1231), .ZN(n1083) );
XNOR2_X1 U939 ( .A(G113), .B(n1203), .ZN(G15) );
NAND3_X1 U940 ( .A1(n1075), .A2(n1076), .A3(n1248), .ZN(n1203) );
NOR3_X1 U941 ( .A1(n1206), .A2(n1254), .A3(n1231), .ZN(n1248) );
NAND2_X1 U942 ( .A1(n1061), .A2(n1060), .ZN(n1231) );
INV_X1 U943 ( .A(n1249), .ZN(n1061) );
INV_X1 U944 ( .A(n1214), .ZN(n1254) );
INV_X1 U945 ( .A(n1051), .ZN(n1076) );
NAND2_X1 U946 ( .A1(n1053), .A2(n1260), .ZN(n1051) );
XNOR2_X1 U947 ( .A(G110), .B(n1261), .ZN(G12) );
NAND2_X1 U948 ( .A1(n1262), .A2(n1212), .ZN(n1261) );
INV_X1 U949 ( .A(n1206), .ZN(n1212) );
NAND2_X1 U950 ( .A1(n1066), .A2(n1065), .ZN(n1206) );
NAND2_X1 U951 ( .A1(G214), .A2(n1263), .ZN(n1065) );
XOR2_X1 U952 ( .A(n1264), .B(n1196), .Z(n1066) );
NAND2_X1 U953 ( .A1(G210), .A2(n1263), .ZN(n1196) );
NAND2_X1 U954 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
INV_X1 U955 ( .A(G237), .ZN(n1265) );
NAND3_X1 U956 ( .A1(n1267), .A2(n1268), .A3(n1266), .ZN(n1264) );
NAND2_X1 U957 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
INV_X1 U958 ( .A(KEYINPUT63), .ZN(n1270) );
NAND2_X1 U959 ( .A1(n1271), .A2(n1195), .ZN(n1269) );
NAND2_X1 U960 ( .A1(n1137), .A2(n1272), .ZN(n1195) );
INV_X1 U961 ( .A(n1193), .ZN(n1271) );
NOR2_X1 U962 ( .A1(n1272), .A2(n1137), .ZN(n1193) );
NAND2_X1 U963 ( .A1(KEYINPUT63), .A2(n1273), .ZN(n1267) );
XOR2_X1 U964 ( .A(n1137), .B(n1272), .Z(n1273) );
XOR2_X1 U965 ( .A(n1274), .B(n1173), .Z(n1272) );
XNOR2_X1 U966 ( .A(G125), .B(n1275), .ZN(n1274) );
AND2_X1 U967 ( .A1(n1069), .A2(G224), .ZN(n1275) );
XNOR2_X1 U968 ( .A(n1276), .B(n1277), .ZN(n1137) );
XOR2_X1 U969 ( .A(n1278), .B(n1279), .Z(n1276) );
XOR2_X1 U970 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U971 ( .A(KEYINPUT6), .B(KEYINPUT58), .Z(n1280) );
XOR2_X1 U972 ( .A(n1282), .B(n1283), .Z(n1278) );
XNOR2_X1 U973 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND2_X1 U974 ( .A1(KEYINPUT3), .A2(n1286), .ZN(n1284) );
INV_X1 U975 ( .A(G104), .ZN(n1286) );
XNOR2_X1 U976 ( .A(n1287), .B(n1288), .ZN(n1282) );
NAND2_X1 U977 ( .A1(KEYINPUT55), .A2(n1255), .ZN(n1288) );
NAND2_X1 U978 ( .A1(n1289), .A2(KEYINPUT51), .ZN(n1287) );
XNOR2_X1 U979 ( .A(G110), .B(KEYINPUT0), .ZN(n1289) );
XOR2_X1 U980 ( .A(n1216), .B(KEYINPUT16), .Z(n1262) );
NAND4_X1 U981 ( .A1(n1213), .A2(n1239), .A3(n1249), .A4(n1214), .ZN(n1216) );
NAND2_X1 U982 ( .A1(n1043), .A2(n1290), .ZN(n1214) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1136), .ZN(n1290) );
INV_X1 U984 ( .A(G898), .ZN(n1136) );
NAND3_X1 U985 ( .A1(n1251), .A2(n1069), .A3(G952), .ZN(n1043) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1251) );
XNOR2_X1 U987 ( .A(n1088), .B(KEYINPUT30), .ZN(n1249) );
XNOR2_X1 U988 ( .A(G472), .B(n1291), .ZN(n1088) );
NOR2_X1 U989 ( .A1(n1292), .A2(G902), .ZN(n1291) );
NOR2_X1 U990 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U991 ( .A(n1295), .B(KEYINPUT41), .Z(n1294) );
NAND2_X1 U992 ( .A1(n1296), .A2(n1160), .ZN(n1295) );
NOR2_X1 U993 ( .A1(n1296), .A2(n1160), .ZN(n1293) );
XNOR2_X1 U994 ( .A(n1297), .B(G101), .ZN(n1160) );
NAND2_X1 U995 ( .A1(G210), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U996 ( .A(n1299), .B(n1173), .ZN(n1296) );
XNOR2_X1 U997 ( .A(n1300), .B(n1301), .ZN(n1173) );
XNOR2_X1 U998 ( .A(n1302), .B(n1303), .ZN(n1299) );
NAND2_X1 U999 ( .A1(KEYINPUT62), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1000 ( .A1(KEYINPUT33), .A2(n1172), .ZN(n1302) );
XOR2_X1 U1001 ( .A(n1305), .B(n1306), .Z(n1172) );
XNOR2_X1 U1002 ( .A(KEYINPUT32), .B(n1255), .ZN(n1306) );
INV_X1 U1003 ( .A(G119), .ZN(n1255) );
XOR2_X1 U1004 ( .A(n1307), .B(G116), .Z(n1305) );
NAND2_X1 U1005 ( .A1(KEYINPUT54), .A2(n1277), .ZN(n1307) );
INV_X1 U1006 ( .A(G113), .ZN(n1277) );
NOR2_X1 U1007 ( .A1(n1060), .A2(n1056), .ZN(n1239) );
INV_X1 U1008 ( .A(n1052), .ZN(n1056) );
NAND2_X1 U1009 ( .A1(n1308), .A2(n1309), .ZN(n1052) );
OR3_X1 U1010 ( .A1(n1252), .A2(n1094), .A3(KEYINPUT49), .ZN(n1309) );
NAND2_X1 U1011 ( .A1(KEYINPUT49), .A2(n1075), .ZN(n1308) );
NOR2_X1 U1012 ( .A1(n1237), .A2(n1252), .ZN(n1075) );
INV_X1 U1013 ( .A(n1228), .ZN(n1252) );
XOR2_X1 U1014 ( .A(n1310), .B(n1089), .Z(n1228) );
XOR2_X1 U1015 ( .A(n1311), .B(G478), .Z(n1089) );
OR2_X1 U1016 ( .A1(n1151), .A2(G902), .ZN(n1311) );
XNOR2_X1 U1017 ( .A(n1312), .B(n1313), .ZN(n1151) );
XOR2_X1 U1018 ( .A(G107), .B(n1281), .Z(n1313) );
XNOR2_X1 U1019 ( .A(n1314), .B(G116), .ZN(n1281) );
XOR2_X1 U1020 ( .A(n1315), .B(n1316), .Z(n1312) );
NOR2_X1 U1021 ( .A1(n1144), .A2(n1317), .ZN(n1316) );
INV_X1 U1022 ( .A(G217), .ZN(n1144) );
NAND2_X1 U1023 ( .A1(KEYINPUT23), .A2(n1318), .ZN(n1315) );
XOR2_X1 U1024 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1025 ( .A(G134), .B(n1300), .ZN(n1320) );
NOR2_X1 U1026 ( .A1(KEYINPUT10), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1027 ( .A(G143), .B(KEYINPUT53), .ZN(n1321) );
XNOR2_X1 U1028 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n1310) );
INV_X1 U1029 ( .A(n1094), .ZN(n1237) );
XOR2_X1 U1030 ( .A(n1322), .B(n1156), .Z(n1094) );
INV_X1 U1031 ( .A(G475), .ZN(n1156) );
OR2_X1 U1032 ( .A1(n1155), .A2(G902), .ZN(n1322) );
XOR2_X1 U1033 ( .A(n1323), .B(n1188), .Z(n1155) );
INV_X1 U1034 ( .A(n1115), .ZN(n1188) );
XOR2_X1 U1035 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1036 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1037 ( .A(n1111), .B(G113), .ZN(n1327) );
INV_X1 U1038 ( .A(G125), .ZN(n1111) );
XOR2_X1 U1039 ( .A(KEYINPUT28), .B(G131), .Z(n1326) );
XOR2_X1 U1040 ( .A(n1328), .B(n1329), .Z(n1324) );
XNOR2_X1 U1041 ( .A(G104), .B(n1330), .ZN(n1329) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1298), .ZN(n1330) );
NOR2_X1 U1043 ( .A1(G953), .A2(G237), .ZN(n1298) );
XNOR2_X1 U1044 ( .A(n1331), .B(n1301), .ZN(n1328) );
NAND2_X1 U1045 ( .A1(KEYINPUT46), .A2(n1314), .ZN(n1331) );
INV_X1 U1046 ( .A(G122), .ZN(n1314) );
XNOR2_X1 U1047 ( .A(n1332), .B(n1096), .ZN(n1060) );
AND2_X1 U1048 ( .A1(G217), .A2(n1333), .ZN(n1096) );
XNOR2_X1 U1049 ( .A(KEYINPUT5), .B(n1334), .ZN(n1333) );
NAND2_X1 U1050 ( .A1(KEYINPUT48), .A2(n1335), .ZN(n1332) );
INV_X1 U1051 ( .A(n1097), .ZN(n1335) );
NOR2_X1 U1052 ( .A1(n1146), .A2(G902), .ZN(n1097) );
XNOR2_X1 U1053 ( .A(n1336), .B(n1337), .ZN(n1146) );
XNOR2_X1 U1054 ( .A(G137), .B(n1338), .ZN(n1337) );
NAND3_X1 U1055 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NAND2_X1 U1056 ( .A1(KEYINPUT12), .A2(n1342), .ZN(n1341) );
OR3_X1 U1057 ( .A1(n1342), .A2(KEYINPUT12), .A3(n1343), .ZN(n1340) );
NAND2_X1 U1058 ( .A1(n1343), .A2(n1344), .ZN(n1339) );
NAND2_X1 U1059 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
INV_X1 U1060 ( .A(KEYINPUT12), .ZN(n1346) );
XOR2_X1 U1061 ( .A(KEYINPUT52), .B(n1342), .Z(n1345) );
XOR2_X1 U1062 ( .A(G110), .B(n1347), .Z(n1342) );
XNOR2_X1 U1063 ( .A(n1300), .B(G119), .ZN(n1347) );
INV_X1 U1064 ( .A(G128), .ZN(n1300) );
XNOR2_X1 U1065 ( .A(n1348), .B(n1349), .ZN(n1343) );
XNOR2_X1 U1066 ( .A(n1350), .B(G125), .ZN(n1349) );
INV_X1 U1067 ( .A(G146), .ZN(n1350) );
NAND2_X1 U1068 ( .A1(KEYINPUT50), .A2(n1115), .ZN(n1348) );
NAND2_X1 U1069 ( .A1(G221), .A2(n1351), .ZN(n1336) );
INV_X1 U1070 ( .A(n1317), .ZN(n1351) );
NAND2_X1 U1071 ( .A1(G234), .A2(n1069), .ZN(n1317) );
XNOR2_X1 U1072 ( .A(n1086), .B(KEYINPUT36), .ZN(n1213) );
NOR2_X1 U1073 ( .A1(n1053), .A2(n1054), .ZN(n1086) );
INV_X1 U1074 ( .A(n1260), .ZN(n1054) );
NAND2_X1 U1075 ( .A1(G221), .A2(n1334), .ZN(n1260) );
NAND2_X1 U1076 ( .A1(G234), .A2(n1266), .ZN(n1334) );
XNOR2_X1 U1077 ( .A(n1352), .B(n1182), .ZN(n1053) );
INV_X1 U1078 ( .A(G469), .ZN(n1182) );
NAND2_X1 U1079 ( .A1(n1353), .A2(n1266), .ZN(n1352) );
INV_X1 U1080 ( .A(G902), .ZN(n1266) );
XNOR2_X1 U1081 ( .A(n1354), .B(n1355), .ZN(n1353) );
XOR2_X1 U1082 ( .A(n1189), .B(n1356), .Z(n1355) );
NAND2_X1 U1083 ( .A1(n1357), .A2(KEYINPUT17), .ZN(n1356) );
XNOR2_X1 U1084 ( .A(G110), .B(n1115), .ZN(n1357) );
XOR2_X1 U1085 ( .A(G140), .B(KEYINPUT25), .Z(n1115) );
NAND2_X1 U1086 ( .A1(G227), .A2(n1069), .ZN(n1189) );
INV_X1 U1087 ( .A(G953), .ZN(n1069) );
INV_X1 U1088 ( .A(n1178), .ZN(n1354) );
XNOR2_X1 U1089 ( .A(n1358), .B(n1359), .ZN(n1178) );
XNOR2_X1 U1090 ( .A(n1120), .B(n1304), .ZN(n1359) );
INV_X1 U1091 ( .A(n1170), .ZN(n1304) );
NAND2_X1 U1092 ( .A1(n1360), .A2(n1361), .ZN(n1170) );
NAND2_X1 U1093 ( .A1(n1362), .A2(G137), .ZN(n1361) );
NAND2_X1 U1094 ( .A1(n1363), .A2(n1123), .ZN(n1360) );
INV_X1 U1095 ( .A(G137), .ZN(n1123) );
XNOR2_X1 U1096 ( .A(n1362), .B(KEYINPUT4), .ZN(n1363) );
XOR2_X1 U1097 ( .A(G131), .B(G134), .Z(n1362) );
XNOR2_X1 U1098 ( .A(G128), .B(n1364), .ZN(n1120) );
NOR2_X1 U1099 ( .A1(KEYINPUT22), .A2(n1301), .ZN(n1364) );
XNOR2_X1 U1100 ( .A(G143), .B(G146), .ZN(n1301) );
XOR2_X1 U1101 ( .A(n1365), .B(n1285), .Z(n1358) );
XOR2_X1 U1102 ( .A(G107), .B(G101), .Z(n1285) );
XNOR2_X1 U1103 ( .A(G104), .B(KEYINPUT34), .ZN(n1365) );
endmodule


