//Key = 0101110100011101100000010100000111000110010000000101000010000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;

XOR2_X1 U725 ( .A(G107), .B(n1009), .Z(G9) );
NOR3_X1 U726 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1009) );
NOR2_X1 U727 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR3_X1 U728 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NOR2_X1 U729 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U730 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
XOR2_X1 U731 ( .A(KEYINPUT62), .B(n1022), .Z(n1021) );
NOR3_X1 U732 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR2_X1 U733 ( .A1(n1026), .A2(n1023), .ZN(n1020) );
NAND3_X1 U734 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1023) );
NAND3_X1 U735 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1015) );
NAND3_X1 U736 ( .A1(n1033), .A2(n1034), .A3(n1029), .ZN(n1032) );
INV_X1 U737 ( .A(n1035), .ZN(n1029) );
NAND2_X1 U738 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND3_X1 U739 ( .A1(n1027), .A2(n1038), .A3(n1039), .ZN(n1037) );
NAND2_X1 U740 ( .A1(n1010), .A2(n1040), .ZN(n1038) );
NAND2_X1 U741 ( .A1(n1028), .A2(n1041), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U743 ( .A1(n1039), .A2(n1044), .ZN(n1043) );
OR2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U745 ( .A1(n1027), .A2(n1047), .ZN(n1042) );
NAND2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U747 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR3_X1 U748 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1013) );
INV_X1 U749 ( .A(n1030), .ZN(n1052) );
NAND4_X1 U750 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1030) );
NOR4_X1 U751 ( .A1(n1057), .A2(n1050), .A3(n1058), .A4(n1059), .ZN(n1056) );
XNOR2_X1 U752 ( .A(n1060), .B(KEYINPUT42), .ZN(n1059) );
XOR2_X1 U753 ( .A(n1061), .B(n1062), .Z(n1058) );
NOR2_X1 U754 ( .A1(KEYINPUT53), .A2(n1063), .ZN(n1062) );
XNOR2_X1 U755 ( .A(G478), .B(KEYINPUT27), .ZN(n1061) );
INV_X1 U756 ( .A(n1024), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1055) );
XOR2_X1 U758 ( .A(n1051), .B(KEYINPUT33), .Z(n1064) );
XNOR2_X1 U759 ( .A(G475), .B(n1066), .ZN(n1054) );
NOR2_X1 U760 ( .A1(KEYINPUT46), .A2(n1067), .ZN(n1066) );
XOR2_X1 U761 ( .A(KEYINPUT29), .B(n1068), .Z(n1053) );
NOR2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U763 ( .A1(KEYINPUT14), .A2(n1071), .ZN(n1070) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
INV_X1 U765 ( .A(KEYINPUT14), .ZN(n1073) );
NOR2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
XOR2_X1 U767 ( .A(n1076), .B(n1077), .Z(G72) );
NOR2_X1 U768 ( .A1(n1078), .A2(n1031), .ZN(n1077) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1083), .A2(n1031), .ZN(n1082) );
XOR2_X1 U772 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND3_X1 U774 ( .A1(G900), .A2(n1085), .A3(G953), .ZN(n1081) );
XOR2_X1 U775 ( .A(n1088), .B(n1089), .Z(n1085) );
XOR2_X1 U776 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U777 ( .A1(KEYINPUT9), .A2(n1092), .ZN(n1090) );
XOR2_X1 U778 ( .A(n1093), .B(n1094), .Z(n1088) );
NOR2_X1 U779 ( .A1(KEYINPUT17), .A2(n1095), .ZN(n1094) );
XNOR2_X1 U780 ( .A(KEYINPUT51), .B(n1096), .ZN(n1095) );
XOR2_X1 U781 ( .A(n1097), .B(n1098), .Z(G69) );
XOR2_X1 U782 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U783 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1101) );
NAND3_X1 U785 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1099) );
NAND2_X1 U786 ( .A1(G953), .A2(n1105), .ZN(n1104) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
OR2_X1 U789 ( .A1(n1110), .A2(KEYINPUT63), .ZN(n1109) );
INV_X1 U790 ( .A(n1111), .ZN(n1106) );
NAND3_X1 U791 ( .A1(n1112), .A2(n1113), .A3(KEYINPUT63), .ZN(n1102) );
NAND2_X1 U792 ( .A1(KEYINPUT4), .A2(n1114), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1108), .A2(n1111), .ZN(n1114) );
NAND2_X1 U794 ( .A1(n1108), .A2(n1110), .ZN(n1112) );
INV_X1 U795 ( .A(KEYINPUT4), .ZN(n1110) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1108) );
NOR2_X1 U797 ( .A1(n1117), .A2(G953), .ZN(n1097) );
NOR2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U799 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND4_X1 U800 ( .A1(G217), .A2(n1017), .A3(n1122), .A4(n1123), .ZN(n1120) );
NAND2_X1 U801 ( .A1(G902), .A2(n1124), .ZN(n1123) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NAND2_X1 U803 ( .A1(n1127), .A2(n1124), .ZN(n1125) );
INV_X1 U804 ( .A(KEYINPUT23), .ZN(n1124) );
NOR2_X1 U805 ( .A1(n1118), .A2(n1128), .ZN(G63) );
NOR3_X1 U806 ( .A1(n1063), .A2(n1129), .A3(n1130), .ZN(n1128) );
NOR3_X1 U807 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
NOR2_X1 U808 ( .A1(n1134), .A2(n1135), .ZN(n1129) );
NOR2_X1 U809 ( .A1(n1136), .A2(n1132), .ZN(n1135) );
NOR2_X1 U810 ( .A1(n1118), .A2(n1137), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR3_X1 U812 ( .A1(n1126), .A2(n1140), .A3(n1141), .ZN(n1139) );
XNOR2_X1 U813 ( .A(n1136), .B(KEYINPUT11), .ZN(n1140) );
XNOR2_X1 U814 ( .A(n1142), .B(n1143), .ZN(G6) );
NAND2_X1 U815 ( .A1(KEYINPUT15), .A2(n1144), .ZN(n1142) );
INV_X1 U816 ( .A(G104), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1118), .A2(n1145), .ZN(G57) );
XOR2_X1 U818 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U819 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U820 ( .A1(n1150), .A2(KEYINPUT10), .ZN(n1148) );
XOR2_X1 U821 ( .A(n1151), .B(n1152), .Z(n1146) );
XNOR2_X1 U822 ( .A(G101), .B(n1153), .ZN(n1152) );
NAND2_X1 U823 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND4_X1 U824 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
INV_X1 U825 ( .A(KEYINPUT50), .ZN(n1158) );
NAND2_X1 U826 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
NAND2_X1 U827 ( .A1(n1157), .A2(n1162), .ZN(n1161) );
NAND2_X1 U828 ( .A1(KEYINPUT50), .A2(n1163), .ZN(n1162) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1159), .ZN(n1160) );
INV_X1 U830 ( .A(KEYINPUT55), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1164), .A2(n1133), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1118), .A2(n1165), .ZN(G54) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR3_X1 U834 ( .A1(n1075), .A2(n1136), .A3(n1168), .ZN(n1167) );
XNOR2_X1 U835 ( .A(G902), .B(KEYINPUT0), .ZN(n1168) );
INV_X1 U836 ( .A(n1017), .ZN(n1136) );
NOR2_X1 U837 ( .A1(KEYINPUT24), .A2(n1169), .ZN(n1166) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U839 ( .A(n1172), .B(n1091), .Z(n1171) );
XNOR2_X1 U840 ( .A(n1173), .B(n1092), .ZN(n1172) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1170) );
XNOR2_X1 U842 ( .A(n1176), .B(KEYINPUT31), .ZN(n1175) );
NAND2_X1 U843 ( .A1(n1177), .A2(KEYINPUT37), .ZN(n1176) );
XOR2_X1 U844 ( .A(n1093), .B(KEYINPUT54), .Z(n1177) );
NOR2_X1 U845 ( .A1(n1118), .A2(n1178), .ZN(G51) );
XNOR2_X1 U846 ( .A(n1179), .B(n1180), .ZN(n1178) );
XNOR2_X1 U847 ( .A(n1156), .B(n1181), .ZN(n1180) );
NOR2_X1 U848 ( .A1(n1182), .A2(n1133), .ZN(n1181) );
NAND2_X1 U849 ( .A1(G902), .A2(n1017), .ZN(n1133) );
NAND3_X1 U850 ( .A1(n1117), .A2(n1086), .A3(n1183), .ZN(n1017) );
XOR2_X1 U851 ( .A(n1087), .B(KEYINPUT8), .Z(n1183) );
AND4_X1 U852 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1086) );
NOR4_X1 U853 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NOR4_X1 U856 ( .A1(n1196), .A2(n1197), .A3(n1048), .A4(n1198), .ZN(n1194) );
AND2_X1 U857 ( .A1(KEYINPUT16), .A2(n1199), .ZN(n1189) );
NOR3_X1 U858 ( .A1(KEYINPUT16), .A2(n1200), .A3(n1019), .ZN(n1188) );
AND2_X1 U859 ( .A1(n1201), .A2(n1202), .ZN(n1117) );
AND4_X1 U860 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1143), .ZN(n1202) );
NAND3_X1 U861 ( .A1(n1027), .A2(n1206), .A3(n1207), .ZN(n1143) );
NOR4_X1 U862 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1201) );
NOR3_X1 U863 ( .A1(n1198), .A2(n1212), .A3(n1011), .ZN(n1211) );
NOR4_X1 U864 ( .A1(n1213), .A2(n1214), .A3(n1012), .A4(n1010), .ZN(n1210) );
INV_X1 U865 ( .A(n1215), .ZN(n1010) );
INV_X1 U866 ( .A(n1027), .ZN(n1012) );
NOR2_X1 U867 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
INV_X1 U868 ( .A(KEYINPUT40), .ZN(n1217) );
NOR3_X1 U869 ( .A1(n1026), .A2(n1218), .A3(n1219), .ZN(n1216) );
NOR2_X1 U870 ( .A1(KEYINPUT40), .A2(n1206), .ZN(n1213) );
AND2_X1 U871 ( .A1(n1220), .A2(G953), .ZN(n1118) );
XNOR2_X1 U872 ( .A(G952), .B(KEYINPUT57), .ZN(n1220) );
XOR2_X1 U873 ( .A(G146), .B(n1221), .Z(G48) );
NOR2_X1 U874 ( .A1(KEYINPUT52), .A2(n1087), .ZN(n1221) );
NAND3_X1 U875 ( .A1(n1207), .A2(n1218), .A3(n1222), .ZN(n1087) );
XNOR2_X1 U876 ( .A(G143), .B(n1223), .ZN(G45) );
NAND3_X1 U877 ( .A1(n1224), .A2(n1218), .A3(n1225), .ZN(n1223) );
NOR3_X1 U878 ( .A1(n1197), .A2(KEYINPUT21), .A3(n1196), .ZN(n1225) );
INV_X1 U879 ( .A(n1226), .ZN(n1196) );
XOR2_X1 U880 ( .A(n1227), .B(G140), .Z(G42) );
NAND2_X1 U881 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
OR4_X1 U882 ( .A1(n1230), .A2(n1026), .A3(n1231), .A4(KEYINPUT41), .ZN(n1229) );
NAND3_X1 U883 ( .A1(n1195), .A2(n1232), .A3(KEYINPUT41), .ZN(n1228) );
INV_X1 U884 ( .A(n1230), .ZN(n1195) );
NAND3_X1 U885 ( .A1(n1207), .A2(n1046), .A3(n1039), .ZN(n1230) );
XOR2_X1 U886 ( .A(n1186), .B(n1233), .Z(G39) );
XNOR2_X1 U887 ( .A(G137), .B(KEYINPUT44), .ZN(n1233) );
NAND3_X1 U888 ( .A1(n1222), .A2(n1028), .A3(n1039), .ZN(n1186) );
XOR2_X1 U889 ( .A(G134), .B(n1190), .Z(G36) );
AND3_X1 U890 ( .A1(n1039), .A2(n1215), .A3(n1224), .ZN(n1190) );
XNOR2_X1 U891 ( .A(G131), .B(n1234), .ZN(G33) );
NOR2_X1 U892 ( .A1(n1199), .A2(KEYINPUT30), .ZN(n1234) );
AND2_X1 U893 ( .A1(n1200), .A2(n1039), .ZN(n1199) );
INV_X1 U894 ( .A(n1019), .ZN(n1039) );
NAND2_X1 U895 ( .A1(n1051), .A2(n1235), .ZN(n1019) );
AND2_X1 U896 ( .A1(n1224), .A2(n1207), .ZN(n1200) );
NOR2_X1 U897 ( .A1(n1193), .A2(n1198), .ZN(n1224) );
INV_X1 U898 ( .A(n1232), .ZN(n1193) );
XNOR2_X1 U899 ( .A(G128), .B(n1184), .ZN(G30) );
NAND3_X1 U900 ( .A1(n1215), .A2(n1218), .A3(n1222), .ZN(n1184) );
AND3_X1 U901 ( .A1(n1236), .A2(n1237), .A3(n1232), .ZN(n1222) );
NOR2_X1 U902 ( .A1(n1026), .A2(n1238), .ZN(n1232) );
NAND2_X1 U903 ( .A1(KEYINPUT2), .A2(n1198), .ZN(n1237) );
NAND2_X1 U904 ( .A1(n1239), .A2(n1240), .ZN(n1236) );
INV_X1 U905 ( .A(KEYINPUT2), .ZN(n1240) );
NAND2_X1 U906 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
XOR2_X1 U907 ( .A(n1243), .B(n1244), .Z(G3) );
XNOR2_X1 U908 ( .A(KEYINPUT26), .B(n1245), .ZN(n1244) );
NOR4_X1 U909 ( .A1(KEYINPUT20), .A2(n1212), .A3(n1011), .A4(n1198), .ZN(n1243) );
INV_X1 U910 ( .A(n1045), .ZN(n1198) );
INV_X1 U911 ( .A(n1206), .ZN(n1011) );
INV_X1 U912 ( .A(n1028), .ZN(n1212) );
XOR2_X1 U913 ( .A(n1185), .B(n1246), .Z(G27) );
XNOR2_X1 U914 ( .A(G125), .B(KEYINPUT19), .ZN(n1246) );
NAND4_X1 U915 ( .A1(n1207), .A2(n1033), .A3(n1247), .A4(n1046), .ZN(n1185) );
NOR2_X1 U916 ( .A1(n1238), .A2(n1048), .ZN(n1247) );
INV_X1 U917 ( .A(n1231), .ZN(n1238) );
NAND2_X1 U918 ( .A1(n1035), .A2(n1248), .ZN(n1231) );
NAND4_X1 U919 ( .A1(G953), .A2(G902), .A3(n1249), .A4(n1080), .ZN(n1248) );
INV_X1 U920 ( .A(G900), .ZN(n1080) );
XOR2_X1 U921 ( .A(G122), .B(n1209), .Z(G24) );
AND4_X1 U922 ( .A1(n1250), .A2(n1027), .A3(n1251), .A4(n1226), .ZN(n1209) );
NOR2_X1 U923 ( .A1(n1242), .A2(n1241), .ZN(n1027) );
XOR2_X1 U924 ( .A(G119), .B(n1208), .Z(G21) );
AND4_X1 U925 ( .A1(n1252), .A2(n1250), .A3(n1241), .A4(n1028), .ZN(n1208) );
XNOR2_X1 U926 ( .A(n1060), .B(KEYINPUT2), .ZN(n1252) );
XNOR2_X1 U927 ( .A(G116), .B(n1205), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1045), .A2(n1215), .A3(n1250), .ZN(n1205) );
XNOR2_X1 U929 ( .A(G113), .B(n1204), .ZN(G15) );
NAND3_X1 U930 ( .A1(n1045), .A2(n1207), .A3(n1250), .ZN(n1204) );
AND3_X1 U931 ( .A1(n1218), .A2(n1253), .A3(n1033), .ZN(n1250) );
AND2_X1 U932 ( .A1(n1071), .A2(n1254), .ZN(n1033) );
INV_X1 U933 ( .A(n1040), .ZN(n1207) );
NAND2_X1 U934 ( .A1(n1255), .A2(n1226), .ZN(n1040) );
XNOR2_X1 U935 ( .A(KEYINPUT43), .B(n1251), .ZN(n1255) );
NOR2_X1 U936 ( .A1(n1256), .A2(n1242), .ZN(n1045) );
XNOR2_X1 U937 ( .A(G110), .B(n1203), .ZN(G12) );
NAND3_X1 U938 ( .A1(n1206), .A2(n1028), .A3(n1046), .ZN(n1203) );
NOR2_X1 U939 ( .A1(n1241), .A2(n1060), .ZN(n1046) );
INV_X1 U940 ( .A(n1242), .ZN(n1060) );
NAND3_X1 U941 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1242) );
OR2_X1 U942 ( .A1(n1260), .A2(n1121), .ZN(n1259) );
NAND3_X1 U943 ( .A1(n1121), .A2(n1260), .A3(n1126), .ZN(n1258) );
NAND2_X1 U944 ( .A1(G217), .A2(n1127), .ZN(n1260) );
XOR2_X1 U945 ( .A(n1261), .B(n1262), .Z(n1121) );
XOR2_X1 U946 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U947 ( .A(n1265), .B(n1266), .Z(n1264) );
NOR2_X1 U948 ( .A1(G119), .A2(KEYINPUT61), .ZN(n1266) );
NOR2_X1 U949 ( .A1(n1267), .A2(n1268), .ZN(n1265) );
XOR2_X1 U950 ( .A(n1269), .B(KEYINPUT1), .Z(n1268) );
NAND2_X1 U951 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NOR2_X1 U952 ( .A1(n1270), .A2(n1271), .ZN(n1267) );
XOR2_X1 U953 ( .A(KEYINPUT59), .B(G146), .Z(n1271) );
XNOR2_X1 U954 ( .A(G125), .B(n1272), .ZN(n1270) );
XOR2_X1 U955 ( .A(KEYINPUT12), .B(G140), .Z(n1272) );
AND2_X1 U956 ( .A1(n1273), .A2(G221), .ZN(n1263) );
XNOR2_X1 U957 ( .A(G110), .B(n1274), .ZN(n1261) );
XNOR2_X1 U958 ( .A(G137), .B(n1275), .ZN(n1274) );
NAND2_X1 U959 ( .A1(G902), .A2(G217), .ZN(n1257) );
INV_X1 U960 ( .A(n1256), .ZN(n1241) );
XOR2_X1 U961 ( .A(n1065), .B(KEYINPUT5), .Z(n1256) );
XOR2_X1 U962 ( .A(n1276), .B(n1164), .Z(n1065) );
INV_X1 U963 ( .A(G472), .ZN(n1164) );
NAND2_X1 U964 ( .A1(n1277), .A2(n1126), .ZN(n1276) );
XOR2_X1 U965 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U966 ( .A(n1157), .B(n1149), .Z(n1279) );
XNOR2_X1 U967 ( .A(n1280), .B(n1281), .ZN(n1149) );
NOR2_X1 U968 ( .A1(G113), .A2(KEYINPUT18), .ZN(n1281) );
XNOR2_X1 U969 ( .A(n1156), .B(n1282), .ZN(n1278) );
NAND2_X1 U970 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U971 ( .A1(G101), .A2(n1150), .ZN(n1284) );
INV_X1 U972 ( .A(n1285), .ZN(n1150) );
XOR2_X1 U973 ( .A(n1286), .B(KEYINPUT47), .Z(n1283) );
NAND2_X1 U974 ( .A1(n1245), .A2(n1285), .ZN(n1286) );
NAND3_X1 U975 ( .A1(n1287), .A2(n1031), .A3(G210), .ZN(n1285) );
INV_X1 U976 ( .A(n1163), .ZN(n1156) );
NAND2_X1 U977 ( .A1(n1288), .A2(n1289), .ZN(n1028) );
OR3_X1 U978 ( .A1(n1226), .A2(n1251), .A3(KEYINPUT43), .ZN(n1289) );
INV_X1 U979 ( .A(n1197), .ZN(n1251) );
NAND2_X1 U980 ( .A1(KEYINPUT43), .A2(n1215), .ZN(n1288) );
NOR2_X1 U981 ( .A1(n1226), .A2(n1197), .ZN(n1215) );
XOR2_X1 U982 ( .A(n1063), .B(n1132), .Z(n1197) );
INV_X1 U983 ( .A(G478), .ZN(n1132) );
NOR2_X1 U984 ( .A1(n1134), .A2(G902), .ZN(n1063) );
INV_X1 U985 ( .A(n1131), .ZN(n1134) );
NAND2_X1 U986 ( .A1(n1290), .A2(n1291), .ZN(n1131) );
NAND3_X1 U987 ( .A1(n1292), .A2(n1273), .A3(G217), .ZN(n1291) );
NAND2_X1 U988 ( .A1(n1293), .A2(n1294), .ZN(n1290) );
NAND2_X1 U989 ( .A1(G217), .A2(n1273), .ZN(n1294) );
NOR2_X1 U990 ( .A1(n1127), .A2(G953), .ZN(n1273) );
INV_X1 U991 ( .A(G234), .ZN(n1127) );
XOR2_X1 U992 ( .A(n1292), .B(KEYINPUT32), .Z(n1293) );
XOR2_X1 U993 ( .A(n1295), .B(n1296), .Z(n1292) );
XOR2_X1 U994 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U995 ( .A(n1299), .B(G134), .ZN(n1298) );
INV_X1 U996 ( .A(G143), .ZN(n1299) );
XOR2_X1 U997 ( .A(KEYINPUT60), .B(KEYINPUT28), .Z(n1297) );
XOR2_X1 U998 ( .A(n1300), .B(n1301), .Z(n1295) );
XOR2_X1 U999 ( .A(G122), .B(G116), .Z(n1301) );
XOR2_X1 U1000 ( .A(n1302), .B(G107), .Z(n1300) );
NAND2_X1 U1001 ( .A1(KEYINPUT49), .A2(G128), .ZN(n1302) );
XOR2_X1 U1002 ( .A(n1067), .B(n1141), .Z(n1226) );
INV_X1 U1003 ( .A(G475), .ZN(n1141) );
NAND2_X1 U1004 ( .A1(n1138), .A2(n1126), .ZN(n1067) );
XNOR2_X1 U1005 ( .A(n1303), .B(n1304), .ZN(n1138) );
XOR2_X1 U1006 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1007 ( .A(n1307), .B(G104), .ZN(n1306) );
XNOR2_X1 U1008 ( .A(KEYINPUT59), .B(n1096), .ZN(n1305) );
XOR2_X1 U1009 ( .A(n1308), .B(n1309), .Z(n1303) );
XNOR2_X1 U1010 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR4_X1 U1011 ( .A1(KEYINPUT35), .A2(G953), .A3(G237), .A4(n1312), .ZN(n1311) );
INV_X1 U1012 ( .A(G214), .ZN(n1312) );
NAND2_X1 U1013 ( .A1(KEYINPUT56), .A2(G122), .ZN(n1310) );
XNOR2_X1 U1014 ( .A(n1091), .B(n1313), .ZN(n1308) );
XOR2_X1 U1015 ( .A(G131), .B(G140), .Z(n1091) );
NOR3_X1 U1016 ( .A1(n1048), .A2(n1219), .A3(n1026), .ZN(n1206) );
NAND2_X1 U1017 ( .A1(n1254), .A2(n1025), .ZN(n1026) );
INV_X1 U1018 ( .A(n1071), .ZN(n1025) );
XOR2_X1 U1019 ( .A(n1074), .B(n1075), .Z(n1071) );
INV_X1 U1020 ( .A(G469), .ZN(n1075) );
AND2_X1 U1021 ( .A1(n1314), .A2(n1126), .ZN(n1074) );
XOR2_X1 U1022 ( .A(n1174), .B(n1315), .Z(n1314) );
XOR2_X1 U1023 ( .A(G140), .B(n1316), .Z(n1315) );
NOR2_X1 U1024 ( .A1(KEYINPUT45), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1025 ( .A(n1157), .B(n1318), .Z(n1317) );
XOR2_X1 U1026 ( .A(n1093), .B(n1173), .Z(n1318) );
XNOR2_X1 U1027 ( .A(G101), .B(n1319), .ZN(n1173) );
NAND2_X1 U1028 ( .A1(n1320), .A2(n1321), .ZN(n1093) );
NAND2_X1 U1029 ( .A1(G128), .A2(n1313), .ZN(n1321) );
XOR2_X1 U1030 ( .A(n1322), .B(KEYINPUT36), .Z(n1320) );
NAND2_X1 U1031 ( .A1(n1323), .A2(n1275), .ZN(n1322) );
XNOR2_X1 U1032 ( .A(n1324), .B(n1325), .ZN(n1157) );
INV_X1 U1033 ( .A(n1092), .ZN(n1325) );
XNOR2_X1 U1034 ( .A(G134), .B(G137), .ZN(n1092) );
INV_X1 U1035 ( .A(G131), .ZN(n1324) );
XNOR2_X1 U1036 ( .A(G110), .B(n1326), .ZN(n1174) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1079), .ZN(n1326) );
INV_X1 U1038 ( .A(G227), .ZN(n1079) );
XNOR2_X1 U1039 ( .A(n1024), .B(KEYINPUT7), .ZN(n1254) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1327), .ZN(n1024) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1126), .ZN(n1327) );
INV_X1 U1042 ( .A(n1253), .ZN(n1219) );
NAND2_X1 U1043 ( .A1(n1035), .A2(n1328), .ZN(n1253) );
NAND4_X1 U1044 ( .A1(G953), .A2(G902), .A3(n1249), .A4(n1105), .ZN(n1328) );
INV_X1 U1045 ( .A(G898), .ZN(n1105) );
NAND3_X1 U1046 ( .A1(n1249), .A2(n1031), .A3(G952), .ZN(n1035) );
NAND2_X1 U1047 ( .A1(G237), .A2(G234), .ZN(n1249) );
INV_X1 U1048 ( .A(n1218), .ZN(n1048) );
NOR2_X1 U1049 ( .A1(n1051), .A2(n1050), .ZN(n1218) );
INV_X1 U1050 ( .A(n1235), .ZN(n1050) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1329), .ZN(n1235) );
XNOR2_X1 U1052 ( .A(n1330), .B(n1182), .ZN(n1051) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1329), .ZN(n1182) );
NAND2_X1 U1054 ( .A1(n1287), .A2(n1126), .ZN(n1329) );
INV_X1 U1055 ( .A(G237), .ZN(n1287) );
NAND2_X1 U1056 ( .A1(n1331), .A2(n1126), .ZN(n1330) );
INV_X1 U1057 ( .A(G902), .ZN(n1126) );
XNOR2_X1 U1058 ( .A(n1332), .B(n1333), .ZN(n1331) );
XOR2_X1 U1059 ( .A(KEYINPUT13), .B(n1334), .Z(n1333) );
NOR2_X1 U1060 ( .A1(KEYINPUT48), .A2(n1163), .ZN(n1334) );
NAND2_X1 U1061 ( .A1(n1335), .A2(n1336), .ZN(n1163) );
NAND2_X1 U1062 ( .A1(n1323), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1063 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND2_X1 U1064 ( .A1(G128), .A2(n1340), .ZN(n1339) );
INV_X1 U1065 ( .A(n1313), .ZN(n1323) );
NAND2_X1 U1066 ( .A1(n1341), .A2(n1275), .ZN(n1335) );
INV_X1 U1067 ( .A(G128), .ZN(n1275) );
NAND2_X1 U1068 ( .A1(n1340), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1069 ( .A1(n1313), .A2(n1338), .ZN(n1342) );
INV_X1 U1070 ( .A(KEYINPUT58), .ZN(n1338) );
XOR2_X1 U1071 ( .A(G143), .B(G146), .Z(n1313) );
INV_X1 U1072 ( .A(KEYINPUT34), .ZN(n1340) );
INV_X1 U1073 ( .A(n1179), .ZN(n1332) );
XNOR2_X1 U1074 ( .A(n1343), .B(n1344), .ZN(n1179) );
XNOR2_X1 U1075 ( .A(n1096), .B(n1345), .ZN(n1344) );
NOR2_X1 U1076 ( .A1(KEYINPUT6), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1077 ( .A(n1347), .B(n1115), .ZN(n1346) );
NAND3_X1 U1078 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1115) );
NAND2_X1 U1079 ( .A1(n1319), .A2(n1351), .ZN(n1350) );
NAND2_X1 U1080 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1081 ( .A(KEYINPUT22), .ZN(n1353) );
XNOR2_X1 U1082 ( .A(KEYINPUT38), .B(n1245), .ZN(n1352) );
INV_X1 U1083 ( .A(G101), .ZN(n1245) );
OR3_X1 U1084 ( .A1(n1319), .A2(G101), .A3(KEYINPUT22), .ZN(n1349) );
XOR2_X1 U1085 ( .A(G104), .B(G107), .Z(n1319) );
NAND2_X1 U1086 ( .A1(KEYINPUT22), .A2(G101), .ZN(n1348) );
NAND2_X1 U1087 ( .A1(KEYINPUT3), .A2(n1116), .ZN(n1347) );
XOR2_X1 U1088 ( .A(n1280), .B(n1354), .Z(n1116) );
NOR2_X1 U1089 ( .A1(KEYINPUT39), .A2(n1307), .ZN(n1354) );
INV_X1 U1090 ( .A(G113), .ZN(n1307) );
XNOR2_X1 U1091 ( .A(G116), .B(G119), .ZN(n1280) );
INV_X1 U1092 ( .A(G125), .ZN(n1096) );
XNOR2_X1 U1093 ( .A(n1111), .B(n1355), .ZN(n1343) );
AND2_X1 U1094 ( .A1(n1031), .A2(G224), .ZN(n1355) );
INV_X1 U1095 ( .A(G953), .ZN(n1031) );
XNOR2_X1 U1096 ( .A(n1356), .B(G122), .ZN(n1111) );
NAND2_X1 U1097 ( .A1(KEYINPUT25), .A2(n1357), .ZN(n1356) );
INV_X1 U1098 ( .A(G110), .ZN(n1357) );
endmodule


