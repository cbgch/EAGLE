//Key = 0111100000110010100111100101001101110100011110111100011010101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274;

XNOR2_X1 U702 ( .A(G107), .B(n976), .ZN(G9) );
NOR2_X1 U703 ( .A1(n977), .A2(n978), .ZN(G75) );
NOR3_X1 U704 ( .A1(n979), .A2(n980), .A3(n981), .ZN(n978) );
NOR3_X1 U705 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n980) );
NOR4_X1 U706 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n984) );
XOR2_X1 U707 ( .A(KEYINPUT51), .B(n989), .Z(n988) );
NOR4_X1 U708 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n989) );
XOR2_X1 U709 ( .A(n994), .B(KEYINPUT25), .Z(n987) );
NAND2_X1 U710 ( .A1(n995), .A2(n996), .ZN(n994) );
AND3_X1 U711 ( .A1(n997), .A2(n995), .A3(n998), .ZN(n986) );
NOR3_X1 U712 ( .A1(n993), .A2(n999), .A3(n992), .ZN(n985) );
NOR2_X1 U713 ( .A1(n1000), .A2(n1001), .ZN(n999) );
AND2_X1 U714 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U715 ( .A1(n1004), .A2(n1005), .ZN(n1000) );
NOR2_X1 U716 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NAND3_X1 U717 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n979) );
NAND3_X1 U718 ( .A1(n1011), .A2(n1012), .A3(n995), .ZN(n1010) );
NOR3_X1 U719 ( .A1(n1005), .A2(n990), .A3(n993), .ZN(n995) );
NAND2_X1 U720 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U721 ( .A1(n983), .A2(n1015), .ZN(n1014) );
NOR3_X1 U722 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n977) );
INV_X1 U723 ( .A(n1008), .ZN(n1016) );
NAND4_X1 U724 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1008) );
NOR4_X1 U725 ( .A1(n997), .A2(n983), .A3(n1021), .A4(n1022), .ZN(n1020) );
XOR2_X1 U726 ( .A(n1023), .B(n1024), .Z(n1022) );
XOR2_X1 U727 ( .A(KEYINPUT7), .B(G469), .Z(n1024) );
NAND2_X1 U728 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
XNOR2_X1 U729 ( .A(KEYINPUT16), .B(KEYINPUT1), .ZN(n1025) );
XOR2_X1 U730 ( .A(n1027), .B(n1028), .Z(n1021) );
NAND2_X1 U731 ( .A1(KEYINPUT44), .A2(n1029), .ZN(n1027) );
INV_X1 U732 ( .A(n1030), .ZN(n983) );
NOR2_X1 U733 ( .A1(n1031), .A2(n1032), .ZN(n1019) );
XOR2_X1 U734 ( .A(n1033), .B(n1034), .Z(n1032) );
XOR2_X1 U735 ( .A(n1035), .B(n1036), .Z(n1018) );
XOR2_X1 U736 ( .A(n1037), .B(KEYINPUT26), .Z(n1017) );
NAND2_X1 U737 ( .A1(n1038), .A2(n1039), .ZN(G72) );
NAND2_X1 U738 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XOR2_X1 U739 ( .A(KEYINPUT24), .B(n1042), .Z(n1041) );
XOR2_X1 U740 ( .A(KEYINPUT49), .B(n1043), .Z(n1038) );
NOR2_X1 U741 ( .A1(n1042), .A2(n1040), .ZN(n1043) );
AND2_X1 U742 ( .A1(G953), .A2(n1044), .ZN(n1040) );
NAND2_X1 U743 ( .A1(G900), .A2(G227), .ZN(n1044) );
AND2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1042) );
NAND3_X1 U745 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U746 ( .A1(G953), .A2(n1050), .ZN(n1047) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NAND2_X1 U748 ( .A1(n1049), .A2(n1009), .ZN(n1052) );
XNOR2_X1 U749 ( .A(n1053), .B(n1054), .ZN(n1049) );
XOR2_X1 U750 ( .A(n1055), .B(n1056), .Z(n1054) );
XOR2_X1 U751 ( .A(G140), .B(n1057), .Z(n1056) );
NOR2_X1 U752 ( .A1(G131), .A2(KEYINPUT61), .ZN(n1057) );
NOR2_X1 U753 ( .A1(KEYINPUT40), .A2(n1058), .ZN(n1055) );
INV_X1 U754 ( .A(G125), .ZN(n1058) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(n1053) );
XNOR2_X1 U756 ( .A(KEYINPUT57), .B(n1048), .ZN(n1051) );
NAND2_X1 U757 ( .A1(n1009), .A2(n1061), .ZN(n1048) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XNOR2_X1 U759 ( .A(KEYINPUT41), .B(n1064), .ZN(n1063) );
XOR2_X1 U760 ( .A(n1065), .B(n1066), .Z(G69) );
NOR2_X1 U761 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR3_X1 U762 ( .A1(n1009), .A2(n1069), .A3(n1070), .ZN(n1068) );
XNOR2_X1 U763 ( .A(G898), .B(KEYINPUT0), .ZN(n1069) );
NOR3_X1 U764 ( .A1(G953), .A2(n1071), .A3(n1072), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
XOR2_X1 U766 ( .A(n1075), .B(n1076), .Z(n1074) );
XOR2_X1 U767 ( .A(G122), .B(G110), .Z(n1076) );
NAND2_X1 U768 ( .A1(KEYINPUT37), .A2(n1077), .ZN(n1075) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U770 ( .A1(KEYINPUT13), .A2(n1080), .ZN(n1078) );
NOR2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(G66) );
XOR2_X1 U772 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND3_X1 U773 ( .A1(n1085), .A2(n1086), .A3(KEYINPUT34), .ZN(n1083) );
INV_X1 U774 ( .A(n1034), .ZN(n1086) );
NOR2_X1 U775 ( .A1(n1081), .A2(n1087), .ZN(G63) );
NOR3_X1 U776 ( .A1(n1028), .A2(n1088), .A3(n1089), .ZN(n1087) );
AND3_X1 U777 ( .A1(n1090), .A2(G478), .A3(n1085), .ZN(n1089) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
AND2_X1 U779 ( .A1(n981), .A2(G478), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1081), .A2(n1092), .ZN(G60) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1092) );
AND2_X1 U782 ( .A1(G475), .A2(n1085), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(G6) );
NAND2_X1 U784 ( .A1(KEYINPUT19), .A2(n1071), .ZN(n1096) );
NOR2_X1 U785 ( .A1(n1081), .A2(n1097), .ZN(G57) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U787 ( .A1(n1085), .A2(G472), .A3(KEYINPUT53), .ZN(n1098) );
NOR2_X1 U788 ( .A1(n1081), .A2(n1100), .ZN(G54) );
XOR2_X1 U789 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U790 ( .A(n1060), .B(n1103), .ZN(n1102) );
XOR2_X1 U791 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1101) );
XOR2_X1 U793 ( .A(n1108), .B(n1109), .Z(n1107) );
AND2_X1 U794 ( .A1(G469), .A2(n1085), .ZN(n1108) );
INV_X1 U795 ( .A(n1110), .ZN(n1085) );
XNOR2_X1 U796 ( .A(KEYINPUT52), .B(KEYINPUT23), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1081), .A2(n1111), .ZN(G51) );
XOR2_X1 U798 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR3_X1 U800 ( .A1(n1110), .A2(KEYINPUT63), .A3(n1116), .ZN(n1114) );
NAND2_X1 U801 ( .A1(G902), .A2(n981), .ZN(n1110) );
NAND4_X1 U802 ( .A1(n1062), .A2(n1117), .A3(n1118), .A4(n1064), .ZN(n981) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1064) );
XNOR2_X1 U804 ( .A(KEYINPUT15), .B(n1121), .ZN(n1120) );
XOR2_X1 U805 ( .A(KEYINPUT2), .B(n1071), .Z(n1118) );
AND3_X1 U806 ( .A1(n1122), .A2(n1003), .A3(n1123), .ZN(n1071) );
INV_X1 U807 ( .A(n1072), .ZN(n1117) );
NAND4_X1 U808 ( .A1(n1124), .A2(n976), .A3(n1125), .A4(n1126), .ZN(n1072) );
NOR3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1119), .A2(n1130), .ZN(n1125) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U812 ( .A(KEYINPUT42), .B(n1133), .ZN(n1132) );
XOR2_X1 U813 ( .A(n1134), .B(KEYINPUT50), .Z(n1131) );
NAND3_X1 U814 ( .A1(n1003), .A2(n1002), .A3(n1122), .ZN(n976) );
AND4_X1 U815 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1062) );
NOR4_X1 U816 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1138) );
INV_X1 U817 ( .A(n1143), .ZN(n1142) );
XNOR2_X1 U818 ( .A(KEYINPUT5), .B(KEYINPUT32), .ZN(n1112) );
NOR2_X1 U819 ( .A1(n1009), .A2(G952), .ZN(n1081) );
XNOR2_X1 U820 ( .A(n1137), .B(n1144), .ZN(G48) );
NOR2_X1 U821 ( .A1(KEYINPUT17), .A2(n1145), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1123), .A2(n1146), .ZN(n1137) );
XOR2_X1 U823 ( .A(n1147), .B(n1135), .Z(G45) );
NAND4_X1 U824 ( .A1(n1148), .A2(n1007), .A3(n1149), .A4(n1031), .ZN(n1135) );
INV_X1 U825 ( .A(n1150), .ZN(n1149) );
XNOR2_X1 U826 ( .A(G140), .B(n1136), .ZN(G42) );
NAND3_X1 U827 ( .A1(n1123), .A2(n1151), .A3(n1006), .ZN(n1136) );
XOR2_X1 U828 ( .A(n1152), .B(n1140), .Z(G39) );
AND4_X1 U829 ( .A1(n1153), .A2(n1151), .A3(n1154), .A4(n1155), .ZN(n1140) );
XNOR2_X1 U830 ( .A(G137), .B(KEYINPUT58), .ZN(n1152) );
XNOR2_X1 U831 ( .A(G134), .B(n1156), .ZN(G36) );
NAND2_X1 U832 ( .A1(KEYINPUT11), .A2(n1139), .ZN(n1156) );
AND3_X1 U833 ( .A1(n1151), .A2(n1002), .A3(n1007), .ZN(n1139) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(G33) );
NOR2_X1 U835 ( .A1(KEYINPUT62), .A2(n1143), .ZN(n1158) );
NAND3_X1 U836 ( .A1(n1007), .A2(n1151), .A3(n1123), .ZN(n1143) );
AND4_X1 U837 ( .A1(n996), .A2(n1015), .A3(n1159), .A4(n1030), .ZN(n1151) );
INV_X1 U838 ( .A(n982), .ZN(n1015) );
XOR2_X1 U839 ( .A(n1160), .B(KEYINPUT21), .Z(n1157) );
XOR2_X1 U840 ( .A(G128), .B(n1141), .Z(G30) );
AND2_X1 U841 ( .A1(n1146), .A2(n1002), .ZN(n1141) );
AND3_X1 U842 ( .A1(n1154), .A2(n1155), .A3(n1148), .ZN(n1146) );
AND3_X1 U843 ( .A1(n1119), .A2(n1159), .A3(n996), .ZN(n1148) );
INV_X1 U844 ( .A(n1161), .ZN(n1155) );
XOR2_X1 U845 ( .A(G101), .B(n1162), .Z(G3) );
NOR3_X1 U846 ( .A1(KEYINPUT9), .A2(n1163), .A3(n1164), .ZN(n1162) );
NOR2_X1 U847 ( .A1(KEYINPUT48), .A2(n1165), .ZN(n1164) );
NOR3_X1 U848 ( .A1(n1166), .A2(n1167), .A3(n1005), .ZN(n1165) );
NAND3_X1 U849 ( .A1(n1168), .A2(n1169), .A3(n1119), .ZN(n1166) );
INV_X1 U850 ( .A(n1013), .ZN(n1119) );
NOR2_X1 U851 ( .A1(n1127), .A2(n1170), .ZN(n1163) );
INV_X1 U852 ( .A(KEYINPUT48), .ZN(n1170) );
AND3_X1 U853 ( .A1(n1007), .A2(n1122), .A3(n1153), .ZN(n1127) );
INV_X1 U854 ( .A(n1167), .ZN(n1007) );
XOR2_X1 U855 ( .A(G125), .B(n1171), .Z(G27) );
NOR2_X1 U856 ( .A1(n1013), .A2(n1121), .ZN(n1171) );
NAND4_X1 U857 ( .A1(n1011), .A2(n1006), .A3(n1123), .A4(n1159), .ZN(n1121) );
NAND2_X1 U858 ( .A1(n993), .A2(n1172), .ZN(n1159) );
NAND4_X1 U859 ( .A1(G902), .A2(G953), .A3(n1173), .A4(n1050), .ZN(n1172) );
INV_X1 U860 ( .A(G900), .ZN(n1050) );
XOR2_X1 U861 ( .A(G122), .B(n1174), .Z(G24) );
NOR2_X1 U862 ( .A1(n1013), .A2(n1134), .ZN(n1174) );
NAND3_X1 U863 ( .A1(n1011), .A2(n1003), .A3(n1175), .ZN(n1134) );
NOR3_X1 U864 ( .A1(n1150), .A2(n1176), .A3(n1177), .ZN(n1175) );
INV_X1 U865 ( .A(n990), .ZN(n1003) );
NAND2_X1 U866 ( .A1(n1161), .A2(n1037), .ZN(n990) );
XOR2_X1 U867 ( .A(G119), .B(n1178), .Z(G21) );
NOR2_X1 U868 ( .A1(n1013), .A2(n1133), .ZN(n1178) );
NAND3_X1 U869 ( .A1(n1011), .A2(n1153), .A3(n1179), .ZN(n1133) );
NOR3_X1 U870 ( .A1(n1037), .A2(n1176), .A3(n1161), .ZN(n1179) );
INV_X1 U871 ( .A(n992), .ZN(n1011) );
XOR2_X1 U872 ( .A(G116), .B(n1129), .Z(G18) );
AND2_X1 U873 ( .A1(n1180), .A2(n1002), .ZN(n1129) );
NOR2_X1 U874 ( .A1(n1031), .A2(n1150), .ZN(n1002) );
XOR2_X1 U875 ( .A(G113), .B(n1128), .Z(G15) );
AND2_X1 U876 ( .A1(n1180), .A2(n1123), .ZN(n1128) );
INV_X1 U877 ( .A(n991), .ZN(n1123) );
NAND2_X1 U878 ( .A1(n1150), .A2(n1031), .ZN(n991) );
INV_X1 U879 ( .A(n1177), .ZN(n1031) );
NOR4_X1 U880 ( .A1(n992), .A2(n1167), .A3(n1013), .A4(n1176), .ZN(n1180) );
NAND2_X1 U881 ( .A1(n1161), .A2(n1154), .ZN(n1167) );
NAND2_X1 U882 ( .A1(n998), .A2(n1181), .ZN(n992) );
XOR2_X1 U883 ( .A(n1182), .B(n1124), .Z(G12) );
NAND3_X1 U884 ( .A1(n1153), .A2(n1122), .A3(n1006), .ZN(n1124) );
NOR2_X1 U885 ( .A1(n1154), .A2(n1161), .ZN(n1006) );
XOR2_X1 U886 ( .A(n1033), .B(n1183), .Z(n1161) );
NOR2_X1 U887 ( .A1(KEYINPUT29), .A2(n1034), .ZN(n1183) );
NAND2_X1 U888 ( .A1(G217), .A2(n1184), .ZN(n1034) );
NAND2_X1 U889 ( .A1(n1084), .A2(n1185), .ZN(n1033) );
XOR2_X1 U890 ( .A(KEYINPUT14), .B(G902), .Z(n1185) );
XOR2_X1 U891 ( .A(n1186), .B(n1187), .Z(n1084) );
XOR2_X1 U892 ( .A(KEYINPUT33), .B(G137), .Z(n1187) );
XNOR2_X1 U893 ( .A(n1188), .B(n1189), .ZN(n1186) );
NOR2_X1 U894 ( .A1(KEYINPUT45), .A2(n1190), .ZN(n1189) );
XOR2_X1 U895 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U896 ( .A(G146), .B(G140), .Z(n1192) );
XOR2_X1 U897 ( .A(n1193), .B(n1194), .Z(n1191) );
NAND2_X1 U898 ( .A1(KEYINPUT56), .A2(n1195), .ZN(n1193) );
XOR2_X1 U899 ( .A(G128), .B(G119), .Z(n1195) );
NOR4_X1 U900 ( .A1(KEYINPUT6), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1188) );
INV_X1 U901 ( .A(G221), .ZN(n1198) );
INV_X1 U902 ( .A(G234), .ZN(n1197) );
XOR2_X1 U903 ( .A(n1009), .B(KEYINPUT4), .Z(n1196) );
INV_X1 U904 ( .A(n1037), .ZN(n1154) );
XOR2_X1 U905 ( .A(n1199), .B(G472), .Z(n1037) );
NAND2_X1 U906 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U907 ( .A(n1099), .B(KEYINPUT28), .Z(n1200) );
XOR2_X1 U908 ( .A(n1202), .B(n1203), .Z(n1099) );
XNOR2_X1 U909 ( .A(n1080), .B(n1204), .ZN(n1203) );
XOR2_X1 U910 ( .A(G101), .B(n1205), .Z(n1204) );
AND3_X1 U911 ( .A1(G210), .A2(n1009), .A3(n1206), .ZN(n1205) );
XOR2_X1 U912 ( .A(n1207), .B(n1208), .Z(n1202) );
NOR3_X1 U913 ( .A1(n1013), .A2(n1176), .A3(n1169), .ZN(n1122) );
INV_X1 U914 ( .A(n996), .ZN(n1169) );
NOR2_X1 U915 ( .A1(n998), .A2(n997), .ZN(n996) );
INV_X1 U916 ( .A(n1181), .ZN(n997) );
NAND2_X1 U917 ( .A1(G221), .A2(n1184), .ZN(n1181) );
NAND2_X1 U918 ( .A1(G234), .A2(n1201), .ZN(n1184) );
XOR2_X1 U919 ( .A(n1026), .B(G469), .Z(n998) );
NAND2_X1 U920 ( .A1(n1209), .A2(n1201), .ZN(n1026) );
XNOR2_X1 U921 ( .A(n1210), .B(n1109), .ZN(n1209) );
XNOR2_X1 U922 ( .A(n1211), .B(n1212), .ZN(n1109) );
XOR2_X1 U923 ( .A(G140), .B(G110), .Z(n1212) );
NAND2_X1 U924 ( .A1(G227), .A2(n1009), .ZN(n1211) );
NAND2_X1 U925 ( .A1(n1213), .A2(KEYINPUT46), .ZN(n1210) );
XOR2_X1 U926 ( .A(n1214), .B(n1104), .Z(n1213) );
XNOR2_X1 U927 ( .A(n1207), .B(KEYINPUT30), .ZN(n1104) );
XOR2_X1 U928 ( .A(n1215), .B(n1059), .Z(n1207) );
XOR2_X1 U929 ( .A(G137), .B(G134), .Z(n1059) );
XOR2_X1 U930 ( .A(n1160), .B(KEYINPUT55), .Z(n1215) );
INV_X1 U931 ( .A(G131), .ZN(n1160) );
NAND2_X1 U932 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND2_X1 U933 ( .A1(n1060), .A2(n1105), .ZN(n1217) );
XOR2_X1 U934 ( .A(KEYINPUT22), .B(n1218), .Z(n1216) );
NOR2_X1 U935 ( .A1(n1060), .A2(n1105), .ZN(n1218) );
XNOR2_X1 U936 ( .A(n1219), .B(n1220), .ZN(n1105) );
NAND2_X1 U937 ( .A1(KEYINPUT10), .A2(n1095), .ZN(n1219) );
XOR2_X1 U938 ( .A(n1221), .B(n1222), .Z(n1060) );
XOR2_X1 U939 ( .A(n1145), .B(G143), .Z(n1221) );
INV_X1 U940 ( .A(n1168), .ZN(n1176) );
NAND2_X1 U941 ( .A1(n993), .A2(n1223), .ZN(n1168) );
NAND3_X1 U942 ( .A1(n1073), .A2(n1173), .A3(G902), .ZN(n1223) );
NOR2_X1 U943 ( .A1(n1009), .A2(G898), .ZN(n1073) );
NAND3_X1 U944 ( .A1(n1173), .A2(n1009), .A3(G952), .ZN(n993) );
NAND2_X1 U945 ( .A1(G237), .A2(n1224), .ZN(n1173) );
XOR2_X1 U946 ( .A(KEYINPUT12), .B(G234), .Z(n1224) );
NAND2_X1 U947 ( .A1(n982), .A2(n1030), .ZN(n1013) );
NAND2_X1 U948 ( .A1(G214), .A2(n1225), .ZN(n1030) );
XOR2_X1 U949 ( .A(n1035), .B(n1226), .Z(n982) );
NOR2_X1 U950 ( .A1(n1036), .A2(KEYINPUT36), .ZN(n1226) );
INV_X1 U951 ( .A(n1116), .ZN(n1036) );
NAND2_X1 U952 ( .A1(G210), .A2(n1225), .ZN(n1116) );
NAND2_X1 U953 ( .A1(n1206), .A2(n1201), .ZN(n1225) );
NAND2_X1 U954 ( .A1(n1115), .A2(n1201), .ZN(n1035) );
INV_X1 U955 ( .A(G902), .ZN(n1201) );
XNOR2_X1 U956 ( .A(n1227), .B(n1228), .ZN(n1115) );
XNOR2_X1 U957 ( .A(n1080), .B(n1229), .ZN(n1228) );
XOR2_X1 U958 ( .A(G122), .B(n1230), .Z(n1229) );
NOR2_X1 U959 ( .A1(G953), .A2(n1070), .ZN(n1230) );
INV_X1 U960 ( .A(G224), .ZN(n1070) );
XNOR2_X1 U961 ( .A(G113), .B(n1231), .ZN(n1080) );
XOR2_X1 U962 ( .A(G119), .B(G116), .Z(n1231) );
XOR2_X1 U963 ( .A(n1232), .B(n1079), .Z(n1227) );
XNOR2_X1 U964 ( .A(n1233), .B(n1220), .ZN(n1079) );
XOR2_X1 U965 ( .A(G101), .B(G107), .Z(n1220) );
NAND2_X1 U966 ( .A1(KEYINPUT54), .A2(n1095), .ZN(n1233) );
XNOR2_X1 U967 ( .A(n1194), .B(n1208), .ZN(n1232) );
XNOR2_X1 U968 ( .A(n1234), .B(n1222), .ZN(n1208) );
XOR2_X1 U969 ( .A(G128), .B(KEYINPUT39), .Z(n1222) );
NAND3_X1 U970 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1234) );
NAND2_X1 U971 ( .A1(KEYINPUT59), .A2(G143), .ZN(n1237) );
NAND3_X1 U972 ( .A1(n1147), .A2(n1238), .A3(G146), .ZN(n1236) );
NAND2_X1 U973 ( .A1(n1239), .A2(n1145), .ZN(n1235) );
NAND2_X1 U974 ( .A1(n1240), .A2(n1238), .ZN(n1239) );
INV_X1 U975 ( .A(KEYINPUT59), .ZN(n1238) );
XOR2_X1 U976 ( .A(KEYINPUT20), .B(G143), .Z(n1240) );
XNOR2_X1 U977 ( .A(n1182), .B(G125), .ZN(n1194) );
INV_X1 U978 ( .A(n1005), .ZN(n1153) );
NAND2_X1 U979 ( .A1(n1150), .A2(n1177), .ZN(n1005) );
XOR2_X1 U980 ( .A(n1241), .B(G475), .Z(n1177) );
OR2_X1 U981 ( .A1(n1094), .A2(G902), .ZN(n1241) );
XNOR2_X1 U982 ( .A(n1242), .B(n1243), .ZN(n1094) );
XOR2_X1 U983 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U984 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U985 ( .A1(n1248), .A2(n1147), .ZN(n1247) );
XOR2_X1 U986 ( .A(n1249), .B(KEYINPUT38), .Z(n1246) );
OR2_X1 U987 ( .A1(n1248), .A2(n1147), .ZN(n1249) );
INV_X1 U988 ( .A(G143), .ZN(n1147) );
NAND3_X1 U989 ( .A1(n1206), .A2(n1009), .A3(G214), .ZN(n1248) );
INV_X1 U990 ( .A(G237), .ZN(n1206) );
NAND2_X1 U991 ( .A1(KEYINPUT43), .A2(n1250), .ZN(n1244) );
XOR2_X1 U992 ( .A(n1145), .B(n1251), .Z(n1250) );
NAND2_X1 U993 ( .A1(KEYINPUT35), .A2(n1252), .ZN(n1251) );
XOR2_X1 U994 ( .A(G140), .B(G125), .Z(n1252) );
INV_X1 U995 ( .A(G146), .ZN(n1145) );
XOR2_X1 U996 ( .A(n1253), .B(G131), .Z(n1242) );
NAND3_X1 U997 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1253) );
OR2_X1 U998 ( .A1(n1095), .A2(KEYINPUT31), .ZN(n1256) );
NAND3_X1 U999 ( .A1(KEYINPUT31), .A2(n1257), .A3(n1258), .ZN(n1255) );
OR2_X1 U1000 ( .A1(n1258), .A2(n1257), .ZN(n1254) );
AND2_X1 U1001 ( .A1(KEYINPUT60), .A2(n1095), .ZN(n1257) );
INV_X1 U1002 ( .A(G104), .ZN(n1095) );
XOR2_X1 U1003 ( .A(G113), .B(G122), .Z(n1258) );
XOR2_X1 U1004 ( .A(n1029), .B(n1028), .Z(n1150) );
NOR2_X1 U1005 ( .A1(n1090), .A2(G902), .ZN(n1028) );
AND2_X1 U1006 ( .A1(n1259), .A2(n1260), .ZN(n1090) );
NAND2_X1 U1007 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U1008 ( .A(KEYINPUT3), .B(n1263), .Z(n1259) );
NOR2_X1 U1009 ( .A1(n1262), .A2(n1261), .ZN(n1263) );
AND2_X1 U1010 ( .A1(n1264), .A2(n1265), .ZN(n1261) );
NAND2_X1 U1011 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n1268), .Z(n1264) );
NOR2_X1 U1013 ( .A1(n1266), .A2(n1267), .ZN(n1268) );
NAND2_X1 U1014 ( .A1(n1269), .A2(n1270), .ZN(n1267) );
OR2_X1 U1015 ( .A1(n1271), .A2(G134), .ZN(n1270) );
XOR2_X1 U1016 ( .A(n1272), .B(KEYINPUT8), .Z(n1269) );
NAND2_X1 U1017 ( .A1(G134), .A2(n1271), .ZN(n1272) );
XOR2_X1 U1018 ( .A(G128), .B(G143), .Z(n1271) );
XNOR2_X1 U1019 ( .A(n1273), .B(G107), .ZN(n1266) );
NAND2_X1 U1020 ( .A1(KEYINPUT27), .A2(n1274), .ZN(n1273) );
XOR2_X1 U1021 ( .A(G122), .B(G116), .Z(n1274) );
AND3_X1 U1022 ( .A1(G234), .A2(n1009), .A3(G217), .ZN(n1262) );
INV_X1 U1023 ( .A(G953), .ZN(n1009) );
XNOR2_X1 U1024 ( .A(G478), .B(KEYINPUT18), .ZN(n1029) );
INV_X1 U1025 ( .A(G110), .ZN(n1182) );
endmodule


