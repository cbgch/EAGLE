//Key = 0111101110011011101010000000010000000000011110111010101010011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331;

XOR2_X1 U738 ( .A(n1011), .B(n1012), .Z(G9) );
NOR2_X1 U739 ( .A1(G107), .A2(KEYINPUT53), .ZN(n1012) );
NOR2_X1 U740 ( .A1(n1013), .A2(n1014), .ZN(G75) );
XOR2_X1 U741 ( .A(n1015), .B(KEYINPUT60), .Z(n1014) );
NAND3_X1 U742 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NAND2_X1 U743 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U744 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NAND3_X1 U745 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U746 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
OR2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U749 ( .A1(n1032), .A2(n1033), .ZN(n1026) );
NAND2_X1 U750 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U751 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U752 ( .A1(n1032), .A2(n1038), .A3(n1028), .ZN(n1021) );
NAND2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U754 ( .A1(n1025), .A2(n1041), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1023), .A2(n1044), .ZN(n1039) );
NAND2_X1 U757 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U758 ( .A1(G214), .A2(n1047), .A3(n1048), .ZN(n1046) );
INV_X1 U759 ( .A(n1049), .ZN(n1016) );
NOR2_X1 U760 ( .A1(G952), .A2(n1049), .ZN(n1013) );
NAND2_X1 U761 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND4_X1 U762 ( .A1(n1037), .A2(n1052), .A3(n1025), .A4(n1053), .ZN(n1051) );
NOR4_X1 U763 ( .A1(n1036), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1053) );
XNOR2_X1 U764 ( .A(G475), .B(n1057), .ZN(n1056) );
NOR2_X1 U765 ( .A1(n1058), .A2(KEYINPUT40), .ZN(n1057) );
XOR2_X1 U766 ( .A(n1059), .B(G472), .Z(n1055) );
NAND2_X1 U767 ( .A1(KEYINPUT46), .A2(n1060), .ZN(n1059) );
XNOR2_X1 U768 ( .A(n1061), .B(n1062), .ZN(n1054) );
XOR2_X1 U769 ( .A(n1063), .B(n1064), .Z(G72) );
NOR2_X1 U770 ( .A1(n1065), .A2(n1050), .ZN(n1064) );
AND2_X1 U771 ( .A1(G227), .A2(G900), .ZN(n1065) );
NAND2_X1 U772 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NAND3_X1 U773 ( .A1(n1068), .A2(n1050), .A3(n1069), .ZN(n1067) );
XOR2_X1 U774 ( .A(n1070), .B(KEYINPUT36), .Z(n1066) );
NAND2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U776 ( .A1(n1068), .A2(n1050), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1069), .B(KEYINPUT63), .Z(n1071) );
NAND2_X1 U778 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
XOR2_X1 U779 ( .A(n1075), .B(n1076), .Z(n1074) );
XOR2_X1 U780 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U781 ( .A(n1079), .B(n1080), .Z(n1075) );
XNOR2_X1 U782 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR3_X1 U783 ( .A1(KEYINPUT19), .A2(n1083), .A3(n1084), .ZN(n1082) );
NOR2_X1 U784 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U785 ( .A(KEYINPUT43), .ZN(n1085) );
NOR2_X1 U786 ( .A1(KEYINPUT43), .A2(n1087), .ZN(n1083) );
NOR2_X1 U787 ( .A1(G137), .A2(n1088), .ZN(n1087) );
NAND2_X1 U788 ( .A1(KEYINPUT2), .A2(n1089), .ZN(n1081) );
XOR2_X1 U789 ( .A(n1090), .B(KEYINPUT30), .Z(n1073) );
NAND2_X1 U790 ( .A1(G953), .A2(n1091), .ZN(n1090) );
XOR2_X1 U791 ( .A(n1092), .B(n1093), .Z(G69) );
XOR2_X1 U792 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U793 ( .A1(n1096), .A2(G953), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U795 ( .A(KEYINPUT39), .B(n1099), .ZN(n1098) );
NOR2_X1 U796 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
XOR2_X1 U797 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U798 ( .A(G122), .B(n1104), .Z(n1103) );
NAND2_X1 U799 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U801 ( .A(n1109), .ZN(n1108) );
XNOR2_X1 U802 ( .A(n1110), .B(KEYINPUT41), .ZN(n1107) );
NAND2_X1 U803 ( .A1(n1111), .A2(n1109), .ZN(n1105) );
XNOR2_X1 U804 ( .A(KEYINPUT7), .B(n1112), .ZN(n1111) );
INV_X1 U805 ( .A(n1110), .ZN(n1112) );
XOR2_X1 U806 ( .A(G116), .B(n1113), .Z(n1110) );
NOR2_X1 U807 ( .A1(G898), .A2(n1050), .ZN(n1100) );
NOR2_X1 U808 ( .A1(n1114), .A2(n1050), .ZN(n1092) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U810 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XOR2_X1 U811 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U812 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NOR2_X1 U813 ( .A1(n1117), .A2(n1123), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1061), .A2(n1124), .A3(n1125), .ZN(n1123) );
AND3_X1 U815 ( .A1(n1126), .A2(G478), .A3(n1121), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1127), .A2(n1126), .ZN(n1124) );
AND2_X1 U817 ( .A1(n1128), .A2(G478), .ZN(n1127) );
NOR2_X1 U818 ( .A1(n1117), .A2(n1129), .ZN(G60) );
XOR2_X1 U819 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U820 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1130) );
NAND2_X1 U821 ( .A1(n1121), .A2(G475), .ZN(n1132) );
XNOR2_X1 U822 ( .A(G104), .B(n1099), .ZN(G6) );
NOR2_X1 U823 ( .A1(n1117), .A2(n1133), .ZN(G57) );
XOR2_X1 U824 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U825 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND2_X1 U826 ( .A1(KEYINPUT12), .A2(n1138), .ZN(n1136) );
XOR2_X1 U827 ( .A(n1139), .B(n1140), .Z(n1134) );
NAND2_X1 U828 ( .A1(n1121), .A2(G472), .ZN(n1140) );
NAND2_X1 U829 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND2_X1 U830 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U831 ( .A(n1145), .B(KEYINPUT37), .Z(n1141) );
NAND2_X1 U832 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U833 ( .A(KEYINPUT62), .B(n1143), .Z(n1146) );
XNOR2_X1 U834 ( .A(n1148), .B(KEYINPUT23), .ZN(n1143) );
NOR2_X1 U835 ( .A1(n1117), .A2(n1149), .ZN(G54) );
XOR2_X1 U836 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U837 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U838 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U839 ( .A1(n1121), .A2(G469), .ZN(n1154) );
NOR2_X1 U840 ( .A1(n1156), .A2(n1018), .ZN(n1121) );
XOR2_X1 U841 ( .A(n1157), .B(n1158), .Z(n1150) );
XNOR2_X1 U842 ( .A(G110), .B(G140), .ZN(n1158) );
NAND2_X1 U843 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
XOR2_X1 U844 ( .A(n1078), .B(n1161), .Z(n1160) );
XNOR2_X1 U845 ( .A(G146), .B(n1162), .ZN(n1161) );
XOR2_X1 U846 ( .A(KEYINPUT27), .B(G128), .Z(n1078) );
XNOR2_X1 U847 ( .A(KEYINPUT8), .B(KEYINPUT20), .ZN(n1159) );
NOR2_X1 U848 ( .A1(n1117), .A2(n1163), .ZN(G51) );
NOR2_X1 U849 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U850 ( .A(KEYINPUT35), .B(n1166), .Z(n1165) );
NOR2_X1 U851 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
AND2_X1 U852 ( .A1(n1168), .A2(n1167), .ZN(n1164) );
NAND3_X1 U853 ( .A1(n1169), .A2(n1128), .A3(n1170), .ZN(n1167) );
XNOR2_X1 U854 ( .A(G902), .B(KEYINPUT61), .ZN(n1170) );
INV_X1 U855 ( .A(n1018), .ZN(n1128) );
NOR3_X1 U856 ( .A1(n1068), .A2(n1171), .A3(n1097), .ZN(n1018) );
NAND4_X1 U857 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1097) );
AND4_X1 U858 ( .A1(n1011), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1175) );
NAND3_X1 U859 ( .A1(n1031), .A2(n1023), .A3(n1179), .ZN(n1011) );
NOR2_X1 U860 ( .A1(n1180), .A2(n1181), .ZN(n1174) );
NOR2_X1 U861 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
INV_X1 U862 ( .A(KEYINPUT50), .ZN(n1182) );
NOR2_X1 U863 ( .A1(KEYINPUT50), .A2(n1184), .ZN(n1180) );
NAND4_X1 U864 ( .A1(n1185), .A2(n1186), .A3(n1023), .A4(n1187), .ZN(n1184) );
NOR3_X1 U865 ( .A1(n1188), .A2(n1028), .A3(n1189), .ZN(n1187) );
INV_X1 U866 ( .A(n1099), .ZN(n1171) );
NAND3_X1 U867 ( .A1(n1179), .A2(n1023), .A3(n1030), .ZN(n1099) );
NAND4_X1 U868 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1068) );
NOR4_X1 U869 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
INV_X1 U870 ( .A(n1198), .ZN(n1195) );
NAND2_X1 U871 ( .A1(n1199), .A2(n1200), .ZN(n1192) );
INV_X1 U872 ( .A(KEYINPUT31), .ZN(n1200) );
NAND3_X1 U873 ( .A1(n1201), .A2(n1032), .A3(n1202), .ZN(n1191) );
NAND2_X1 U874 ( .A1(n1030), .A2(n1203), .ZN(n1190) );
NAND3_X1 U875 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NAND2_X1 U876 ( .A1(n1207), .A2(n1201), .ZN(n1206) );
NAND3_X1 U877 ( .A1(n1208), .A2(n1045), .A3(KEYINPUT31), .ZN(n1205) );
NAND2_X1 U878 ( .A1(n1202), .A2(n1209), .ZN(n1204) );
NAND2_X1 U879 ( .A1(n1210), .A2(n1211), .ZN(n1168) );
NAND2_X1 U880 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U881 ( .A(n1214), .B(KEYINPUT55), .Z(n1210) );
OR2_X1 U882 ( .A1(n1212), .A2(n1213), .ZN(n1214) );
XOR2_X1 U883 ( .A(n1215), .B(n1216), .Z(n1212) );
NAND2_X1 U884 ( .A1(KEYINPUT42), .A2(n1217), .ZN(n1215) );
INV_X1 U885 ( .A(n1089), .ZN(n1217) );
NOR2_X1 U886 ( .A1(n1050), .A2(G952), .ZN(n1117) );
XOR2_X1 U887 ( .A(G146), .B(n1218), .Z(G48) );
NOR3_X1 U888 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1218) );
XNOR2_X1 U889 ( .A(n1201), .B(KEYINPUT51), .ZN(n1220) );
XNOR2_X1 U890 ( .A(n1162), .B(n1197), .ZN(G45) );
NOR4_X1 U891 ( .A1(n1219), .A2(n1043), .A3(n1222), .A4(n1188), .ZN(n1197) );
NAND2_X1 U892 ( .A1(n1223), .A2(n1224), .ZN(G42) );
NAND2_X1 U893 ( .A1(G140), .A2(n1225), .ZN(n1224) );
XOR2_X1 U894 ( .A(n1226), .B(KEYINPUT28), .Z(n1223) );
OR2_X1 U895 ( .A1(n1225), .A2(G140), .ZN(n1226) );
INV_X1 U896 ( .A(n1196), .ZN(n1225) );
NOR3_X1 U897 ( .A1(n1042), .A2(n1221), .A3(n1227), .ZN(n1196) );
XOR2_X1 U898 ( .A(G137), .B(n1228), .Z(G39) );
NOR3_X1 U899 ( .A1(n1227), .A2(n1229), .A3(n1230), .ZN(n1228) );
INV_X1 U900 ( .A(n1201), .ZN(n1230) );
XNOR2_X1 U901 ( .A(n1032), .B(KEYINPUT9), .ZN(n1229) );
XNOR2_X1 U902 ( .A(G134), .B(n1198), .ZN(G36) );
NAND3_X1 U903 ( .A1(n1209), .A2(n1031), .A3(n1202), .ZN(n1198) );
XOR2_X1 U904 ( .A(n1231), .B(n1232), .Z(G33) );
XOR2_X1 U905 ( .A(KEYINPUT59), .B(G131), .Z(n1232) );
NAND3_X1 U906 ( .A1(n1202), .A2(n1030), .A3(n1233), .ZN(n1231) );
XNOR2_X1 U907 ( .A(n1209), .B(KEYINPUT11), .ZN(n1233) );
INV_X1 U908 ( .A(n1227), .ZN(n1202) );
NAND3_X1 U909 ( .A1(n1234), .A2(n1235), .A3(n1025), .ZN(n1227) );
AND2_X1 U910 ( .A1(n1048), .A2(n1236), .ZN(n1025) );
INV_X1 U911 ( .A(n1237), .ZN(n1048) );
XOR2_X1 U912 ( .A(G128), .B(n1194), .Z(G30) );
AND3_X1 U913 ( .A1(n1201), .A2(n1031), .A3(n1207), .ZN(n1194) );
INV_X1 U914 ( .A(n1219), .ZN(n1207) );
NAND3_X1 U915 ( .A1(n1234), .A2(n1235), .A3(n1185), .ZN(n1219) );
XNOR2_X1 U916 ( .A(G101), .B(n1172), .ZN(G3) );
NAND3_X1 U917 ( .A1(n1032), .A2(n1179), .A3(n1209), .ZN(n1172) );
XOR2_X1 U918 ( .A(n1238), .B(n1199), .Z(G27) );
AND3_X1 U919 ( .A1(n1185), .A2(n1030), .A3(n1208), .ZN(n1199) );
AND3_X1 U920 ( .A1(n1239), .A2(n1235), .A3(n1028), .ZN(n1208) );
NAND2_X1 U921 ( .A1(n1240), .A2(n1241), .ZN(n1235) );
NAND2_X1 U922 ( .A1(n1242), .A2(n1091), .ZN(n1241) );
INV_X1 U923 ( .A(G900), .ZN(n1091) );
NAND2_X1 U924 ( .A1(KEYINPUT14), .A2(n1243), .ZN(n1238) );
INV_X1 U925 ( .A(G125), .ZN(n1243) );
XOR2_X1 U926 ( .A(n1183), .B(n1244), .Z(G24) );
XNOR2_X1 U927 ( .A(G122), .B(KEYINPUT25), .ZN(n1244) );
NAND4_X1 U928 ( .A1(n1245), .A2(n1246), .A3(n1186), .A4(n1023), .ZN(n1183) );
AND2_X1 U929 ( .A1(n1052), .A2(n1247), .ZN(n1023) );
XNOR2_X1 U930 ( .A(G119), .B(n1173), .ZN(G21) );
NAND3_X1 U931 ( .A1(n1246), .A2(n1032), .A3(n1201), .ZN(n1173) );
NOR2_X1 U932 ( .A1(n1248), .A2(n1052), .ZN(n1201) );
XOR2_X1 U933 ( .A(KEYINPUT45), .B(n1247), .Z(n1248) );
XNOR2_X1 U934 ( .A(G116), .B(n1178), .ZN(G18) );
NAND3_X1 U935 ( .A1(n1209), .A2(n1031), .A3(n1246), .ZN(n1178) );
AND3_X1 U936 ( .A1(n1028), .A2(n1249), .A3(n1185), .ZN(n1246) );
INV_X1 U937 ( .A(n1045), .ZN(n1185) );
XNOR2_X1 U938 ( .A(n1250), .B(KEYINPUT6), .ZN(n1045) );
NOR2_X1 U939 ( .A1(n1222), .A2(n1245), .ZN(n1031) );
XOR2_X1 U940 ( .A(n1251), .B(G113), .Z(G15) );
NAND2_X1 U941 ( .A1(KEYINPUT56), .A2(n1177), .ZN(n1251) );
NAND3_X1 U942 ( .A1(n1028), .A2(n1209), .A3(n1252), .ZN(n1177) );
NOR3_X1 U943 ( .A1(n1221), .A2(n1189), .A3(n1250), .ZN(n1252) );
INV_X1 U944 ( .A(n1030), .ZN(n1221) );
NOR2_X1 U945 ( .A1(n1188), .A2(n1186), .ZN(n1030) );
INV_X1 U946 ( .A(n1043), .ZN(n1209) );
NAND2_X1 U947 ( .A1(n1052), .A2(n1253), .ZN(n1043) );
XNOR2_X1 U948 ( .A(KEYINPUT45), .B(n1247), .ZN(n1253) );
AND2_X1 U949 ( .A1(n1254), .A2(n1037), .ZN(n1028) );
XNOR2_X1 U950 ( .A(n1036), .B(KEYINPUT34), .ZN(n1254) );
XOR2_X1 U951 ( .A(n1176), .B(n1255), .Z(G12) );
XNOR2_X1 U952 ( .A(G110), .B(KEYINPUT0), .ZN(n1255) );
NAND3_X1 U953 ( .A1(n1239), .A2(n1179), .A3(n1032), .ZN(n1176) );
NOR2_X1 U954 ( .A1(n1245), .A2(n1186), .ZN(n1032) );
INV_X1 U955 ( .A(n1222), .ZN(n1186) );
XNOR2_X1 U956 ( .A(n1256), .B(n1061), .ZN(n1222) );
NOR2_X1 U957 ( .A1(n1126), .A2(G902), .ZN(n1061) );
XOR2_X1 U958 ( .A(n1257), .B(n1258), .Z(n1126) );
XNOR2_X1 U959 ( .A(n1088), .B(n1259), .ZN(n1258) );
NOR2_X1 U960 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U961 ( .A(n1262), .B(KEYINPUT16), .Z(n1261) );
NAND2_X1 U962 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U963 ( .A(KEYINPUT52), .B(n1265), .Z(n1263) );
AND2_X1 U964 ( .A1(n1265), .A2(G107), .ZN(n1260) );
INV_X1 U965 ( .A(G134), .ZN(n1088) );
XOR2_X1 U966 ( .A(n1266), .B(n1267), .Z(n1257) );
AND2_X1 U967 ( .A1(n1268), .A2(G217), .ZN(n1267) );
NAND3_X1 U968 ( .A1(n1269), .A2(n1270), .A3(KEYINPUT15), .ZN(n1266) );
NAND2_X1 U969 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U970 ( .A(G128), .B(n1273), .Z(n1271) );
NOR2_X1 U971 ( .A1(G143), .A2(KEYINPUT13), .ZN(n1273) );
OR3_X1 U972 ( .A1(n1162), .A2(G128), .A3(n1272), .ZN(n1269) );
INV_X1 U973 ( .A(KEYINPUT26), .ZN(n1272) );
NAND2_X1 U974 ( .A1(KEYINPUT54), .A2(n1062), .ZN(n1256) );
XOR2_X1 U975 ( .A(G478), .B(KEYINPUT1), .Z(n1062) );
INV_X1 U976 ( .A(n1188), .ZN(n1245) );
XOR2_X1 U977 ( .A(n1058), .B(n1274), .Z(n1188) );
XOR2_X1 U978 ( .A(KEYINPUT29), .B(G475), .Z(n1274) );
NOR2_X1 U979 ( .A1(n1131), .A2(G902), .ZN(n1058) );
XOR2_X1 U980 ( .A(n1275), .B(n1276), .Z(n1131) );
XNOR2_X1 U981 ( .A(n1277), .B(n1278), .ZN(n1276) );
XOR2_X1 U982 ( .A(G122), .B(G113), .Z(n1278) );
XOR2_X1 U983 ( .A(n1279), .B(n1077), .Z(n1275) );
XOR2_X1 U984 ( .A(G131), .B(G143), .Z(n1077) );
XOR2_X1 U985 ( .A(n1280), .B(n1281), .Z(n1279) );
NAND2_X1 U986 ( .A1(n1282), .A2(G214), .ZN(n1280) );
NOR3_X1 U987 ( .A1(n1034), .A2(n1189), .A3(n1250), .ZN(n1179) );
NAND2_X1 U988 ( .A1(n1237), .A2(n1236), .ZN(n1250) );
NAND2_X1 U989 ( .A1(G214), .A2(n1047), .ZN(n1236) );
XNOR2_X1 U990 ( .A(n1283), .B(n1169), .ZN(n1237) );
AND2_X1 U991 ( .A1(G210), .A2(n1047), .ZN(n1169) );
OR2_X1 U992 ( .A1(G902), .A2(G237), .ZN(n1047) );
NAND2_X1 U993 ( .A1(n1284), .A2(n1156), .ZN(n1283) );
XNOR2_X1 U994 ( .A(n1285), .B(n1213), .ZN(n1284) );
XNOR2_X1 U995 ( .A(n1286), .B(n1287), .ZN(n1213) );
XOR2_X1 U996 ( .A(n1113), .B(n1104), .Z(n1287) );
XNOR2_X1 U997 ( .A(n1288), .B(KEYINPUT17), .ZN(n1104) );
INV_X1 U998 ( .A(G110), .ZN(n1288) );
XNOR2_X1 U999 ( .A(n1289), .B(n1290), .ZN(n1113) );
NOR2_X1 U1000 ( .A1(KEYINPUT21), .A2(G113), .ZN(n1290) );
XNOR2_X1 U1001 ( .A(G119), .B(KEYINPUT24), .ZN(n1289) );
XNOR2_X1 U1002 ( .A(n1109), .B(n1265), .ZN(n1286) );
XOR2_X1 U1003 ( .A(G116), .B(G122), .Z(n1265) );
XNOR2_X1 U1004 ( .A(n1291), .B(n1292), .ZN(n1109) );
NAND2_X1 U1005 ( .A1(KEYINPUT44), .A2(n1277), .ZN(n1291) );
INV_X1 U1006 ( .A(G104), .ZN(n1277) );
NAND2_X1 U1007 ( .A1(KEYINPUT3), .A2(n1293), .ZN(n1285) );
XNOR2_X1 U1008 ( .A(n1216), .B(n1089), .ZN(n1293) );
XNOR2_X1 U1009 ( .A(n1148), .B(n1294), .ZN(n1216) );
NOR2_X1 U1010 ( .A1(n1115), .A2(n1295), .ZN(n1294) );
XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n1050), .ZN(n1295) );
INV_X1 U1012 ( .A(G224), .ZN(n1115) );
INV_X1 U1013 ( .A(n1249), .ZN(n1189) );
NAND2_X1 U1014 ( .A1(n1240), .A2(n1296), .ZN(n1249) );
NAND2_X1 U1015 ( .A1(n1242), .A2(n1116), .ZN(n1296) );
INV_X1 U1016 ( .A(G898), .ZN(n1116) );
AND3_X1 U1017 ( .A1(G953), .A2(n1020), .A3(G902), .ZN(n1242) );
NAND3_X1 U1018 ( .A1(n1020), .A2(n1050), .A3(G952), .ZN(n1240) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1297), .ZN(n1020) );
XOR2_X1 U1020 ( .A(KEYINPUT58), .B(G237), .Z(n1297) );
INV_X1 U1021 ( .A(n1234), .ZN(n1034) );
NOR2_X1 U1022 ( .A1(n1037), .A2(n1036), .ZN(n1234) );
AND2_X1 U1023 ( .A1(G221), .A2(n1298), .ZN(n1036) );
XOR2_X1 U1024 ( .A(n1299), .B(G469), .Z(n1037) );
NAND2_X1 U1025 ( .A1(n1300), .A2(n1156), .ZN(n1299) );
XOR2_X1 U1026 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1027 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1028 ( .A(KEYINPUT27), .B(n1162), .ZN(n1304) );
NOR2_X1 U1029 ( .A1(KEYINPUT5), .A2(n1155), .ZN(n1303) );
XNOR2_X1 U1030 ( .A(G104), .B(n1292), .ZN(n1155) );
XNOR2_X1 U1031 ( .A(G101), .B(n1264), .ZN(n1292) );
INV_X1 U1032 ( .A(G107), .ZN(n1264) );
XNOR2_X1 U1033 ( .A(n1152), .B(n1305), .ZN(n1301) );
XOR2_X1 U1034 ( .A(n1306), .B(n1079), .Z(n1305) );
XOR2_X1 U1035 ( .A(n1307), .B(n1147), .Z(n1152) );
NAND2_X1 U1036 ( .A1(G227), .A2(n1050), .ZN(n1307) );
INV_X1 U1037 ( .A(n1042), .ZN(n1239) );
NAND2_X1 U1038 ( .A1(n1308), .A2(n1247), .ZN(n1042) );
XOR2_X1 U1039 ( .A(n1060), .B(G472), .Z(n1247) );
NAND2_X1 U1040 ( .A1(n1309), .A2(n1156), .ZN(n1060) );
XOR2_X1 U1041 ( .A(n1310), .B(n1138), .Z(n1309) );
XOR2_X1 U1042 ( .A(n1311), .B(G101), .Z(n1138) );
NAND2_X1 U1043 ( .A1(n1282), .A2(G210), .ZN(n1311) );
NOR2_X1 U1044 ( .A1(G953), .A2(G237), .ZN(n1282) );
NAND2_X1 U1045 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
OR2_X1 U1046 ( .A1(n1137), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1047 ( .A(n1315), .B(KEYINPUT57), .Z(n1312) );
NAND2_X1 U1048 ( .A1(n1314), .A2(n1137), .ZN(n1315) );
XOR2_X1 U1049 ( .A(G113), .B(n1316), .Z(n1137) );
NOR2_X1 U1050 ( .A1(KEYINPUT32), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1051 ( .A(n1318), .B(n1319), .ZN(n1317) );
NOR2_X1 U1052 ( .A1(G116), .A2(KEYINPUT38), .ZN(n1319) );
XOR2_X1 U1053 ( .A(n1148), .B(n1147), .Z(n1314) );
INV_X1 U1054 ( .A(n1144), .ZN(n1147) );
XNOR2_X1 U1055 ( .A(n1086), .B(n1320), .ZN(n1144) );
NOR2_X1 U1056 ( .A1(G131), .A2(KEYINPUT10), .ZN(n1320) );
XNOR2_X1 U1057 ( .A(G134), .B(G137), .ZN(n1086) );
NAND2_X1 U1058 ( .A1(n1321), .A2(n1322), .ZN(n1148) );
NAND2_X1 U1059 ( .A1(n1323), .A2(n1162), .ZN(n1322) );
INV_X1 U1060 ( .A(G143), .ZN(n1162) );
XOR2_X1 U1061 ( .A(KEYINPUT33), .B(n1324), .Z(n1323) );
NAND2_X1 U1062 ( .A1(n1325), .A2(G143), .ZN(n1321) );
XOR2_X1 U1063 ( .A(KEYINPUT18), .B(n1324), .Z(n1325) );
XOR2_X1 U1064 ( .A(G146), .B(G128), .Z(n1324) );
XOR2_X1 U1065 ( .A(n1052), .B(KEYINPUT47), .Z(n1308) );
XOR2_X1 U1066 ( .A(n1326), .B(n1122), .Z(n1052) );
AND2_X1 U1067 ( .A1(G217), .A2(n1298), .ZN(n1122) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1156), .ZN(n1298) );
NAND2_X1 U1069 ( .A1(n1120), .A2(n1156), .ZN(n1326) );
INV_X1 U1070 ( .A(G902), .ZN(n1156) );
XOR2_X1 U1071 ( .A(n1327), .B(n1328), .Z(n1120) );
XOR2_X1 U1072 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1073 ( .A(n1331), .B(G137), .Z(n1330) );
NAND2_X1 U1074 ( .A1(KEYINPUT4), .A2(n1318), .ZN(n1331) );
INV_X1 U1075 ( .A(G119), .ZN(n1318) );
NAND2_X1 U1076 ( .A1(n1268), .A2(G221), .ZN(n1329) );
AND2_X1 U1077 ( .A1(G234), .A2(n1050), .ZN(n1268) );
INV_X1 U1078 ( .A(G953), .ZN(n1050) );
XNOR2_X1 U1079 ( .A(n1306), .B(n1281), .ZN(n1327) );
XOR2_X1 U1080 ( .A(n1079), .B(n1089), .Z(n1281) );
XOR2_X1 U1081 ( .A(G125), .B(KEYINPUT22), .Z(n1089) );
XOR2_X1 U1082 ( .A(G140), .B(G146), .Z(n1079) );
XOR2_X1 U1083 ( .A(G110), .B(G128), .Z(n1306) );
endmodule


