//Key = 1110011010010101001110111001110101000101111010010011111000000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336;

XOR2_X1 U732 ( .A(n1016), .B(n1017), .Z(G9) );
NOR2_X1 U733 ( .A1(KEYINPUT12), .A2(n1018), .ZN(n1017) );
NAND2_X1 U734 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NAND3_X1 U735 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
INV_X1 U736 ( .A(KEYINPUT13), .ZN(n1023) );
NAND3_X1 U737 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1022) );
NAND3_X1 U738 ( .A1(n1027), .A2(n1026), .A3(KEYINPUT13), .ZN(n1019) );
INV_X1 U739 ( .A(n1028), .ZN(n1026) );
NOR2_X1 U740 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U741 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
NOR2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR3_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
INV_X1 U745 ( .A(n1041), .ZN(n1040) );
NOR3_X1 U746 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1039) );
NOR3_X1 U747 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1042) );
NOR2_X1 U749 ( .A1(n1050), .A2(n1024), .ZN(n1048) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U751 ( .A1(n1047), .A2(n1053), .A3(n1049), .ZN(n1036) );
INV_X1 U752 ( .A(n1054), .ZN(n1049) );
NOR3_X1 U753 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1053) );
NOR2_X1 U754 ( .A1(n1058), .A2(n1038), .ZN(n1057) );
AND2_X1 U755 ( .A1(n1041), .A2(n1059), .ZN(n1056) );
NOR3_X1 U756 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U757 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1031) );
NOR4_X1 U758 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XNOR2_X1 U759 ( .A(n1068), .B(KEYINPUT15), .ZN(n1067) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
INV_X1 U761 ( .A(n1045), .ZN(n1064) );
NOR3_X1 U762 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U764 ( .A(KEYINPUT33), .ZN(n1075) );
NOR2_X1 U765 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
AND3_X1 U766 ( .A1(KEYINPUT19), .A2(n1070), .A3(n1069), .ZN(n1077) );
NOR2_X1 U767 ( .A1(KEYINPUT19), .A2(n1069), .ZN(n1076) );
NOR2_X1 U768 ( .A1(KEYINPUT33), .A2(n1078), .ZN(n1072) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U770 ( .A(KEYINPUT19), .B(n1081), .ZN(n1080) );
XNOR2_X1 U771 ( .A(KEYINPUT49), .B(n1082), .ZN(n1071) );
XNOR2_X1 U772 ( .A(KEYINPUT0), .B(n1083), .ZN(n1061) );
XOR2_X1 U773 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U774 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U776 ( .A1(G953), .A2(n1090), .ZN(n1089) );
XOR2_X1 U777 ( .A(n1091), .B(n1092), .Z(n1088) );
XOR2_X1 U778 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U779 ( .A(G131), .B(n1095), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1096), .A2(KEYINPUT56), .ZN(n1095) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U782 ( .A(n1099), .B(KEYINPUT31), .Z(n1098) );
NAND2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U784 ( .A(n1102), .B(KEYINPUT43), .Z(n1100) );
NOR2_X1 U785 ( .A1(n1102), .A2(n1101), .ZN(n1097) );
INV_X1 U786 ( .A(G134), .ZN(n1101) );
XNOR2_X1 U787 ( .A(G137), .B(KEYINPUT24), .ZN(n1102) );
NAND2_X1 U788 ( .A1(n1103), .A2(n1104), .ZN(n1086) );
XNOR2_X1 U789 ( .A(G953), .B(KEYINPUT36), .ZN(n1103) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1084) );
AND2_X1 U791 ( .A1(G227), .A2(G900), .ZN(n1105) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(G69) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1111), .A2(n1106), .ZN(n1110) );
XOR2_X1 U795 ( .A(KEYINPUT62), .B(n1112), .Z(n1111) );
NAND3_X1 U796 ( .A1(G898), .A2(G224), .A3(G953), .ZN(n1109) );
OR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(G66) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1118) );
AND2_X1 U801 ( .A1(n1121), .A2(KEYINPUT27), .ZN(n1120) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
NOR2_X1 U803 ( .A1(KEYINPUT27), .A2(n1121), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1124), .ZN(G63) );
XNOR2_X1 U805 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U806 ( .A1(n1122), .A2(G478), .ZN(n1125) );
NOR2_X1 U807 ( .A1(n1115), .A2(n1127), .ZN(G60) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U810 ( .A1(n1122), .A2(G475), .ZN(n1131) );
NAND2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1128) );
INV_X1 U813 ( .A(KEYINPUT57), .ZN(n1133) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(G6) );
NAND2_X1 U815 ( .A1(G104), .A2(n1136), .ZN(n1135) );
XOR2_X1 U816 ( .A(KEYINPUT8), .B(n1137), .Z(n1134) );
NOR2_X1 U817 ( .A1(G104), .A2(n1136), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1115), .A2(n1138), .ZN(G57) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U820 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U821 ( .A1(KEYINPUT7), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U822 ( .A(KEYINPUT59), .B(n1144), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
XOR2_X1 U824 ( .A(n1147), .B(KEYINPUT53), .Z(n1146) );
NAND2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1150), .B(KEYINPUT32), .Z(n1148) );
NOR2_X1 U827 ( .A1(n1151), .A2(n1149), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NAND2_X1 U829 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U830 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
XNOR2_X1 U831 ( .A(KEYINPUT60), .B(n1154), .ZN(n1156) );
XOR2_X1 U832 ( .A(n1150), .B(KEYINPUT48), .Z(n1151) );
NAND2_X1 U833 ( .A1(n1122), .A2(G472), .ZN(n1150) );
NOR2_X1 U834 ( .A1(n1115), .A2(n1158), .ZN(G54) );
XOR2_X1 U835 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U836 ( .A1(KEYINPUT35), .A2(n1161), .ZN(n1160) );
XOR2_X1 U837 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U838 ( .A(n1157), .B(n1164), .ZN(n1162) );
NAND2_X1 U839 ( .A1(n1122), .A2(G469), .ZN(n1159) );
NOR2_X1 U840 ( .A1(n1115), .A2(n1165), .ZN(G51) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U843 ( .A1(KEYINPUT10), .A2(n1170), .ZN(n1169) );
NAND2_X1 U844 ( .A1(n1122), .A2(n1079), .ZN(n1168) );
AND2_X1 U845 ( .A1(G902), .A2(n1033), .ZN(n1122) );
NAND2_X1 U846 ( .A1(n1112), .A2(n1171), .ZN(n1033) );
INV_X1 U847 ( .A(n1104), .ZN(n1171) );
NAND4_X1 U848 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1104) );
AND4_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
INV_X1 U850 ( .A(n1180), .ZN(n1178) );
NAND2_X1 U851 ( .A1(n1181), .A2(n1021), .ZN(n1174) );
XOR2_X1 U852 ( .A(n1182), .B(KEYINPUT52), .Z(n1181) );
NAND2_X1 U853 ( .A1(n1054), .A2(n1183), .ZN(n1172) );
NAND2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U857 ( .A1(n1190), .A2(n1191), .A3(KEYINPUT29), .ZN(n1189) );
NAND2_X1 U858 ( .A1(n1192), .A2(n1060), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1193), .A2(n1194), .ZN(n1184) );
INV_X1 U860 ( .A(KEYINPUT29), .ZN(n1194) );
NAND3_X1 U861 ( .A1(n1190), .A2(n1191), .A3(n1186), .ZN(n1193) );
XOR2_X1 U862 ( .A(n1059), .B(KEYINPUT38), .Z(n1190) );
AND4_X1 U863 ( .A1(n1195), .A2(n1136), .A3(n1196), .A4(n1197), .ZN(n1112) );
NOR4_X1 U864 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
INV_X1 U865 ( .A(n1202), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1027), .A2(n1055), .ZN(n1196) );
NAND2_X1 U867 ( .A1(n1028), .A2(n1203), .ZN(n1055) );
NAND2_X1 U868 ( .A1(n1204), .A2(n1060), .ZN(n1203) );
NAND2_X1 U869 ( .A1(n1205), .A2(n1041), .ZN(n1028) );
NAND3_X1 U870 ( .A1(n1059), .A2(n1041), .A3(n1027), .ZN(n1136) );
INV_X1 U871 ( .A(n1206), .ZN(n1027) );
NAND4_X1 U872 ( .A1(n1204), .A2(n1043), .A3(n1205), .A4(n1207), .ZN(n1195) );
XNOR2_X1 U873 ( .A(KEYINPUT1), .B(n1025), .ZN(n1207) );
NOR2_X1 U874 ( .A1(n1106), .A2(G952), .ZN(n1115) );
XNOR2_X1 U875 ( .A(G146), .B(n1173), .ZN(G48) );
NAND2_X1 U876 ( .A1(n1208), .A2(n1059), .ZN(n1173) );
XOR2_X1 U877 ( .A(n1209), .B(n1210), .Z(G45) );
XOR2_X1 U878 ( .A(KEYINPUT45), .B(G143), .Z(n1210) );
NOR2_X1 U879 ( .A1(n1211), .A2(n1182), .ZN(n1209) );
NAND4_X1 U880 ( .A1(n1186), .A2(n1204), .A3(n1212), .A4(n1213), .ZN(n1182) );
XOR2_X1 U881 ( .A(G140), .B(n1214), .Z(G42) );
NOR2_X1 U882 ( .A1(n1058), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U883 ( .A(G137), .B(n1216), .ZN(G39) );
NAND4_X1 U884 ( .A1(n1217), .A2(n1186), .A3(n1060), .A4(n1218), .ZN(n1216) );
XOR2_X1 U885 ( .A(KEYINPUT26), .B(n1192), .Z(n1218) );
XNOR2_X1 U886 ( .A(KEYINPUT41), .B(n1054), .ZN(n1217) );
XNOR2_X1 U887 ( .A(G134), .B(n1179), .ZN(G36) );
NAND4_X1 U888 ( .A1(n1186), .A2(n1204), .A3(n1205), .A4(n1054), .ZN(n1179) );
XNOR2_X1 U889 ( .A(G131), .B(n1219), .ZN(G33) );
NAND2_X1 U890 ( .A1(KEYINPUT6), .A2(n1180), .ZN(n1219) );
NOR2_X1 U891 ( .A1(n1215), .A2(n1220), .ZN(n1180) );
INV_X1 U892 ( .A(n1204), .ZN(n1220) );
NAND3_X1 U893 ( .A1(n1054), .A2(n1059), .A3(n1186), .ZN(n1215) );
NAND2_X1 U894 ( .A1(n1221), .A2(n1222), .ZN(n1054) );
OR2_X1 U895 ( .A1(n1211), .A2(KEYINPUT50), .ZN(n1222) );
NAND3_X1 U896 ( .A1(n1223), .A2(n1045), .A3(KEYINPUT50), .ZN(n1221) );
XOR2_X1 U897 ( .A(n1177), .B(n1224), .Z(G30) );
NOR2_X1 U898 ( .A1(G128), .A2(KEYINPUT21), .ZN(n1224) );
NAND2_X1 U899 ( .A1(n1208), .A2(n1205), .ZN(n1177) );
AND3_X1 U900 ( .A1(n1192), .A2(n1021), .A3(n1186), .ZN(n1208) );
AND2_X1 U901 ( .A1(n1024), .A2(n1225), .ZN(n1186) );
XNOR2_X1 U902 ( .A(G101), .B(n1226), .ZN(G3) );
NAND4_X1 U903 ( .A1(n1227), .A2(n1228), .A3(n1204), .A4(n1229), .ZN(n1226) );
NOR2_X1 U904 ( .A1(KEYINPUT16), .A2(n1038), .ZN(n1229) );
NAND2_X1 U905 ( .A1(KEYINPUT11), .A2(n1206), .ZN(n1228) );
NAND2_X1 U906 ( .A1(n1230), .A2(n1231), .ZN(n1227) );
INV_X1 U907 ( .A(KEYINPUT11), .ZN(n1231) );
NAND3_X1 U908 ( .A1(n1025), .A2(n1211), .A3(n1024), .ZN(n1230) );
XNOR2_X1 U909 ( .A(G125), .B(n1176), .ZN(G27) );
NAND4_X1 U910 ( .A1(n1043), .A2(n1191), .A3(n1059), .A4(n1225), .ZN(n1176) );
NAND2_X1 U911 ( .A1(n1035), .A2(n1232), .ZN(n1225) );
NAND4_X1 U912 ( .A1(G902), .A2(n1233), .A3(n1234), .A4(n1090), .ZN(n1232) );
INV_X1 U913 ( .A(G900), .ZN(n1090) );
XNOR2_X1 U914 ( .A(KEYINPUT14), .B(n1106), .ZN(n1233) );
INV_X1 U915 ( .A(n1058), .ZN(n1191) );
XOR2_X1 U916 ( .A(n1201), .B(n1235), .Z(G24) );
NOR2_X1 U917 ( .A1(KEYINPUT58), .A2(n1236), .ZN(n1235) );
AND4_X1 U918 ( .A1(n1237), .A2(n1041), .A3(n1212), .A4(n1213), .ZN(n1201) );
NAND2_X1 U919 ( .A1(n1238), .A2(n1239), .ZN(n1041) );
OR2_X1 U920 ( .A1(n1058), .A2(KEYINPUT2), .ZN(n1239) );
NAND3_X1 U921 ( .A1(n1082), .A2(n1240), .A3(KEYINPUT2), .ZN(n1238) );
XOR2_X1 U922 ( .A(G119), .B(n1200), .Z(G21) );
AND3_X1 U923 ( .A1(n1237), .A2(n1060), .A3(n1192), .ZN(n1200) );
NOR2_X1 U924 ( .A1(n1240), .A2(n1082), .ZN(n1192) );
INV_X1 U925 ( .A(n1068), .ZN(n1240) );
XNOR2_X1 U926 ( .A(G116), .B(n1241), .ZN(G18) );
NAND4_X1 U927 ( .A1(n1242), .A2(n1204), .A3(n1043), .A4(n1205), .ZN(n1241) );
NOR2_X1 U928 ( .A1(n1213), .A2(n1243), .ZN(n1205) );
XOR2_X1 U929 ( .A(n1025), .B(KEYINPUT17), .Z(n1242) );
XNOR2_X1 U930 ( .A(G113), .B(n1202), .ZN(G15) );
NAND3_X1 U931 ( .A1(n1237), .A2(n1059), .A3(n1204), .ZN(n1202) );
NOR2_X1 U932 ( .A1(n1068), .A2(n1082), .ZN(n1204) );
NAND2_X1 U933 ( .A1(n1244), .A2(n1245), .ZN(n1059) );
OR2_X1 U934 ( .A1(n1038), .A2(KEYINPUT39), .ZN(n1245) );
NAND3_X1 U935 ( .A1(n1213), .A2(n1243), .A3(KEYINPUT39), .ZN(n1244) );
INV_X1 U936 ( .A(n1212), .ZN(n1243) );
AND2_X1 U937 ( .A1(n1043), .A2(n1025), .ZN(n1237) );
NOR2_X1 U938 ( .A1(n1047), .A2(n1211), .ZN(n1043) );
NAND2_X1 U939 ( .A1(n1083), .A2(n1052), .ZN(n1047) );
XOR2_X1 U940 ( .A(G110), .B(n1198), .Z(G12) );
NOR3_X1 U941 ( .A1(n1206), .A2(n1058), .A3(n1038), .ZN(n1198) );
INV_X1 U942 ( .A(n1060), .ZN(n1038) );
NOR2_X1 U943 ( .A1(n1212), .A2(n1213), .ZN(n1060) );
XNOR2_X1 U944 ( .A(n1246), .B(n1247), .ZN(n1213) );
XOR2_X1 U945 ( .A(KEYINPUT3), .B(G475), .Z(n1247) );
NAND2_X1 U946 ( .A1(n1132), .A2(n1248), .ZN(n1246) );
XOR2_X1 U947 ( .A(n1249), .B(n1250), .Z(n1132) );
XOR2_X1 U948 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U949 ( .A(n1236), .B(G113), .ZN(n1252) );
INV_X1 U950 ( .A(G122), .ZN(n1236) );
XNOR2_X1 U951 ( .A(KEYINPUT51), .B(n1253), .ZN(n1251) );
XOR2_X1 U952 ( .A(n1254), .B(n1255), .Z(n1249) );
XOR2_X1 U953 ( .A(n1093), .B(n1256), .Z(n1255) );
XNOR2_X1 U954 ( .A(G104), .B(n1257), .ZN(n1254) );
AND3_X1 U955 ( .A1(G214), .A2(n1106), .A3(n1258), .ZN(n1257) );
XOR2_X1 U956 ( .A(G478), .B(n1259), .Z(n1212) );
NOR2_X1 U957 ( .A1(n1260), .A2(n1126), .ZN(n1259) );
XNOR2_X1 U958 ( .A(n1261), .B(n1262), .ZN(n1126) );
XOR2_X1 U959 ( .A(n1263), .B(n1264), .Z(n1262) );
AND3_X1 U960 ( .A1(G217), .A2(n1106), .A3(G234), .ZN(n1263) );
XOR2_X1 U961 ( .A(n1265), .B(n1266), .Z(n1261) );
NOR2_X1 U962 ( .A1(KEYINPUT63), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U963 ( .A(n1268), .B(n1018), .ZN(n1267) );
NAND2_X1 U964 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U965 ( .A1(G122), .A2(n1271), .ZN(n1270) );
XOR2_X1 U966 ( .A(KEYINPUT37), .B(n1272), .Z(n1269) );
NOR2_X1 U967 ( .A1(G122), .A2(n1271), .ZN(n1272) );
INV_X1 U968 ( .A(G116), .ZN(n1271) );
XNOR2_X1 U969 ( .A(G134), .B(KEYINPUT4), .ZN(n1265) );
XNOR2_X1 U970 ( .A(G902), .B(KEYINPUT23), .ZN(n1260) );
NAND2_X1 U971 ( .A1(n1082), .A2(n1068), .ZN(n1058) );
XNOR2_X1 U972 ( .A(n1273), .B(n1123), .ZN(n1068) );
AND2_X1 U973 ( .A1(G217), .A2(n1274), .ZN(n1123) );
OR2_X1 U974 ( .A1(n1121), .A2(G902), .ZN(n1273) );
XNOR2_X1 U975 ( .A(n1275), .B(n1276), .ZN(n1121) );
XOR2_X1 U976 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U977 ( .A(G137), .B(G146), .ZN(n1278) );
NAND3_X1 U978 ( .A1(G234), .A2(n1106), .A3(G221), .ZN(n1277) );
XOR2_X1 U979 ( .A(n1279), .B(n1280), .Z(n1275) );
XNOR2_X1 U980 ( .A(n1281), .B(n1282), .ZN(n1279) );
NAND2_X1 U981 ( .A1(KEYINPUT40), .A2(n1283), .ZN(n1282) );
NAND2_X1 U982 ( .A1(KEYINPUT44), .A2(n1093), .ZN(n1281) );
XOR2_X1 U983 ( .A(G125), .B(G140), .Z(n1093) );
XOR2_X1 U984 ( .A(n1284), .B(G472), .Z(n1082) );
NAND2_X1 U985 ( .A1(n1248), .A2(n1285), .ZN(n1284) );
NAND2_X1 U986 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U987 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U988 ( .A(n1157), .B(n1154), .ZN(n1289) );
XNOR2_X1 U989 ( .A(n1290), .B(n1144), .ZN(n1288) );
INV_X1 U990 ( .A(G101), .ZN(n1144) );
XOR2_X1 U991 ( .A(n1291), .B(KEYINPUT55), .Z(n1286) );
NAND2_X1 U992 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U993 ( .A(G101), .B(n1290), .ZN(n1293) );
NAND2_X1 U994 ( .A1(KEYINPUT28), .A2(n1141), .ZN(n1290) );
AND3_X1 U995 ( .A1(n1258), .A2(n1106), .A3(G210), .ZN(n1141) );
XNOR2_X1 U996 ( .A(n1154), .B(n1155), .ZN(n1292) );
XOR2_X1 U997 ( .A(n1294), .B(n1295), .Z(n1154) );
XNOR2_X1 U998 ( .A(n1296), .B(n1297), .ZN(n1295) );
XNOR2_X1 U999 ( .A(G119), .B(G113), .ZN(n1294) );
NAND3_X1 U1000 ( .A1(n1024), .A2(n1025), .A3(n1021), .ZN(n1206) );
INV_X1 U1001 ( .A(n1211), .ZN(n1021) );
NAND2_X1 U1002 ( .A1(n1046), .A2(n1045), .ZN(n1211) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1298), .ZN(n1045) );
INV_X1 U1004 ( .A(n1223), .ZN(n1046) );
XOR2_X1 U1005 ( .A(n1069), .B(n1299), .Z(n1223) );
NOR2_X1 U1006 ( .A1(n1079), .A2(KEYINPUT9), .ZN(n1299) );
INV_X1 U1007 ( .A(n1070), .ZN(n1079) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1298), .ZN(n1070) );
NAND2_X1 U1009 ( .A1(n1258), .A2(n1248), .ZN(n1298) );
INV_X1 U1010 ( .A(G237), .ZN(n1258) );
INV_X1 U1011 ( .A(n1081), .ZN(n1069) );
NAND2_X1 U1012 ( .A1(n1300), .A2(n1248), .ZN(n1081) );
XNOR2_X1 U1013 ( .A(n1166), .B(n1170), .ZN(n1300) );
INV_X1 U1014 ( .A(n1113), .ZN(n1170) );
XNOR2_X1 U1015 ( .A(n1301), .B(n1302), .ZN(n1113) );
XOR2_X1 U1016 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1017 ( .A(G122), .B(G101), .ZN(n1304) );
NAND2_X1 U1018 ( .A1(KEYINPUT20), .A2(n1305), .ZN(n1303) );
INV_X1 U1019 ( .A(G113), .ZN(n1305) );
XOR2_X1 U1020 ( .A(n1306), .B(n1307), .Z(n1301) );
XOR2_X1 U1021 ( .A(n1308), .B(n1280), .Z(n1306) );
XOR2_X1 U1022 ( .A(G110), .B(G119), .Z(n1280) );
NAND2_X1 U1023 ( .A1(KEYINPUT61), .A2(n1297), .ZN(n1308) );
XOR2_X1 U1024 ( .A(G116), .B(KEYINPUT47), .Z(n1297) );
XOR2_X1 U1025 ( .A(n1309), .B(n1310), .Z(n1166) );
XOR2_X1 U1026 ( .A(KEYINPUT30), .B(G125), .Z(n1310) );
XOR2_X1 U1027 ( .A(n1296), .B(n1311), .Z(n1309) );
AND2_X1 U1028 ( .A1(n1106), .A2(G224), .ZN(n1311) );
NAND3_X1 U1029 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1296) );
NAND2_X1 U1030 ( .A1(G128), .A2(n1315), .ZN(n1314) );
OR3_X1 U1031 ( .A1(n1315), .A2(G128), .A3(KEYINPUT25), .ZN(n1313) );
NAND2_X1 U1032 ( .A1(KEYINPUT5), .A2(n1256), .ZN(n1315) );
INV_X1 U1033 ( .A(n1316), .ZN(n1256) );
NAND2_X1 U1034 ( .A1(KEYINPUT25), .A2(n1316), .ZN(n1312) );
XNOR2_X1 U1035 ( .A(G143), .B(G146), .ZN(n1316) );
NAND2_X1 U1036 ( .A1(n1035), .A2(n1317), .ZN(n1025) );
NAND3_X1 U1037 ( .A1(n1114), .A2(n1234), .A3(G902), .ZN(n1317) );
NOR2_X1 U1038 ( .A1(n1106), .A2(G898), .ZN(n1114) );
NAND3_X1 U1039 ( .A1(n1234), .A2(n1106), .A3(G952), .ZN(n1035) );
NAND2_X1 U1040 ( .A1(G237), .A2(G234), .ZN(n1234) );
NOR2_X1 U1041 ( .A1(n1083), .A2(n1065), .ZN(n1024) );
INV_X1 U1042 ( .A(n1052), .ZN(n1065) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1274), .ZN(n1052) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1248), .ZN(n1274) );
INV_X1 U1045 ( .A(n1051), .ZN(n1083) );
XNOR2_X1 U1046 ( .A(n1318), .B(G469), .ZN(n1051) );
NAND2_X1 U1047 ( .A1(n1319), .A2(n1248), .ZN(n1318) );
INV_X1 U1048 ( .A(G902), .ZN(n1248) );
XOR2_X1 U1049 ( .A(n1164), .B(n1320), .Z(n1319) );
XOR2_X1 U1050 ( .A(KEYINPUT34), .B(n1321), .Z(n1320) );
NOR2_X1 U1051 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1052 ( .A(n1324), .B(KEYINPUT42), .Z(n1323) );
NAND2_X1 U1053 ( .A1(n1325), .A2(n1155), .ZN(n1324) );
XOR2_X1 U1054 ( .A(KEYINPUT22), .B(n1326), .Z(n1325) );
AND2_X1 U1055 ( .A1(n1326), .A2(n1157), .ZN(n1322) );
INV_X1 U1056 ( .A(n1155), .ZN(n1157) );
NAND2_X1 U1057 ( .A1(n1327), .A2(n1328), .ZN(n1155) );
NAND2_X1 U1058 ( .A1(n1329), .A2(n1253), .ZN(n1328) );
XOR2_X1 U1059 ( .A(KEYINPUT18), .B(n1330), .Z(n1327) );
NOR2_X1 U1060 ( .A1(n1329), .A2(n1253), .ZN(n1330) );
INV_X1 U1061 ( .A(G131), .ZN(n1253) );
XNOR2_X1 U1062 ( .A(G137), .B(G134), .ZN(n1329) );
XOR2_X1 U1063 ( .A(n1163), .B(KEYINPUT46), .Z(n1326) );
XNOR2_X1 U1064 ( .A(n1331), .B(n1094), .ZN(n1163) );
XOR2_X1 U1065 ( .A(G146), .B(n1264), .Z(n1094) );
XNOR2_X1 U1066 ( .A(G143), .B(n1283), .ZN(n1264) );
INV_X1 U1067 ( .A(G128), .ZN(n1283) );
NAND2_X1 U1068 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1069 ( .A1(G101), .A2(n1307), .ZN(n1333) );
XOR2_X1 U1070 ( .A(KEYINPUT54), .B(n1334), .Z(n1332) );
NOR2_X1 U1071 ( .A1(G101), .A2(n1307), .ZN(n1334) );
XNOR2_X1 U1072 ( .A(n1018), .B(G104), .ZN(n1307) );
INV_X1 U1073 ( .A(G107), .ZN(n1018) );
XNOR2_X1 U1074 ( .A(n1335), .B(n1336), .ZN(n1164) );
XOR2_X1 U1075 ( .A(G140), .B(G110), .Z(n1336) );
NAND2_X1 U1076 ( .A1(G227), .A2(n1106), .ZN(n1335) );
INV_X1 U1077 ( .A(G953), .ZN(n1106) );
endmodule


