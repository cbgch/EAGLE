//Key = 1100111000011100111011011010110101100100010001100110111010101001


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
n2182, n2183, n2184, n2185, n2186, n2187, n2188;

XOR2_X2 U1228 ( .A(n2174), .B(KEYINPUT22), .Z(n1917) );
INV_X2 U1229 ( .A(n1790), .ZN(n1776) );
INV_X2 U1230 ( .A(U280), .ZN(n1775) );
NAND2_X1 U1231 ( .A1(n1642), .A2(n1643), .ZN(U344) );
NAND2_X1 U1232 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1644), .ZN(n1643) );
NAND2_X1 U1233 ( .A1(n1645), .A2(DATA_IN_7_), .ZN(n1642) );
NAND2_X1 U1234 ( .A1(n1646), .A2(n1647), .ZN(U343) );
NAND2_X1 U1235 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1644), .ZN(n1647) );
NAND2_X1 U1236 ( .A1(n1645), .A2(DATA_IN_6_), .ZN(n1646) );
NAND2_X1 U1237 ( .A1(n1648), .A2(n1649), .ZN(U342) );
NAND2_X1 U1238 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1644), .ZN(n1649) );
NAND2_X1 U1239 ( .A1(n1645), .A2(DATA_IN_5_), .ZN(n1648) );
NAND2_X1 U1240 ( .A1(n1650), .A2(n1651), .ZN(U341) );
NAND2_X1 U1241 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1644), .ZN(n1651) );
NAND2_X1 U1242 ( .A1(n1645), .A2(DATA_IN_4_), .ZN(n1650) );
NAND2_X1 U1243 ( .A1(n1652), .A2(n1653), .ZN(U340) );
NAND2_X1 U1244 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1644), .ZN(n1653) );
NAND2_X1 U1245 ( .A1(n1645), .A2(DATA_IN_3_), .ZN(n1652) );
NAND2_X1 U1246 ( .A1(n1654), .A2(n1655), .ZN(U339) );
NAND2_X1 U1247 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1644), .ZN(n1655) );
NAND2_X1 U1248 ( .A1(n1645), .A2(DATA_IN_2_), .ZN(n1654) );
NAND2_X1 U1249 ( .A1(n1656), .A2(n1657), .ZN(U338) );
NAND2_X1 U1250 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1644), .ZN(n1657) );
NAND2_X1 U1251 ( .A1(n1645), .A2(DATA_IN_1_), .ZN(n1656) );
NAND2_X1 U1252 ( .A1(n1658), .A2(n1659), .ZN(U337) );
NAND2_X1 U1253 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1644), .ZN(n1659) );
NAND2_X1 U1254 ( .A1(n1645), .A2(DATA_IN_0_), .ZN(n1658) );
INV_X1 U1255 ( .A(n1644), .ZN(n1645) );
NAND2_X1 U1256 ( .A1(n1660), .A2(n1661), .ZN(n1644) );
NAND3_X1 U1257 ( .A1(n1662), .A2(n1663), .A3(n1664), .ZN(n1661) );
NAND2_X1 U1258 ( .A1(n1665), .A2(n1666), .ZN(U336) );
NAND2_X1 U1259 ( .A1(n1667), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1666) );
NAND2_X1 U1260 ( .A1(n1668), .A2(DATA_IN_7_), .ZN(n1665) );
NAND2_X1 U1261 ( .A1(n1669), .A2(n1670), .ZN(U335) );
NAND2_X1 U1262 ( .A1(n1667), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1670) );
NAND2_X1 U1263 ( .A1(n1668), .A2(DATA_IN_6_), .ZN(n1669) );
NAND2_X1 U1264 ( .A1(n1671), .A2(n1672), .ZN(U334) );
NAND2_X1 U1265 ( .A1(n1667), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1672) );
NAND2_X1 U1266 ( .A1(n1668), .A2(DATA_IN_5_), .ZN(n1671) );
NAND2_X1 U1267 ( .A1(n1673), .A2(n1674), .ZN(U333) );
NAND2_X1 U1268 ( .A1(n1667), .A2(RMIN_REG_4__SCAN_IN), .ZN(n1674) );
NAND2_X1 U1269 ( .A1(n1668), .A2(DATA_IN_4_), .ZN(n1673) );
NAND2_X1 U1270 ( .A1(n1675), .A2(n1676), .ZN(U332) );
NAND2_X1 U1271 ( .A1(n1667), .A2(RMIN_REG_3__SCAN_IN), .ZN(n1676) );
NAND2_X1 U1272 ( .A1(n1668), .A2(DATA_IN_3_), .ZN(n1675) );
NAND2_X1 U1273 ( .A1(n1677), .A2(n1678), .ZN(U331) );
NAND2_X1 U1274 ( .A1(n1667), .A2(RMIN_REG_2__SCAN_IN), .ZN(n1678) );
NAND2_X1 U1275 ( .A1(n1668), .A2(DATA_IN_2_), .ZN(n1677) );
NAND2_X1 U1276 ( .A1(n1679), .A2(n1680), .ZN(U330) );
NAND2_X1 U1277 ( .A1(n1667), .A2(RMIN_REG_1__SCAN_IN), .ZN(n1680) );
NAND2_X1 U1278 ( .A1(n1668), .A2(DATA_IN_1_), .ZN(n1679) );
NAND2_X1 U1279 ( .A1(n1681), .A2(n1682), .ZN(U329) );
NAND2_X1 U1280 ( .A1(n1667), .A2(RMIN_REG_0__SCAN_IN), .ZN(n1682) );
AND2_X1 U1281 ( .A1(n1683), .A2(n1684), .ZN(n1667) );
OR3_X1 U1282 ( .A1(n1685), .A2(U375), .A3(KEYINPUT12), .ZN(n1684) );
INV_X1 U1283 ( .A(n1660), .ZN(U375) );
NAND2_X1 U1284 ( .A1(KEYINPUT12), .A2(n1668), .ZN(n1683) );
NAND2_X1 U1285 ( .A1(n1668), .A2(DATA_IN_0_), .ZN(n1681) );
AND2_X1 U1286 ( .A1(n1685), .A2(n1660), .ZN(n1668) );
NAND2_X1 U1287 ( .A1(n1663), .A2(n1686), .ZN(n1685) );
NAND2_X1 U1288 ( .A1(n1687), .A2(n1662), .ZN(n1686) );
NAND3_X1 U1289 ( .A1(n1688), .A2(n1689), .A3(n1690), .ZN(n1662) );
NAND2_X1 U1290 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1691), .ZN(n1690) );
NAND3_X1 U1291 ( .A1(n1692), .A2(n1693), .A3(n1694), .ZN(n1689) );
OR2_X1 U1292 ( .A1(n1691), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1694) );
NAND3_X1 U1293 ( .A1(n1695), .A2(n1696), .A3(n1697), .ZN(n1693) );
NAND2_X1 U1294 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1698), .ZN(n1697) );
NAND3_X1 U1295 ( .A1(n1699), .A2(n1700), .A3(n1701), .ZN(n1696) );
NAND2_X1 U1296 ( .A1(DATA_IN_4_), .A2(n1702), .ZN(n1701) );
NAND3_X1 U1297 ( .A1(n1703), .A2(n1704), .A3(n1705), .ZN(n1700) );
NAND2_X1 U1298 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1706), .ZN(n1705) );
XOR2_X1 U1299 ( .A(KEYINPUT53), .B(DATA_IN_2_), .Z(n1706) );
NAND3_X1 U1300 ( .A1(n1707), .A2(n1708), .A3(n1709), .ZN(n1704) );
OR2_X1 U1301 ( .A1(n1710), .A2(RMAX_REG_2__SCAN_IN), .ZN(n1709) );
NAND3_X1 U1302 ( .A1(n1711), .A2(n1712), .A3(DATA_IN_0_), .ZN(n1708) );
NAND2_X1 U1303 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1713), .ZN(n1711) );
NAND2_X1 U1304 ( .A1(DATA_IN_1_), .A2(n1714), .ZN(n1707) );
NAND2_X1 U1305 ( .A1(n1715), .A2(n1716), .ZN(n1703) );
XOR2_X1 U1306 ( .A(n1717), .B(KEYINPUT0), .Z(n1715) );
NAND2_X1 U1307 ( .A1(DATA_IN_3_), .A2(n1718), .ZN(n1699) );
XOR2_X1 U1308 ( .A(RMAX_REG_3__SCAN_IN), .B(KEYINPUT13), .Z(n1718) );
NAND2_X1 U1309 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1719), .ZN(n1695) );
OR2_X1 U1310 ( .A1(n1698), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1692) );
NAND2_X1 U1311 ( .A1(DATA_IN_7_), .A2(n1720), .ZN(n1688) );
XOR2_X1 U1312 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT11), .Z(n1720) );
NAND2_X1 U1313 ( .A1(n1721), .A2(n1722), .ZN(n1687) );
OR2_X1 U1314 ( .A1(n1723), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1722) );
NAND4_X1 U1315 ( .A1(n1724), .A2(n1725), .A3(n1726), .A4(n1664), .ZN(n1721));
NAND2_X1 U1316 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1723), .ZN(n1664) );
NAND3_X1 U1317 ( .A1(n1727), .A2(n1728), .A3(n1729), .ZN(n1726) );
NAND2_X1 U1318 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1698), .ZN(n1729) );
NAND3_X1 U1319 ( .A1(n1730), .A2(n1731), .A3(n1732), .ZN(n1728) );
OR2_X1 U1320 ( .A1(n1698), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1732) );
NAND3_X1 U1321 ( .A1(n1733), .A2(n1734), .A3(n1735), .ZN(n1731) );
NAND2_X1 U1322 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1719), .ZN(n1735) );
INV_X1 U1323 ( .A(DATA_IN_4_), .ZN(n1719) );
NAND3_X1 U1324 ( .A1(n1736), .A2(n1737), .A3(n1738), .ZN(n1734) );
NAND2_X1 U1325 ( .A1(DATA_IN_3_), .A2(n1739), .ZN(n1738) );
NAND3_X1 U1326 ( .A1(n1740), .A2(n1741), .A3(n1742), .ZN(n1737) );
NAND2_X1 U1327 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1710), .ZN(n1742) );
NAND3_X1 U1328 ( .A1(n1743), .A2(n1744), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1741) );
NAND2_X1 U1329 ( .A1(DATA_IN_1_), .A2(n1745), .ZN(n1743) );
NAND2_X1 U1330 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1713), .ZN(n1740) );
INV_X1 U1331 ( .A(DATA_IN_1_), .ZN(n1713) );
NAND2_X1 U1332 ( .A1(n1746), .A2(DATA_IN_2_), .ZN(n1736) );
XNOR2_X1 U1333 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT42), .ZN(n1746) );
NAND2_X1 U1334 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1716), .ZN(n1733) );
NAND2_X1 U1335 ( .A1(n1747), .A2(DATA_IN_4_), .ZN(n1730) );
XOR2_X1 U1336 ( .A(n1748), .B(KEYINPUT3), .Z(n1747) );
NAND2_X1 U1337 ( .A1(n1749), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1727) );
XOR2_X1 U1338 ( .A(n1691), .B(KEYINPUT39), .Z(n1749) );
OR2_X1 U1339 ( .A1(n1691), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1725) );
INV_X1 U1340 ( .A(DATA_IN_6_), .ZN(n1691) );
NAND2_X1 U1341 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1723), .ZN(n1724) );
NAND2_X1 U1342 ( .A1(n1750), .A2(n1751), .ZN(U328) );
NAND2_X1 U1343 ( .A1(n1752), .A2(DATA_IN_7_), .ZN(n1751) );
XOR2_X1 U1344 ( .A(n1753), .B(KEYINPUT43), .Z(n1750) );
NAND2_X1 U1345 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1754), .ZN(n1753) );
NAND2_X1 U1346 ( .A1(n1755), .A2(n1756), .ZN(U327) );
NAND2_X1 U1347 ( .A1(n1752), .A2(DATA_IN_6_), .ZN(n1756) );
NAND2_X1 U1348 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1754), .ZN(n1755) );
NAND2_X1 U1349 ( .A1(n1757), .A2(n1758), .ZN(U326) );
NAND2_X1 U1350 ( .A1(n1752), .A2(DATA_IN_5_), .ZN(n1758) );
NAND2_X1 U1351 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1754), .ZN(n1757) );
NAND2_X1 U1352 ( .A1(n1759), .A2(n1760), .ZN(U325) );
NAND2_X1 U1353 ( .A1(n1752), .A2(DATA_IN_4_), .ZN(n1760) );
NAND2_X1 U1354 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1754), .ZN(n1759) );
NAND2_X1 U1355 ( .A1(n1761), .A2(n1762), .ZN(U324) );
NAND2_X1 U1356 ( .A1(n1752), .A2(DATA_IN_3_), .ZN(n1762) );
NAND2_X1 U1357 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1754), .ZN(n1761) );
NAND2_X1 U1358 ( .A1(n1763), .A2(n1764), .ZN(U323) );
NAND2_X1 U1359 ( .A1(n1752), .A2(DATA_IN_2_), .ZN(n1764) );
NAND2_X1 U1360 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1754), .ZN(n1763) );
NAND2_X1 U1361 ( .A1(n1765), .A2(n1766), .ZN(U322) );
NAND2_X1 U1362 ( .A1(n1752), .A2(DATA_IN_1_), .ZN(n1766) );
NAND2_X1 U1363 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1754), .ZN(n1765) );
NAND2_X1 U1364 ( .A1(n1767), .A2(n1768), .ZN(U321) );
NAND2_X1 U1365 ( .A1(n1752), .A2(DATA_IN_0_), .ZN(n1768) );
AND2_X1 U1366 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1769), .ZN(n1752) );
NAND2_X1 U1367 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1754), .ZN(n1767) );
NAND2_X1 U1368 ( .A1(n1660), .A2(n1769), .ZN(n1754) );
NAND2_X1 U1369 ( .A1(n1663), .A2(n1770), .ZN(n1769) );
NAND2_X1 U1370 ( .A1(n1771), .A2(n1663), .ZN(n1660) );
NAND2_X1 U1371 ( .A1(n1772), .A2(n1773), .ZN(U320) );
NAND2_X1 U1372 ( .A1(n1774), .A2(n1775), .ZN(n1773) );
XNOR2_X1 U1373 ( .A(REG1_REG_7__SCAN_IN), .B(KEYINPUT49), .ZN(n1774) );
NAND2_X1 U1374 ( .A1(n1776), .A2(DATA_IN_7_), .ZN(n1772) );
NAND2_X1 U1375 ( .A1(n1777), .A2(n1778), .ZN(U319) );
NAND2_X1 U1376 ( .A1(n1779), .A2(n1775), .ZN(n1778) );
XOR2_X1 U1377 ( .A(REG1_REG_6__SCAN_IN), .B(KEYINPUT10), .Z(n1779) );
NAND2_X1 U1378 ( .A1(n1776), .A2(DATA_IN_6_), .ZN(n1777) );
NAND2_X1 U1379 ( .A1(n1780), .A2(n1781), .ZN(U318) );
NAND2_X1 U1380 ( .A1(n1776), .A2(DATA_IN_5_), .ZN(n1781) );
NAND2_X1 U1381 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1775), .ZN(n1780) );
NAND2_X1 U1382 ( .A1(n1782), .A2(n1783), .ZN(U317) );
NAND2_X1 U1383 ( .A1(n1776), .A2(DATA_IN_4_), .ZN(n1783) );
NAND2_X1 U1384 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1775), .ZN(n1782) );
NAND2_X1 U1385 ( .A1(n1784), .A2(n1785), .ZN(U316) );
NAND2_X1 U1386 ( .A1(n1776), .A2(DATA_IN_3_), .ZN(n1785) );
XOR2_X1 U1387 ( .A(KEYINPUT52), .B(n1786), .Z(n1784) );
AND2_X1 U1388 ( .A1(n1775), .A2(REG1_REG_3__SCAN_IN), .ZN(n1786) );
NAND2_X1 U1389 ( .A1(n1787), .A2(n1788), .ZN(U315) );
NAND2_X1 U1390 ( .A1(n1789), .A2(DATA_IN_2_), .ZN(n1788) );
XOR2_X1 U1391 ( .A(n1790), .B(KEYINPUT41), .Z(n1789) );
NAND2_X1 U1392 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1775), .ZN(n1787) );
NAND2_X1 U1393 ( .A1(n1791), .A2(n1792), .ZN(U314) );
NAND2_X1 U1394 ( .A1(n1776), .A2(DATA_IN_1_), .ZN(n1792) );
NAND2_X1 U1395 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1775), .ZN(n1791) );
NAND2_X1 U1396 ( .A1(n1793), .A2(n1794), .ZN(U313) );
NAND2_X1 U1397 ( .A1(n1776), .A2(DATA_IN_0_), .ZN(n1794) );
NAND2_X1 U1398 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1775), .ZN(n1793) );
NAND2_X1 U1399 ( .A1(n1795), .A2(n1796), .ZN(U312) );
NAND2_X1 U1400 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1797), .ZN(n1796) );
XOR2_X1 U1401 ( .A(KEYINPUT2), .B(n1776), .Z(n1797) );
NAND2_X1 U1402 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1775), .ZN(n1795) );
NAND2_X1 U1403 ( .A1(n1798), .A2(n1799), .ZN(U311) );
NAND2_X1 U1404 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1776), .ZN(n1799) );
NAND2_X1 U1405 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1775), .ZN(n1798) );
NAND2_X1 U1406 ( .A1(n1800), .A2(n1801), .ZN(U310) );
NAND2_X1 U1407 ( .A1(n1802), .A2(n1776), .ZN(n1801) );
XNOR2_X1 U1408 ( .A(REG1_REG_5__SCAN_IN), .B(KEYINPUT16), .ZN(n1802) );
XOR2_X1 U1409 ( .A(n1803), .B(KEYINPUT27), .Z(n1800) );
NAND2_X1 U1410 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1775), .ZN(n1803) );
NAND2_X1 U1411 ( .A1(n1804), .A2(n1805), .ZN(U309) );
NAND2_X1 U1412 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1776), .ZN(n1805) );
NAND2_X1 U1413 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1775), .ZN(n1804) );
NAND2_X1 U1414 ( .A1(n1806), .A2(n1807), .ZN(U308) );
NAND2_X1 U1415 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1776), .ZN(n1807) );
XOR2_X1 U1416 ( .A(KEYINPUT45), .B(n1808), .Z(n1806) );
AND2_X1 U1417 ( .A1(n1775), .A2(REG2_REG_3__SCAN_IN), .ZN(n1808) );
NAND2_X1 U1418 ( .A1(n1809), .A2(n1810), .ZN(U307) );
NAND2_X1 U1419 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1776), .ZN(n1810) );
NAND2_X1 U1420 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1775), .ZN(n1809) );
NAND2_X1 U1421 ( .A1(n1811), .A2(n1812), .ZN(U306) );
NAND2_X1 U1422 ( .A1(n1813), .A2(REG1_REG_1__SCAN_IN), .ZN(n1812) );
XOR2_X1 U1423 ( .A(n1790), .B(KEYINPUT60), .Z(n1813) );
NAND2_X1 U1424 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1775), .ZN(n1811) );
NAND2_X1 U1425 ( .A1(n1814), .A2(n1815), .ZN(U305) );
NAND2_X1 U1426 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1776), .ZN(n1815) );
NAND2_X1 U1427 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1775), .ZN(n1814) );
NAND2_X1 U1428 ( .A1(n1816), .A2(n1817), .ZN(U304) );
NAND2_X1 U1429 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1776), .ZN(n1817) );
NAND2_X1 U1430 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1775), .ZN(n1816) );
NAND2_X1 U1431 ( .A1(n1818), .A2(n1819), .ZN(U303) );
NAND2_X1 U1432 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1776), .ZN(n1819) );
NAND2_X1 U1433 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1775), .ZN(n1818) );
NAND2_X1 U1434 ( .A1(n1820), .A2(n1821), .ZN(U302) );
NAND2_X1 U1435 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1776), .ZN(n1821) );
NAND2_X1 U1436 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1775), .ZN(n1820) );
NAND2_X1 U1437 ( .A1(n1822), .A2(n1823), .ZN(U301) );
NAND2_X1 U1438 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1776), .ZN(n1823) );
NAND2_X1 U1439 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1775), .ZN(n1822) );
NAND2_X1 U1440 ( .A1(n1824), .A2(n1825), .ZN(U300) );
NAND2_X1 U1441 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1776), .ZN(n1825) );
XOR2_X1 U1442 ( .A(n1826), .B(KEYINPUT48), .Z(n1824) );
NAND2_X1 U1443 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1775), .ZN(n1826) );
NAND2_X1 U1444 ( .A1(n1827), .A2(n1828), .ZN(U299) );
NAND2_X1 U1445 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1829), .ZN(n1828) );
XOR2_X1 U1446 ( .A(KEYINPUT19), .B(n1775), .Z(n1829) );
NAND2_X1 U1447 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1776), .ZN(n1827) );
NAND2_X1 U1448 ( .A1(n1830), .A2(n1831), .ZN(U298) );
NAND2_X1 U1449 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1776), .ZN(n1831) );
NAND2_X1 U1450 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1775), .ZN(n1830) );
NAND2_X1 U1451 ( .A1(n1832), .A2(n1833), .ZN(U297) );
NAND2_X1 U1452 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1776), .ZN(n1833) );
NAND2_X1 U1453 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1775), .ZN(n1832) );
NAND2_X1 U1454 ( .A1(n1834), .A2(n1835), .ZN(U296) );
NAND2_X1 U1455 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1776), .ZN(n1835) );
NAND2_X1 U1456 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1775), .ZN(n1834) );
NAND2_X1 U1457 ( .A1(n1836), .A2(n1837), .ZN(U295) );
NAND2_X1 U1458 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1776), .ZN(n1837) );
NAND2_X1 U1459 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1775), .ZN(n1836) );
NAND2_X1 U1460 ( .A1(n1838), .A2(n1839), .ZN(U294) );
NAND2_X1 U1461 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1776), .ZN(n1839) );
NAND2_X1 U1462 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1775), .ZN(n1838) );
NAND2_X1 U1463 ( .A1(n1840), .A2(n1841), .ZN(U293) );
NAND2_X1 U1464 ( .A1(n1842), .A2(n1776), .ZN(n1841) );
XNOR2_X1 U1465 ( .A(REG3_REG_4__SCAN_IN), .B(KEYINPUT46), .ZN(n1842) );
NAND2_X1 U1466 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1775), .ZN(n1840) );
NAND2_X1 U1467 ( .A1(n1843), .A2(n1844), .ZN(U292) );
NAND2_X1 U1468 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1845), .ZN(n1844) );
XOR2_X1 U1469 ( .A(KEYINPUT35), .B(n1776), .Z(n1845) );
NAND2_X1 U1470 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1775), .ZN(n1843) );
NAND2_X1 U1471 ( .A1(n1846), .A2(n1847), .ZN(U291) );
NAND2_X1 U1472 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1776), .ZN(n1847) );
NAND2_X1 U1473 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1775), .ZN(n1846) );
NAND2_X1 U1474 ( .A1(n1848), .A2(n1849), .ZN(U290) );
NAND2_X1 U1475 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1776), .ZN(n1849) );
NAND2_X1 U1476 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1775), .ZN(n1848) );
NAND2_X1 U1477 ( .A1(n1850), .A2(n1851), .ZN(U289) );
NAND2_X1 U1478 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1776), .ZN(n1851) );
NAND2_X1 U1479 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1775), .ZN(n1850) );
NAND4_X1 U1480 ( .A1(n1852), .A2(n1853), .A3(n1854), .A4(n1855), .ZN(U288));
NAND2_X1 U1481 ( .A1(n1856), .A2(REG4_REG_7__SCAN_IN), .ZN(n1854) );
NAND2_X1 U1482 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1857), .ZN(n1853) );
NAND2_X1 U1483 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1775), .ZN(n1852) );
NAND4_X1 U1484 ( .A1(n1858), .A2(n1855), .A3(n1859), .A4(n1860), .ZN(U287));
NOR3_X1 U1485 ( .A1(n1861), .A2(n1862), .A3(n1863), .ZN(n1860) );
NOR2_X1 U1486 ( .A1(n1864), .A2(n1865), .ZN(n1863) );
XOR2_X1 U1487 ( .A(REG4_REG_6__SCAN_IN), .B(KEYINPUT23), .Z(n1865) );
NOR3_X1 U1488 ( .A1(n1866), .A2(n1867), .A3(n1868), .ZN(n1862) );
INV_X1 U1489 ( .A(n1869), .ZN(n1867) );
XOR2_X1 U1490 ( .A(KEYINPUT26), .B(n1870), .Z(n1866) );
AND2_X1 U1491 ( .A1(n1857), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1861) );
NAND2_X1 U1492 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1775), .ZN(n1859) );
NAND2_X1 U1493 ( .A1(n1871), .A2(n1872), .ZN(n1855) );
NAND2_X1 U1494 ( .A1(n1873), .A2(n1874), .ZN(n1871) );
NAND3_X1 U1495 ( .A1(n1875), .A2(n1876), .A3(n1877), .ZN(n1874) );
NAND3_X1 U1496 ( .A1(n1878), .A2(n1879), .A3(n1880), .ZN(n1873) );
XNOR2_X1 U1497 ( .A(n1881), .B(KEYINPUT7), .ZN(n1880) );
XNOR2_X1 U1498 ( .A(KEYINPUT57), .B(n1882), .ZN(n1879) );
NAND3_X1 U1499 ( .A1(n1878), .A2(n1881), .A3(n1883), .ZN(n1858) );
NAND4_X1 U1500 ( .A1(n1884), .A2(n1885), .A3(n1886), .A4(n1887), .ZN(U286));
NOR3_X1 U1501 ( .A1(n1888), .A2(n1889), .A3(n1890), .ZN(n1887) );
NOR3_X1 U1502 ( .A1(n1868), .A2(n1870), .A3(n1891), .ZN(n1890) );
NOR2_X1 U1503 ( .A1(n1892), .A2(n1893), .ZN(n1891) );
INV_X1 U1504 ( .A(n1876), .ZN(n1870) );
NAND2_X1 U1505 ( .A1(n1894), .A2(n1892), .ZN(n1876) );
XOR2_X1 U1506 ( .A(n1893), .B(KEYINPUT40), .Z(n1894) );
NAND2_X1 U1507 ( .A1(n1869), .A2(n1895), .ZN(n1893) );
NAND2_X1 U1508 ( .A1(n1883), .A2(n1896), .ZN(n1895) );
INV_X1 U1509 ( .A(n1875), .ZN(n1896) );
NAND2_X1 U1510 ( .A1(n1875), .A2(n1872), .ZN(n1869) );
NOR3_X1 U1511 ( .A1(n1897), .A2(n1881), .A3(n1898), .ZN(n1889) );
NOR2_X1 U1512 ( .A1(n1899), .A2(n1900), .ZN(n1898) );
XOR2_X1 U1513 ( .A(n1901), .B(KEYINPUT44), .Z(n1900) );
AND2_X1 U1514 ( .A1(n1899), .A2(n1901), .ZN(n1881) );
XNOR2_X1 U1515 ( .A(n1902), .B(n1882), .ZN(n1901) );
OR2_X1 U1516 ( .A1(KEYINPUT57), .A2(n1883), .ZN(n1902) );
INV_X1 U1517 ( .A(n1872), .ZN(n1883) );
NOR2_X1 U1518 ( .A1(n1872), .A2(n1903), .ZN(n1888) );
NAND2_X1 U1519 ( .A1(n1904), .A2(n1905), .ZN(n1872) );
NAND3_X1 U1520 ( .A1(n1906), .A2(n1907), .A3(n1908), .ZN(n1905) );
XOR2_X1 U1521 ( .A(n1909), .B(n1910), .Z(n1908) );
NAND2_X1 U1522 ( .A1(n1911), .A2(n1912), .ZN(n1906) );
NAND3_X1 U1523 ( .A1(n1912), .A2(n1913), .A3(n1914), .ZN(n1904) );
XNOR2_X1 U1524 ( .A(n1910), .B(n1909), .ZN(n1914) );
NAND2_X1 U1525 ( .A1(n1915), .A2(n1916), .ZN(n1909) );
NAND2_X1 U1526 ( .A1(n1917), .A2(DATA_IN_6_), .ZN(n1916) );
NAND2_X1 U1527 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1915) );
AND2_X1 U1528 ( .A1(n1918), .A2(n1919), .ZN(n1910) );
NAND2_X1 U1529 ( .A1(n1917), .A2(REG4_REG_6__SCAN_IN), .ZN(n1919) );
NAND2_X1 U1530 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1918) );
NAND2_X1 U1531 ( .A1(n1920), .A2(n1921), .ZN(n1913) );
XNOR2_X1 U1532 ( .A(KEYINPUT6), .B(n1907), .ZN(n1920) );
OR2_X1 U1533 ( .A1(n1922), .A2(n1923), .ZN(n1907) );
NAND2_X1 U1534 ( .A1(n1922), .A2(n1923), .ZN(n1912) );
NAND2_X1 U1535 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1775), .ZN(n1886) );
NAND2_X1 U1536 ( .A1(n1856), .A2(REG4_REG_5__SCAN_IN), .ZN(n1885) );
NAND2_X1 U1537 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1857), .ZN(n1884) );
NAND4_X1 U1538 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .ZN(U285));
NOR3_X1 U1539 ( .A1(n1928), .A2(n1929), .A3(n1930), .ZN(n1927) );
NOR3_X1 U1540 ( .A1(n1868), .A2(n1892), .A3(n1931), .ZN(n1930) );
NOR2_X1 U1541 ( .A1(n1932), .A2(n1933), .ZN(n1931) );
AND2_X1 U1542 ( .A1(n1932), .A2(n1933), .ZN(n1892) );
NAND2_X1 U1543 ( .A1(n1934), .A2(n1935), .ZN(n1933) );
NAND2_X1 U1544 ( .A1(n1936), .A2(n1937), .ZN(n1935) );
XOR2_X1 U1545 ( .A(KEYINPUT54), .B(n1875), .Z(n1934) );
NOR2_X1 U1546 ( .A1(n1937), .A2(n1936), .ZN(n1875) );
NOR3_X1 U1547 ( .A1(n1897), .A2(n1899), .A3(n1938), .ZN(n1929) );
NOR2_X1 U1548 ( .A1(n1939), .A2(n1940), .ZN(n1938) );
AND2_X1 U1549 ( .A1(n1939), .A2(n1940), .ZN(n1899) );
NAND3_X1 U1550 ( .A1(n1941), .A2(n1942), .A3(n1882), .ZN(n1940) );
OR2_X1 U1551 ( .A1(n1943), .A2(n1936), .ZN(n1882) );
NAND3_X1 U1552 ( .A1(KEYINPUT4), .A2(n1936), .A3(n1943), .ZN(n1942) );
INV_X1 U1553 ( .A(n1944), .ZN(n1936) );
OR2_X1 U1554 ( .A1(n1943), .A2(KEYINPUT4), .ZN(n1941) );
NOR2_X1 U1555 ( .A1(n1944), .A2(n1945), .ZN(n1928) );
XOR2_X1 U1556 ( .A(KEYINPUT63), .B(n1946), .Z(n1945) );
XOR2_X1 U1557 ( .A(n1947), .B(n1922), .Z(n1944) );
AND2_X1 U1558 ( .A1(n1948), .A2(n1949), .ZN(n1922) );
NAND2_X1 U1559 ( .A1(RESTART), .A2(n1950), .ZN(n1949) );
XOR2_X1 U1560 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT61), .Z(n1950) );
NAND2_X1 U1561 ( .A1(n1917), .A2(DATA_IN_5_), .ZN(n1948) );
NAND2_X1 U1562 ( .A1(n1951), .A2(n1952), .ZN(n1947) );
NAND2_X1 U1563 ( .A1(n1911), .A2(n1923), .ZN(n1952) );
INV_X1 U1564 ( .A(n1921), .ZN(n1911) );
NAND2_X1 U1565 ( .A1(n1953), .A2(n1921), .ZN(n1951) );
NAND2_X1 U1566 ( .A1(n1954), .A2(n1955), .ZN(n1921) );
NAND2_X1 U1567 ( .A1(n1956), .A2(n1957), .ZN(n1955) );
NAND2_X1 U1568 ( .A1(n1958), .A2(n1959), .ZN(n1957) );
XOR2_X1 U1569 ( .A(n1960), .B(KEYINPUT62), .Z(n1958) );
OR2_X1 U1570 ( .A1(n1960), .A2(n1959), .ZN(n1954) );
NAND2_X1 U1571 ( .A1(KEYINPUT18), .A2(n1923), .ZN(n1953) );
AND2_X1 U1572 ( .A1(n1961), .A2(n1962), .ZN(n1923) );
NAND2_X1 U1573 ( .A1(n1917), .A2(REG4_REG_5__SCAN_IN), .ZN(n1962) );
NAND2_X1 U1574 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1961) );
NAND2_X1 U1575 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1775), .ZN(n1926) );
NAND2_X1 U1576 ( .A1(n1856), .A2(REG4_REG_4__SCAN_IN), .ZN(n1925) );
NAND2_X1 U1577 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1857), .ZN(n1924) );
NAND4_X1 U1578 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(U284));
NOR3_X1 U1579 ( .A1(n1967), .A2(n1968), .A3(n1969), .ZN(n1966) );
NOR3_X1 U1580 ( .A1(n1868), .A2(n1932), .A3(n1970), .ZN(n1969) );
NOR2_X1 U1581 ( .A1(n1971), .A2(n1972), .ZN(n1970) );
AND2_X1 U1582 ( .A1(n1971), .A2(n1972), .ZN(n1932) );
NAND2_X1 U1583 ( .A1(n1937), .A2(n1973), .ZN(n1972) );
NAND2_X1 U1584 ( .A1(n1974), .A2(n1975), .ZN(n1937) );
XOR2_X1 U1585 ( .A(n1976), .B(KEYINPUT17), .Z(n1974) );
NOR3_X1 U1586 ( .A1(n1897), .A2(n1939), .A3(n1977), .ZN(n1968) );
NOR2_X1 U1587 ( .A1(n1978), .A2(n1979), .ZN(n1977) );
AND2_X1 U1588 ( .A1(n1978), .A2(n1979), .ZN(n1939) );
NAND2_X1 U1589 ( .A1(n1943), .A2(n1973), .ZN(n1979) );
NAND2_X1 U1590 ( .A1(n1976), .A2(n1980), .ZN(n1973) );
NAND2_X1 U1591 ( .A1(n1975), .A2(n1981), .ZN(n1943) );
NOR2_X1 U1592 ( .A1(n1981), .A2(n1903), .ZN(n1967) );
INV_X1 U1593 ( .A(n1976), .ZN(n1981) );
NAND3_X1 U1594 ( .A1(n1982), .A2(n1983), .A3(n1984), .ZN(n1976) );
NAND2_X1 U1595 ( .A1(n1959), .A2(n1985), .ZN(n1984) );
NAND3_X1 U1596 ( .A1(n1986), .A2(n1987), .A3(KEYINPUT21), .ZN(n1985) );
NAND2_X1 U1597 ( .A1(KEYINPUT34), .A2(n1988), .ZN(n1987) );
OR3_X1 U1598 ( .A1(n1960), .A2(n1956), .A3(KEYINPUT34), .ZN(n1986) );
INV_X1 U1599 ( .A(n1989), .ZN(n1959) );
NAND3_X1 U1600 ( .A1(KEYINPUT21), .A2(n1989), .A3(n1990), .ZN(n1983) );
NAND2_X1 U1601 ( .A1(n1991), .A2(n1992), .ZN(n1989) );
NAND2_X1 U1602 ( .A1(n1993), .A2(n1994), .ZN(n1992) );
OR2_X1 U1603 ( .A1(n1995), .A2(n1996), .ZN(n1994) );
NAND2_X1 U1604 ( .A1(n1996), .A2(n1995), .ZN(n1991) );
OR2_X1 U1605 ( .A1(n1990), .A2(KEYINPUT21), .ZN(n1982) );
INV_X1 U1606 ( .A(n1988), .ZN(n1990) );
XOR2_X1 U1607 ( .A(n1956), .B(n1960), .Z(n1988) );
NAND2_X1 U1608 ( .A1(n1997), .A2(n1998), .ZN(n1960) );
NAND2_X1 U1609 ( .A1(n1917), .A2(DATA_IN_4_), .ZN(n1998) );
NAND2_X1 U1610 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1997) );
AND2_X1 U1611 ( .A1(n1999), .A2(n2000), .ZN(n1956) );
NAND2_X1 U1612 ( .A1(REG4_REG_4__SCAN_IN), .A2(n2001), .ZN(n2000) );
XOR2_X1 U1613 ( .A(KEYINPUT50), .B(n2002), .Z(n2001) );
NAND2_X1 U1614 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n1999) );
NAND2_X1 U1615 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1775), .ZN(n1965) );
NAND2_X1 U1616 ( .A1(n1856), .A2(REG4_REG_3__SCAN_IN), .ZN(n1964) );
NAND2_X1 U1617 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1857), .ZN(n1963) );
NAND4_X1 U1618 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .ZN(U283));
NOR3_X1 U1619 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n2006) );
XOR2_X1 U1620 ( .A(KEYINPUT25), .B(n2010), .Z(n2009) );
NOR2_X1 U1621 ( .A1(n2011), .A2(n1864), .ZN(n2010) );
XOR2_X1 U1622 ( .A(KEYINPUT47), .B(n2012), .Z(n2008) );
NOR3_X1 U1623 ( .A1(n1868), .A2(n1971), .A3(n2013), .ZN(n2012) );
NOR2_X1 U1624 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
AND2_X1 U1625 ( .A1(n2016), .A2(n2017), .ZN(n2014) );
AND3_X1 U1626 ( .A1(n2015), .A2(n2016), .A3(n2018), .ZN(n1971) );
XNOR2_X1 U1627 ( .A(KEYINPUT31), .B(n2017), .ZN(n2018) );
XOR2_X1 U1628 ( .A(KEYINPUT51), .B(n2019), .Z(n2007) );
NOR3_X1 U1629 ( .A1(n1897), .A2(n1978), .A3(n2020), .ZN(n2019) );
NOR2_X1 U1630 ( .A1(n2021), .A2(n2015), .ZN(n2020) );
XOR2_X1 U1631 ( .A(n2022), .B(KEYINPUT29), .Z(n2021) );
NAND2_X1 U1632 ( .A1(n2017), .A2(n2023), .ZN(n2022) );
AND3_X1 U1633 ( .A1(n2017), .A2(n2015), .A3(n2023), .ZN(n1978) );
NAND2_X1 U1634 ( .A1(n1980), .A2(n2024), .ZN(n2015) );
NAND2_X1 U1635 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
INV_X1 U1636 ( .A(n1975), .ZN(n1980) );
NOR2_X1 U1637 ( .A1(n2026), .A2(n2025), .ZN(n1975) );
NAND2_X1 U1638 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1775), .ZN(n2005) );
NAND2_X1 U1639 ( .A1(n1946), .A2(n2025), .ZN(n2004) );
NAND2_X1 U1640 ( .A1(n2027), .A2(n2028), .ZN(n2025) );
NAND2_X1 U1641 ( .A1(n2029), .A2(n2030), .ZN(n2028) );
NAND2_X1 U1642 ( .A1(KEYINPUT20), .A2(n1995), .ZN(n2030) );
XOR2_X1 U1643 ( .A(n1996), .B(n2031), .Z(n2029) );
NAND3_X1 U1644 ( .A1(n2032), .A2(n2033), .A3(n1995), .ZN(n2027) );
NAND2_X1 U1645 ( .A1(n2034), .A2(n2035), .ZN(n1995) );
NAND2_X1 U1646 ( .A1(n2036), .A2(n2037), .ZN(n2035) );
NAND2_X1 U1647 ( .A1(n2038), .A2(n2039), .ZN(n2036) );
OR2_X1 U1648 ( .A1(n2038), .A2(n2039), .ZN(n2034) );
NAND2_X1 U1649 ( .A1(n1996), .A2(n1993), .ZN(n2033) );
INV_X1 U1650 ( .A(n2031), .ZN(n1993) );
NAND2_X1 U1651 ( .A1(n2040), .A2(n2031), .ZN(n2032) );
NAND2_X1 U1652 ( .A1(n2041), .A2(n2042), .ZN(n2031) );
NAND2_X1 U1653 ( .A1(n2043), .A2(DATA_IN_3_), .ZN(n2042) );
XOR2_X1 U1654 ( .A(n1917), .B(KEYINPUT14), .Z(n2043) );
NAND2_X1 U1655 ( .A1(RESTART), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2041) );
NAND2_X1 U1656 ( .A1(KEYINPUT20), .A2(n1996), .ZN(n2040) );
AND2_X1 U1657 ( .A1(n2044), .A2(n2045), .ZN(n1996) );
NAND2_X1 U1658 ( .A1(n1917), .A2(REG4_REG_3__SCAN_IN), .ZN(n2045) );
XOR2_X1 U1659 ( .A(n2046), .B(KEYINPUT32), .Z(n2044) );
NAND2_X1 U1660 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2046) );
NAND2_X1 U1661 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1857), .ZN(n2003) );
NAND4_X1 U1662 ( .A1(n2047), .A2(n2048), .A3(n2049), .A4(n2050), .ZN(U282));
NOR3_X1 U1663 ( .A1(n2051), .A2(n2052), .A3(n2053), .ZN(n2050) );
NOR2_X1 U1664 ( .A1(n2054), .A2(n1897), .ZN(n2053) );
INV_X1 U1665 ( .A(n1878), .ZN(n1897) );
NOR2_X1 U1666 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
XOR2_X1 U1667 ( .A(n2057), .B(KEYINPUT5), .Z(n2056) );
NAND2_X1 U1668 ( .A1(n2058), .A2(n2017), .ZN(n2057) );
NOR2_X1 U1669 ( .A1(n2058), .A2(n2017), .ZN(n2055) );
INV_X1 U1670 ( .A(n2023), .ZN(n2058) );
NAND2_X1 U1671 ( .A1(n2026), .A2(n2059), .ZN(n2023) );
NAND2_X1 U1672 ( .A1(n2060), .A2(n2061), .ZN(n2059) );
NOR2_X1 U1673 ( .A1(n2062), .A2(n2063), .ZN(n2052) );
XOR2_X1 U1674 ( .A(n1868), .B(KEYINPUT38), .Z(n2063) );
XNOR2_X1 U1675 ( .A(n2016), .B(n2017), .ZN(n2062) );
NAND3_X1 U1676 ( .A1(n2064), .A2(n2065), .A3(n2026), .ZN(n2016) );
OR2_X1 U1677 ( .A1(n2061), .A2(n2060), .ZN(n2026) );
NAND3_X1 U1678 ( .A1(n2060), .A2(n2061), .A3(n2066), .ZN(n2065) );
OR2_X1 U1679 ( .A1(n2066), .A2(n2061), .ZN(n2064) );
INV_X1 U1680 ( .A(KEYINPUT8), .ZN(n2066) );
AND2_X1 U1681 ( .A1(n2060), .A2(n1946), .ZN(n2051) );
INV_X1 U1682 ( .A(n1903), .ZN(n1946) );
XNOR2_X1 U1683 ( .A(n2037), .B(n2067), .ZN(n2060) );
XOR2_X1 U1684 ( .A(n2038), .B(n2039), .Z(n2067) );
NAND2_X1 U1685 ( .A1(n2068), .A2(n2069), .ZN(n2039) );
NAND2_X1 U1686 ( .A1(n1917), .A2(REG4_REG_2__SCAN_IN), .ZN(n2069) );
NAND2_X1 U1687 ( .A1(RESTART), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2068) );
NAND2_X1 U1688 ( .A1(n2070), .A2(n2071), .ZN(n2038) );
NAND2_X1 U1689 ( .A1(n1917), .A2(DATA_IN_2_), .ZN(n2071) );
NAND2_X1 U1690 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2070) );
NAND2_X1 U1691 ( .A1(n2072), .A2(n2073), .ZN(n2037) );
NAND2_X1 U1692 ( .A1(n2074), .A2(n2075), .ZN(n2073) );
NAND2_X1 U1693 ( .A1(n2076), .A2(n2077), .ZN(n2075) );
XOR2_X1 U1694 ( .A(KEYINPUT59), .B(n2078), .Z(n2074) );
OR2_X1 U1695 ( .A1(n2079), .A2(n2076), .ZN(n2072) );
NAND2_X1 U1696 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1775), .ZN(n2049) );
NAND2_X1 U1697 ( .A1(n1856), .A2(REG4_REG_1__SCAN_IN), .ZN(n2048) );
NAND2_X1 U1698 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1857), .ZN(n2047) );
NAND3_X1 U1699 ( .A1(n2080), .A2(n2081), .A3(n2082), .ZN(U281) );
NOR3_X1 U1700 ( .A1(n2083), .A2(n2084), .A3(n2085), .ZN(n2082) );
NOR2_X1 U1701 ( .A1(n2086), .A2(n2087), .ZN(n2085) );
XOR2_X1 U1702 ( .A(n1864), .B(KEYINPUT30), .Z(n2086) );
INV_X1 U1703 ( .A(n1856), .ZN(n1864) );
NOR2_X1 U1704 ( .A1(n2088), .A2(n2089), .ZN(n1856) );
NOR2_X1 U1705 ( .A1(n2090), .A2(n2017), .ZN(n2084) );
NAND2_X1 U1706 ( .A1(n2061), .A2(n2091), .ZN(n2017) );
NAND3_X1 U1707 ( .A1(n2092), .A2(n2093), .A3(n2094), .ZN(n2091) );
NAND2_X1 U1708 ( .A1(n2095), .A2(n2096), .ZN(n2061) );
NAND2_X1 U1709 ( .A1(n2093), .A2(n2094), .ZN(n2096) );
NAND2_X1 U1710 ( .A1(n2097), .A2(n2098), .ZN(n2094) );
NAND2_X1 U1711 ( .A1(n1917), .A2(n2099), .ZN(n2098) );
NAND2_X1 U1712 ( .A1(n2087), .A2(n1744), .ZN(n2099) );
NAND2_X1 U1713 ( .A1(RESTART), .A2(n2100), .ZN(n2097) );
NAND2_X1 U1714 ( .A1(n2101), .A2(n1712), .ZN(n2100) );
NOR2_X1 U1715 ( .A1(n1878), .A2(n1877), .ZN(n2090) );
INV_X1 U1716 ( .A(n1868), .ZN(n1877) );
NAND3_X1 U1717 ( .A1(RESTART), .A2(n2102), .A3(n2103), .ZN(n1868) );
NOR3_X1 U1718 ( .A1(n2104), .A2(AVERAGE), .A3(n2089), .ZN(n1878) );
NOR2_X1 U1719 ( .A1(n2095), .A2(n1903), .ZN(n2083) );
NAND3_X1 U1720 ( .A1(n2105), .A2(n2106), .A3(n2103), .ZN(n1903) );
NAND2_X1 U1721 ( .A1(n1917), .A2(n2107), .ZN(n2106) );
NAND3_X1 U1722 ( .A1(n2104), .A2(n2088), .A3(ENABLE), .ZN(n2107) );
INV_X1 U1723 ( .A(AVERAGE), .ZN(n2088) );
NAND2_X1 U1724 ( .A1(n2108), .A2(n2109), .ZN(n2104) );
NAND2_X1 U1725 ( .A1(n2110), .A2(n2111), .ZN(n2109) );
INV_X1 U1726 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2111) );
OR2_X1 U1727 ( .A1(n2112), .A2(n1723), .ZN(n2110) );
NAND2_X1 U1728 ( .A1(n2112), .A2(n1723), .ZN(n2108) );
INV_X1 U1729 ( .A(DATA_IN_7_), .ZN(n1723) );
NAND2_X1 U1730 ( .A1(n2113), .A2(n2114), .ZN(n2112) );
NAND2_X1 U1731 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2115), .ZN(n2114) );
OR2_X1 U1732 ( .A1(n2116), .A2(DATA_IN_6_), .ZN(n2115) );
NAND2_X1 U1733 ( .A1(DATA_IN_6_), .A2(n2116), .ZN(n2113) );
NAND3_X1 U1734 ( .A1(n2117), .A2(n2118), .A3(n2119), .ZN(n2116) );
NAND2_X1 U1735 ( .A1(DATA_IN_5_), .A2(n2120), .ZN(n2119) );
NAND2_X1 U1736 ( .A1(KEYINPUT15), .A2(n2121), .ZN(n2118) );
NAND2_X1 U1737 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2121) );
NAND2_X1 U1738 ( .A1(REG4_REG_5__SCAN_IN), .A2(n2122), .ZN(n2117) );
NAND2_X1 U1739 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
OR2_X1 U1740 ( .A1(n1698), .A2(KEYINPUT15), .ZN(n2124) );
INV_X1 U1741 ( .A(DATA_IN_5_), .ZN(n1698) );
INV_X1 U1742 ( .A(n2120), .ZN(n2123) );
NAND2_X1 U1743 ( .A1(n2125), .A2(n2126), .ZN(n2120) );
NAND2_X1 U1744 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2126) );
NAND3_X1 U1745 ( .A1(n2127), .A2(n2128), .A3(n2129), .ZN(n2125) );
XOR2_X1 U1746 ( .A(KEYINPUT24), .B(n2130), .Z(n2129) );
NOR3_X1 U1747 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n2130) );
NOR2_X1 U1748 ( .A1(n1716), .A2(n2134), .ZN(n2133) );
NOR3_X1 U1749 ( .A1(n2135), .A2(n2136), .A3(n2137), .ZN(n2132) );
NOR2_X1 U1750 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2137) );
NOR2_X1 U1751 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2136) );
NOR2_X1 U1752 ( .A1(n2138), .A2(n2139), .ZN(n2135) );
AND2_X1 U1753 ( .A1(DATA_IN_1_), .A2(REG4_REG_1__SCAN_IN), .ZN(n2139) );
NOR2_X1 U1754 ( .A1(n1744), .A2(n2087), .ZN(n2138) );
NOR2_X1 U1755 ( .A1(n1710), .A2(n2011), .ZN(n2131) );
INV_X1 U1756 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2011) );
INV_X1 U1757 ( .A(DATA_IN_2_), .ZN(n1710) );
NAND2_X1 U1758 ( .A1(n1716), .A2(n2134), .ZN(n2128) );
INV_X1 U1759 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2134) );
INV_X1 U1760 ( .A(DATA_IN_3_), .ZN(n1716) );
OR2_X1 U1761 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2127) );
NAND2_X1 U1762 ( .A1(RESTART), .A2(n2102), .ZN(n2105) );
NAND2_X1 U1763 ( .A1(n2140), .A2(n2141), .ZN(n2102) );
NAND2_X1 U1764 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2141) );
XOR2_X1 U1765 ( .A(n2142), .B(KEYINPUT55), .Z(n2140) );
NAND3_X1 U1766 ( .A1(n2143), .A2(n2144), .A3(n2145), .ZN(n2142) );
OR2_X1 U1767 ( .A1(RMAX_REG_7__SCAN_IN), .A2(RMIN_REG_7__SCAN_IN), .ZN(n2145) );
NAND2_X1 U1768 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2146), .ZN(n2144) );
OR2_X1 U1769 ( .A1(n2147), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2146) );
NAND2_X1 U1770 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2147), .ZN(n2143) );
NAND2_X1 U1771 ( .A1(n2148), .A2(n2149), .ZN(n2147) );
NAND2_X1 U1772 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n2150), .ZN(n2149) );
OR2_X1 U1773 ( .A1(n2151), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2150) );
NAND2_X1 U1774 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2151), .ZN(n2148) );
NAND2_X1 U1775 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
NAND3_X1 U1776 ( .A1(n2154), .A2(n2155), .A3(n2156), .ZN(n2153) );
NAND2_X1 U1777 ( .A1(n1702), .A2(n1748), .ZN(n2156) );
NAND3_X1 U1778 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n2155) );
XOR2_X1 U1779 ( .A(KEYINPUT56), .B(n2160), .Z(n2159) );
NOR2_X1 U1780 ( .A1(n1717), .A2(n1739), .ZN(n2160) );
NAND3_X1 U1781 ( .A1(n2161), .A2(n2162), .A3(n2163), .ZN(n2158) );
OR2_X1 U1782 ( .A1(RMAX_REG_2__SCAN_IN), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2163) );
NAND2_X1 U1783 ( .A1(n2164), .A2(n1745), .ZN(n2162) );
OR2_X1 U1784 ( .A1(n2165), .A2(n1714), .ZN(n2164) );
NAND2_X1 U1785 ( .A1(n2165), .A2(n1714), .ZN(n2161) );
INV_X1 U1786 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1714) );
NAND2_X1 U1787 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2157) );
NAND2_X1 U1788 ( .A1(n1717), .A2(n1739), .ZN(n2154) );
INV_X1 U1789 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1739) );
INV_X1 U1790 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1717) );
XOR2_X1 U1791 ( .A(KEYINPUT1), .B(n2166), .Z(n2152) );
NOR2_X1 U1792 ( .A1(n1702), .A2(n1748), .ZN(n2166) );
INV_X1 U1793 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1748) );
INV_X1 U1794 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1702) );
INV_X1 U1795 ( .A(n2092), .ZN(n2095) );
NAND2_X1 U1796 ( .A1(n2167), .A2(n2168), .ZN(n2092) );
NAND2_X1 U1797 ( .A1(n2169), .A2(n2077), .ZN(n2168) );
XOR2_X1 U1798 ( .A(KEYINPUT33), .B(n2170), .Z(n2167) );
NOR2_X1 U1799 ( .A1(n2079), .A2(n2169), .ZN(n2170) );
XOR2_X1 U1800 ( .A(n2076), .B(n2078), .Z(n2169) );
AND2_X1 U1801 ( .A1(n2171), .A2(n2172), .ZN(n2078) );
NAND2_X1 U1802 ( .A1(n1917), .A2(REG4_REG_1__SCAN_IN), .ZN(n2172) );
XOR2_X1 U1803 ( .A(KEYINPUT28), .B(n2173), .Z(n2171) );
NOR2_X1 U1804 ( .A1(n1745), .A2(n2174), .ZN(n2173) );
INV_X1 U1805 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1745) );
INV_X1 U1806 ( .A(n2093), .ZN(n2076) );
NAND4_X1 U1807 ( .A1(n2175), .A2(n2176), .A3(n2177), .A4(n2178), .ZN(n2093));
NAND2_X1 U1808 ( .A1(n2179), .A2(n2174), .ZN(n2178) );
NAND3_X1 U1809 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .A3(n1917), .ZN(n2179) );
NAND2_X1 U1810 ( .A1(n2002), .A2(n2165), .ZN(n2177) );
NAND2_X1 U1811 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2165) );
NAND2_X1 U1812 ( .A1(n1744), .A2(n1712), .ZN(n2176) );
INV_X1 U1813 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1712) );
INV_X1 U1814 ( .A(DATA_IN_0_), .ZN(n1744) );
NAND2_X1 U1815 ( .A1(n2087), .A2(n2101), .ZN(n2175) );
INV_X1 U1816 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2101) );
INV_X1 U1817 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2087) );
XNOR2_X1 U1818 ( .A(n2077), .B(KEYINPUT37), .ZN(n2079) );
NAND2_X1 U1819 ( .A1(n2180), .A2(n2181), .ZN(n2077) );
NAND2_X1 U1820 ( .A1(n1917), .A2(DATA_IN_1_), .ZN(n2181) );
NAND2_X1 U1821 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2180) );
NAND2_X1 U1822 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1857), .ZN(n2081) );
NAND2_X1 U1823 ( .A1(n2182), .A2(n2183), .ZN(n1857) );
NAND3_X1 U1824 ( .A1(n2184), .A2(n1770), .A3(n2185), .ZN(n2183) );
INV_X1 U1825 ( .A(ENABLE), .ZN(n1770) );
OR2_X1 U1826 ( .A1(n2185), .A2(n2089), .ZN(n2182) );
NAND2_X1 U1827 ( .A1(ENABLE), .A2(n2184), .ZN(n2089) );
AND2_X1 U1828 ( .A1(n2103), .A2(n2186), .ZN(n2184) );
XOR2_X1 U1829 ( .A(KEYINPUT58), .B(n2002), .Z(n2186) );
INV_X1 U1830 ( .A(n1917), .ZN(n2002) );
INV_X1 U1831 ( .A(RESTART), .ZN(n2174) );
NOR2_X1 U1832 ( .A1(n1771), .A2(n1775), .ZN(n2103) );
INV_X1 U1833 ( .A(KEYINPUT9), .ZN(n2185) );
NAND2_X1 U1834 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1775), .ZN(n2080) );
NAND2_X1 U1835 ( .A1(n1790), .A2(n2187), .ZN(U280) );
NAND2_X1 U1836 ( .A1(n2188), .A2(STATO_REG_0__SCAN_IN), .ZN(n2187) );
XOR2_X1 U1837 ( .A(n1771), .B(KEYINPUT36), .Z(n2188) );
INV_X1 U1838 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1771) );
NAND2_X1 U1839 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1663), .ZN(n1790) );
INV_X1 U1840 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1663) );
endmodule


