//Key = 0100101001000011101001010011110010110110011110100000010100101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337;

XOR2_X1 U735 ( .A(n1012), .B(n1013), .Z(G9) );
XNOR2_X1 U736 ( .A(KEYINPUT2), .B(n1014), .ZN(n1013) );
NOR2_X1 U737 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NOR3_X1 U739 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR3_X1 U741 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
XOR2_X1 U742 ( .A(n1028), .B(KEYINPUT54), .Z(n1027) );
XNOR2_X1 U743 ( .A(n1029), .B(KEYINPUT40), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1023) );
NAND3_X1 U745 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1017) );
NAND3_X1 U746 ( .A1(n1035), .A2(n1036), .A3(n1029), .ZN(n1034) );
INV_X1 U747 ( .A(n1031), .ZN(n1029) );
NAND2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1037) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U753 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1045) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
AND3_X1 U758 ( .A1(n1032), .A2(n1033), .A3(n1058), .ZN(n1015) );
NAND4_X1 U759 ( .A1(n1059), .A2(n1054), .A3(n1060), .A4(n1061), .ZN(n1032) );
NOR3_X1 U760 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
XNOR2_X1 U761 ( .A(n1065), .B(n1066), .ZN(n1064) );
NAND2_X1 U762 ( .A1(KEYINPUT9), .A2(n1067), .ZN(n1065) );
XOR2_X1 U763 ( .A(n1068), .B(n1069), .Z(n1063) );
NOR2_X1 U764 ( .A1(n1070), .A2(KEYINPUT31), .ZN(n1069) );
XNOR2_X1 U765 ( .A(n1071), .B(G478), .ZN(n1060) );
XNOR2_X1 U766 ( .A(n1072), .B(n1073), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(G72) );
NAND2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U769 ( .A1(G953), .A2(n1078), .ZN(n1077) );
NAND3_X1 U770 ( .A1(G953), .A2(n1079), .A3(n1080), .ZN(n1074) );
INV_X1 U771 ( .A(n1076), .ZN(n1080) );
XNOR2_X1 U772 ( .A(n1081), .B(n1082), .ZN(n1076) );
NOR3_X1 U773 ( .A1(n1083), .A2(KEYINPUT56), .A3(G953), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U775 ( .A(n1086), .B(KEYINPUT3), .Z(n1084) );
NAND2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
NAND2_X1 U777 ( .A1(G953), .A2(n1089), .ZN(n1088) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1087) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U780 ( .A(n1094), .B(KEYINPUT45), .Z(n1090) );
NAND3_X1 U781 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
NAND2_X1 U782 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
OR3_X1 U783 ( .A1(n1099), .A2(n1100), .A3(G134), .ZN(n1096) );
INV_X1 U784 ( .A(KEYINPUT42), .ZN(n1099) );
NAND2_X1 U785 ( .A1(G134), .A2(n1100), .ZN(n1095) );
NAND2_X1 U786 ( .A1(KEYINPUT53), .A2(n1101), .ZN(n1100) );
NAND2_X1 U787 ( .A1(G900), .A2(G227), .ZN(n1079) );
XOR2_X1 U788 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U789 ( .A1(n1104), .A2(n1033), .ZN(n1103) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U791 ( .A(KEYINPUT27), .B(n1107), .ZN(n1106) );
INV_X1 U792 ( .A(G224), .ZN(n1105) );
NOR3_X1 U793 ( .A1(KEYINPUT17), .A2(n1108), .A3(n1109), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
INV_X1 U796 ( .A(n1114), .ZN(n1113) );
NOR2_X1 U797 ( .A1(G898), .A2(n1033), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
INV_X1 U799 ( .A(n1111), .ZN(n1116) );
NOR2_X1 U800 ( .A1(G953), .A2(n1114), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NOR2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XNOR2_X1 U803 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1125), .ZN(G63) );
NOR3_X1 U806 ( .A1(n1071), .A2(n1126), .A3(n1127), .ZN(n1125) );
AND3_X1 U807 ( .A1(n1128), .A2(G478), .A3(n1129), .ZN(n1127) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1128), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1133), .ZN(G60) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U812 ( .A1(n1129), .A2(G475), .ZN(n1135) );
NAND2_X1 U813 ( .A1(KEYINPUT23), .A2(n1136), .ZN(n1134) );
XOR2_X1 U814 ( .A(n1137), .B(n1138), .Z(G6) );
NAND2_X1 U815 ( .A1(KEYINPUT15), .A2(n1139), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1119), .A2(n1140), .ZN(G57) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1141) );
NOR2_X1 U820 ( .A1(n1067), .A2(n1124), .ZN(n1146) );
NAND2_X1 U821 ( .A1(KEYINPUT55), .A2(n1147), .ZN(n1145) );
NOR3_X1 U822 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(G54) );
AND2_X1 U823 ( .A1(KEYINPUT41), .A2(n1119), .ZN(n1150) );
NOR3_X1 U824 ( .A1(KEYINPUT41), .A2(n1033), .A3(n1058), .ZN(n1149) );
INV_X1 U825 ( .A(G952), .ZN(n1058) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1148) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND3_X1 U829 ( .A1(n1157), .A2(n1019), .A3(G469), .ZN(n1156) );
INV_X1 U830 ( .A(n1131), .ZN(n1019) );
XNOR2_X1 U831 ( .A(KEYINPUT51), .B(n1158), .ZN(n1157) );
NAND3_X1 U832 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1155) );
NAND2_X1 U833 ( .A1(n1092), .A2(n1162), .ZN(n1161) );
OR3_X1 U834 ( .A1(n1162), .A2(n1092), .A3(n1163), .ZN(n1160) );
INV_X1 U835 ( .A(KEYINPUT34), .ZN(n1162) );
NAND2_X1 U836 ( .A1(n1163), .A2(n1164), .ZN(n1159) );
NAND2_X1 U837 ( .A1(KEYINPUT34), .A2(n1165), .ZN(n1164) );
XOR2_X1 U838 ( .A(KEYINPUT16), .B(n1092), .Z(n1165) );
XOR2_X1 U839 ( .A(n1166), .B(n1167), .Z(n1151) );
NOR2_X1 U840 ( .A1(G140), .A2(KEYINPUT47), .ZN(n1167) );
XOR2_X1 U841 ( .A(n1168), .B(KEYINPUT46), .Z(n1166) );
NOR2_X1 U842 ( .A1(n1119), .A2(n1169), .ZN(G51) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1124), .ZN(n1172) );
INV_X1 U846 ( .A(n1129), .ZN(n1124) );
NOR2_X1 U847 ( .A1(n1158), .A2(n1131), .ZN(n1129) );
NOR4_X1 U848 ( .A1(n1175), .A2(n1086), .A3(n1117), .A4(n1085), .ZN(n1131) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1085) );
NOR4_X1 U850 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
AND2_X1 U851 ( .A1(n1183), .A2(KEYINPUT14), .ZN(n1182) );
NOR3_X1 U852 ( .A1(KEYINPUT14), .A2(n1184), .A3(n1030), .ZN(n1181) );
NOR4_X1 U853 ( .A1(n1185), .A2(n1050), .A3(n1042), .A4(n1186), .ZN(n1184) );
AND2_X1 U854 ( .A1(KEYINPUT21), .A2(n1187), .ZN(n1180) );
NOR3_X1 U855 ( .A1(KEYINPUT21), .A2(n1188), .A3(n1189), .ZN(n1179) );
NAND4_X1 U856 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1117) );
NOR4_X1 U857 ( .A1(n1138), .A2(n1194), .A3(n1012), .A4(n1195), .ZN(n1193) );
INV_X1 U858 ( .A(n1196), .ZN(n1195) );
AND2_X1 U859 ( .A1(n1197), .A2(n1198), .ZN(n1012) );
INV_X1 U860 ( .A(n1199), .ZN(n1194) );
AND2_X1 U861 ( .A1(n1200), .A2(n1198), .ZN(n1138) );
AND4_X1 U862 ( .A1(n1201), .A2(n1202), .A3(n1049), .A4(n1047), .ZN(n1198) );
OR2_X1 U863 ( .A1(n1203), .A2(n1030), .ZN(n1192) );
NAND3_X1 U864 ( .A1(n1204), .A2(n1202), .A3(n1039), .ZN(n1190) );
NAND4_X1 U865 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1086) );
OR4_X1 U866 ( .A1(n1209), .A2(n1204), .A3(n1057), .A4(KEYINPUT28), .ZN(n1208) );
NAND2_X1 U867 ( .A1(n1210), .A2(KEYINPUT28), .ZN(n1207) );
NAND2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U870 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U871 ( .A(KEYINPUT30), .B(n1041), .ZN(n1216) );
NAND2_X1 U872 ( .A1(n1043), .A2(n1217), .ZN(n1213) );
XOR2_X1 U873 ( .A(n1118), .B(KEYINPUT63), .Z(n1175) );
XOR2_X1 U874 ( .A(n1218), .B(KEYINPUT19), .Z(n1170) );
NOR2_X1 U875 ( .A1(n1033), .A2(G952), .ZN(n1119) );
XOR2_X1 U876 ( .A(G146), .B(n1219), .Z(G48) );
NOR3_X1 U877 ( .A1(n1186), .A2(n1041), .A3(n1209), .ZN(n1219) );
XNOR2_X1 U878 ( .A(n1220), .B(n1210), .ZN(G45) );
NOR3_X1 U879 ( .A1(n1221), .A2(n1209), .A3(n1057), .ZN(n1210) );
XNOR2_X1 U880 ( .A(G140), .B(n1206), .ZN(G42) );
NAND3_X1 U881 ( .A1(n1217), .A2(n1200), .A3(n1188), .ZN(n1206) );
XOR2_X1 U882 ( .A(G137), .B(n1222), .Z(G39) );
NOR3_X1 U883 ( .A1(n1223), .A2(n1022), .A3(n1186), .ZN(n1222) );
INV_X1 U884 ( .A(n1043), .ZN(n1022) );
NAND3_X1 U885 ( .A1(n1201), .A2(n1224), .A3(n1035), .ZN(n1223) );
XNOR2_X1 U886 ( .A(KEYINPUT38), .B(n1225), .ZN(n1224) );
XNOR2_X1 U887 ( .A(G134), .B(n1176), .ZN(G36) );
NAND3_X1 U888 ( .A1(n1217), .A2(n1197), .A3(n1226), .ZN(n1176) );
XNOR2_X1 U889 ( .A(G131), .B(n1177), .ZN(G33) );
NAND3_X1 U890 ( .A1(n1217), .A2(n1200), .A3(n1226), .ZN(n1177) );
NOR3_X1 U891 ( .A1(n1050), .A2(n1185), .A3(n1062), .ZN(n1217) );
INV_X1 U892 ( .A(n1035), .ZN(n1062) );
NOR2_X1 U893 ( .A1(n1025), .A2(n1227), .ZN(n1035) );
INV_X1 U894 ( .A(n1028), .ZN(n1227) );
NAND2_X1 U895 ( .A1(n1228), .A2(n1229), .ZN(G30) );
NAND2_X1 U896 ( .A1(n1183), .A2(n1230), .ZN(n1229) );
XOR2_X1 U897 ( .A(n1231), .B(KEYINPUT8), .Z(n1228) );
OR2_X1 U898 ( .A1(n1230), .A2(n1183), .ZN(n1231) );
NOR3_X1 U899 ( .A1(n1209), .A2(n1042), .A3(n1186), .ZN(n1183) );
INV_X1 U900 ( .A(n1197), .ZN(n1042) );
INV_X1 U901 ( .A(n1215), .ZN(n1209) );
NOR3_X1 U902 ( .A1(n1030), .A2(n1185), .A3(n1050), .ZN(n1215) );
INV_X1 U903 ( .A(n1201), .ZN(n1050) );
INV_X1 U904 ( .A(n1225), .ZN(n1185) );
NAND2_X1 U905 ( .A1(n1232), .A2(n1233), .ZN(G3) );
OR2_X1 U906 ( .A1(n1191), .A2(G101), .ZN(n1233) );
XOR2_X1 U907 ( .A(n1234), .B(KEYINPUT0), .Z(n1232) );
NAND2_X1 U908 ( .A1(G101), .A2(n1191), .ZN(n1234) );
NAND4_X1 U909 ( .A1(n1226), .A2(n1043), .A3(n1201), .A4(n1202), .ZN(n1191) );
XOR2_X1 U910 ( .A(G125), .B(n1187), .Z(G27) );
NOR2_X1 U911 ( .A1(n1189), .A2(n1056), .ZN(n1187) );
NAND4_X1 U912 ( .A1(n1200), .A2(n1054), .A3(n1235), .A4(n1225), .ZN(n1189) );
NAND2_X1 U913 ( .A1(n1236), .A2(n1031), .ZN(n1225) );
NAND4_X1 U914 ( .A1(G953), .A2(G902), .A3(n1237), .A4(n1089), .ZN(n1236) );
INV_X1 U915 ( .A(G900), .ZN(n1089) );
XNOR2_X1 U916 ( .A(G122), .B(n1238), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1039), .A2(n1204), .A3(n1239), .A4(n1240), .ZN(n1238) );
XNOR2_X1 U918 ( .A(KEYINPUT22), .B(n1030), .ZN(n1239) );
INV_X1 U919 ( .A(n1221), .ZN(n1204) );
NAND2_X1 U920 ( .A1(n1241), .A2(n1242), .ZN(n1221) );
INV_X1 U921 ( .A(n1020), .ZN(n1039) );
NAND3_X1 U922 ( .A1(n1049), .A2(n1047), .A3(n1054), .ZN(n1020) );
XOR2_X1 U923 ( .A(n1243), .B(KEYINPUT5), .Z(n1049) );
XNOR2_X1 U924 ( .A(G119), .B(n1244), .ZN(G21) );
NAND2_X1 U925 ( .A1(KEYINPUT58), .A2(n1118), .ZN(n1244) );
AND4_X1 U926 ( .A1(n1211), .A2(n1043), .A3(n1054), .A4(n1202), .ZN(n1118) );
INV_X1 U927 ( .A(n1186), .ZN(n1211) );
NAND2_X1 U928 ( .A1(n1245), .A2(n1246), .ZN(n1186) );
XNOR2_X1 U929 ( .A(G116), .B(n1196), .ZN(G18) );
NAND4_X1 U930 ( .A1(n1226), .A2(n1054), .A3(n1197), .A4(n1202), .ZN(n1196) );
NOR2_X1 U931 ( .A1(n1242), .A2(n1247), .ZN(n1197) );
XOR2_X1 U932 ( .A(n1248), .B(G113), .Z(G15) );
NAND2_X1 U933 ( .A1(KEYINPUT35), .A2(n1199), .ZN(n1248) );
NAND4_X1 U934 ( .A1(n1226), .A2(n1200), .A3(n1054), .A4(n1202), .ZN(n1199) );
AND2_X1 U935 ( .A1(n1235), .A2(n1240), .ZN(n1202) );
NOR2_X1 U936 ( .A1(n1249), .A2(n1052), .ZN(n1054) );
INV_X1 U937 ( .A(n1041), .ZN(n1200) );
NAND2_X1 U938 ( .A1(n1247), .A2(n1242), .ZN(n1041) );
INV_X1 U939 ( .A(n1057), .ZN(n1226) );
NAND2_X1 U940 ( .A1(n1243), .A2(n1246), .ZN(n1057) );
XNOR2_X1 U941 ( .A(KEYINPUT20), .B(n1047), .ZN(n1246) );
XOR2_X1 U942 ( .A(n1245), .B(KEYINPUT6), .Z(n1243) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1251), .ZN(G12) );
NAND2_X1 U944 ( .A1(KEYINPUT48), .A2(n1252), .ZN(n1251) );
XOR2_X1 U945 ( .A(n1253), .B(n1254), .Z(n1250) );
NAND2_X1 U946 ( .A1(n1255), .A2(n1235), .ZN(n1254) );
INV_X1 U947 ( .A(n1030), .ZN(n1235) );
NAND2_X1 U948 ( .A1(n1028), .A2(n1025), .ZN(n1030) );
NAND3_X1 U949 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1025) );
NAND2_X1 U950 ( .A1(G210), .A2(G902), .ZN(n1258) );
NAND3_X1 U951 ( .A1(n1259), .A2(n1158), .A3(n1260), .ZN(n1257) );
OR2_X1 U952 ( .A1(n1260), .A2(n1259), .ZN(n1256) );
XOR2_X1 U953 ( .A(n1173), .B(n1261), .Z(n1259) );
NOR2_X1 U954 ( .A1(KEYINPUT52), .A2(n1218), .ZN(n1261) );
NAND2_X1 U955 ( .A1(G224), .A2(n1033), .ZN(n1218) );
XOR2_X1 U956 ( .A(n1111), .B(n1262), .Z(n1173) );
XOR2_X1 U957 ( .A(G125), .B(n1092), .Z(n1262) );
XNOR2_X1 U958 ( .A(n1263), .B(n1264), .ZN(n1111) );
XOR2_X1 U959 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1266) );
NOR2_X1 U961 ( .A1(G113), .A2(KEYINPUT11), .ZN(n1267) );
XOR2_X1 U962 ( .A(n1269), .B(n1270), .Z(n1263) );
XNOR2_X1 U963 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U964 ( .A1(G116), .A2(KEYINPUT61), .ZN(n1272) );
INV_X1 U965 ( .A(G101), .ZN(n1271) );
XNOR2_X1 U966 ( .A(G122), .B(KEYINPUT60), .ZN(n1269) );
NAND2_X1 U967 ( .A1(G210), .A2(G237), .ZN(n1260) );
NAND2_X1 U968 ( .A1(G214), .A2(n1273), .ZN(n1028) );
NAND2_X1 U969 ( .A1(n1274), .A2(n1158), .ZN(n1273) );
XOR2_X1 U970 ( .A(n1203), .B(KEYINPUT37), .Z(n1255) );
NAND4_X1 U971 ( .A1(n1043), .A2(n1188), .A3(n1201), .A4(n1240), .ZN(n1203) );
NAND2_X1 U972 ( .A1(n1031), .A2(n1275), .ZN(n1240) );
NAND4_X1 U973 ( .A1(G953), .A2(G902), .A3(n1237), .A4(n1107), .ZN(n1275) );
INV_X1 U974 ( .A(G898), .ZN(n1107) );
NAND3_X1 U975 ( .A1(n1237), .A2(n1033), .A3(G952), .ZN(n1031) );
NAND2_X1 U976 ( .A1(G237), .A2(G234), .ZN(n1237) );
NOR2_X1 U977 ( .A1(n1053), .A2(n1052), .ZN(n1201) );
AND2_X1 U978 ( .A1(G221), .A2(n1276), .ZN(n1052) );
INV_X1 U979 ( .A(n1249), .ZN(n1053) );
XNOR2_X1 U980 ( .A(n1277), .B(G469), .ZN(n1249) );
NAND2_X1 U981 ( .A1(n1278), .A2(n1158), .ZN(n1277) );
XOR2_X1 U982 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U983 ( .A(n1143), .B(n1281), .Z(n1280) );
XNOR2_X1 U984 ( .A(KEYINPUT18), .B(n1282), .ZN(n1281) );
INV_X1 U985 ( .A(G140), .ZN(n1282) );
XNOR2_X1 U986 ( .A(n1153), .B(n1163), .ZN(n1279) );
XOR2_X1 U987 ( .A(G101), .B(n1283), .Z(n1163) );
NOR2_X1 U988 ( .A1(KEYINPUT12), .A2(n1265), .ZN(n1283) );
XNOR2_X1 U989 ( .A(n1284), .B(n1285), .ZN(n1265) );
XNOR2_X1 U990 ( .A(G107), .B(KEYINPUT26), .ZN(n1284) );
XOR2_X1 U991 ( .A(G110), .B(n1286), .Z(n1153) );
NOR2_X1 U992 ( .A1(G953), .A2(n1078), .ZN(n1286) );
INV_X1 U993 ( .A(G227), .ZN(n1078) );
INV_X1 U994 ( .A(n1056), .ZN(n1188) );
NAND2_X1 U995 ( .A1(n1047), .A2(n1245), .ZN(n1056) );
XOR2_X1 U996 ( .A(n1068), .B(n1287), .Z(n1245) );
NOR2_X1 U997 ( .A1(n1070), .A2(KEYINPUT10), .ZN(n1287) );
INV_X1 U998 ( .A(n1123), .ZN(n1070) );
NAND2_X1 U999 ( .A1(G217), .A2(n1276), .ZN(n1123) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1158), .ZN(n1276) );
NAND2_X1 U1001 ( .A1(n1288), .A2(n1121), .ZN(n1068) );
XNOR2_X1 U1002 ( .A(n1289), .B(n1290), .ZN(n1121) );
XOR2_X1 U1003 ( .A(n1291), .B(n1268), .Z(n1290) );
XNOR2_X1 U1004 ( .A(n1292), .B(G119), .ZN(n1268) );
INV_X1 U1005 ( .A(G110), .ZN(n1292) );
XNOR2_X1 U1006 ( .A(n1293), .B(n1101), .ZN(n1289) );
XOR2_X1 U1007 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U1009 ( .A(KEYINPUT29), .B(n1158), .ZN(n1288) );
XNOR2_X1 U1010 ( .A(n1066), .B(n1067), .ZN(n1047) );
INV_X1 U1011 ( .A(G472), .ZN(n1067) );
NAND2_X1 U1012 ( .A1(n1297), .A2(n1158), .ZN(n1066) );
INV_X1 U1013 ( .A(G902), .ZN(n1158) );
XOR2_X1 U1014 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U1015 ( .A(n1144), .B(n1147), .Z(n1299) );
XNOR2_X1 U1016 ( .A(G101), .B(n1300), .ZN(n1147) );
NOR3_X1 U1017 ( .A1(n1174), .A2(G953), .A3(G237), .ZN(n1300) );
INV_X1 U1018 ( .A(G210), .ZN(n1174) );
XNOR2_X1 U1019 ( .A(n1301), .B(n1302), .ZN(n1144) );
NOR2_X1 U1020 ( .A1(G113), .A2(KEYINPUT50), .ZN(n1302) );
NAND2_X1 U1021 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U1022 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1023 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND2_X1 U1024 ( .A1(KEYINPUT43), .A2(n1309), .ZN(n1308) );
INV_X1 U1025 ( .A(G119), .ZN(n1309) );
NAND2_X1 U1026 ( .A1(G119), .A2(n1310), .ZN(n1303) );
NAND2_X1 U1027 ( .A1(KEYINPUT43), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1028 ( .A1(G116), .A2(n1307), .ZN(n1311) );
INV_X1 U1029 ( .A(KEYINPUT25), .ZN(n1307) );
XNOR2_X1 U1030 ( .A(KEYINPUT7), .B(n1312), .ZN(n1298) );
NOR2_X1 U1031 ( .A1(KEYINPUT62), .A2(n1143), .ZN(n1312) );
XNOR2_X1 U1032 ( .A(n1168), .B(n1092), .ZN(n1143) );
XOR2_X1 U1033 ( .A(G143), .B(n1295), .Z(n1092) );
XNOR2_X1 U1034 ( .A(G146), .B(n1230), .ZN(n1295) );
INV_X1 U1035 ( .A(G128), .ZN(n1230) );
NAND2_X1 U1036 ( .A1(n1313), .A2(n1314), .ZN(n1168) );
NAND2_X1 U1037 ( .A1(G131), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1038 ( .A(n1316), .B(KEYINPUT59), .Z(n1313) );
OR2_X1 U1039 ( .A1(n1315), .A2(G131), .ZN(n1316) );
XNOR2_X1 U1040 ( .A(G134), .B(n1101), .ZN(n1315) );
INV_X1 U1041 ( .A(n1098), .ZN(n1101) );
XOR2_X1 U1042 ( .A(G137), .B(KEYINPUT39), .Z(n1098) );
NOR2_X1 U1043 ( .A1(n1242), .A2(n1241), .ZN(n1043) );
INV_X1 U1044 ( .A(n1247), .ZN(n1241) );
XNOR2_X1 U1045 ( .A(n1317), .B(n1071), .ZN(n1247) );
NOR2_X1 U1046 ( .A1(n1128), .A2(G902), .ZN(n1071) );
XNOR2_X1 U1047 ( .A(n1318), .B(n1319), .ZN(n1128) );
XOR2_X1 U1048 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1049 ( .A(n1014), .B(n1322), .ZN(n1321) );
NOR2_X1 U1050 ( .A1(KEYINPUT33), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1051 ( .A(n1324), .B(G122), .Z(n1323) );
NAND2_X1 U1052 ( .A1(KEYINPUT1), .A2(n1306), .ZN(n1324) );
INV_X1 U1053 ( .A(G116), .ZN(n1306) );
INV_X1 U1054 ( .A(G107), .ZN(n1014) );
AND2_X1 U1055 ( .A1(n1296), .A2(G217), .ZN(n1320) );
AND2_X1 U1056 ( .A1(G234), .A2(n1033), .ZN(n1296) );
XNOR2_X1 U1057 ( .A(G128), .B(n1325), .ZN(n1318) );
XNOR2_X1 U1058 ( .A(n1220), .B(G134), .ZN(n1325) );
NAND2_X1 U1059 ( .A1(KEYINPUT32), .A2(n1132), .ZN(n1317) );
INV_X1 U1060 ( .A(G478), .ZN(n1132) );
XNOR2_X1 U1061 ( .A(n1326), .B(n1072), .ZN(n1242) );
NOR2_X1 U1062 ( .A1(n1136), .A2(n1327), .ZN(n1072) );
XNOR2_X1 U1063 ( .A(KEYINPUT44), .B(G902), .ZN(n1327) );
XNOR2_X1 U1064 ( .A(n1328), .B(n1329), .ZN(n1136) );
XOR2_X1 U1065 ( .A(n1093), .B(n1330), .Z(n1329) );
XOR2_X1 U1066 ( .A(n1331), .B(n1285), .Z(n1330) );
XNOR2_X1 U1067 ( .A(n1139), .B(KEYINPUT36), .ZN(n1285) );
INV_X1 U1068 ( .A(G104), .ZN(n1139) );
NOR2_X1 U1069 ( .A1(G113), .A2(KEYINPUT13), .ZN(n1331) );
XOR2_X1 U1070 ( .A(G131), .B(n1291), .Z(n1093) );
XOR2_X1 U1071 ( .A(G125), .B(G140), .Z(n1291) );
XOR2_X1 U1072 ( .A(n1332), .B(n1333), .Z(n1328) );
XOR2_X1 U1073 ( .A(G146), .B(G122), .Z(n1333) );
NAND2_X1 U1074 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
NAND4_X1 U1075 ( .A1(G214), .A2(G143), .A3(n1274), .A4(n1033), .ZN(n1335) );
XOR2_X1 U1076 ( .A(n1336), .B(KEYINPUT49), .Z(n1334) );
NAND2_X1 U1077 ( .A1(n1220), .A2(n1337), .ZN(n1336) );
NAND3_X1 U1078 ( .A1(n1274), .A2(n1033), .A3(G214), .ZN(n1337) );
INV_X1 U1079 ( .A(G953), .ZN(n1033) );
INV_X1 U1080 ( .A(G237), .ZN(n1274) );
INV_X1 U1081 ( .A(G143), .ZN(n1220) );
NAND2_X1 U1082 ( .A1(KEYINPUT4), .A2(n1073), .ZN(n1326) );
XOR2_X1 U1083 ( .A(G475), .B(KEYINPUT24), .Z(n1073) );
OR2_X1 U1084 ( .A1(n1252), .A2(KEYINPUT48), .ZN(n1253) );
XOR2_X1 U1085 ( .A(G110), .B(KEYINPUT57), .Z(n1252) );
endmodule


