//Key = 0000011111101010010111100011110010010111111000110101100000010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371;

XNOR2_X1 U760 ( .A(G107), .B(n1040), .ZN(G9) );
NOR2_X1 U761 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
XOR2_X1 U763 ( .A(n1047), .B(KEYINPUT31), .Z(n1046) );
NAND2_X1 U764 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U765 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND2_X1 U766 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND3_X1 U767 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND3_X1 U769 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U770 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND4_X1 U771 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1061) );
INV_X1 U772 ( .A(KEYINPUT18), .ZN(n1068) );
NAND2_X1 U773 ( .A1(KEYINPUT18), .A2(n1055), .ZN(n1060) );
NAND2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1048) );
INV_X1 U775 ( .A(n1071), .ZN(n1069) );
NOR2_X1 U776 ( .A1(n1072), .A2(n1071), .ZN(n1045) );
NAND3_X1 U777 ( .A1(n1055), .A2(n1058), .A3(n1052), .ZN(n1071) );
NAND3_X1 U778 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1043) );
NAND3_X1 U779 ( .A1(n1050), .A2(n1076), .A3(n1052), .ZN(n1075) );
INV_X1 U780 ( .A(n1077), .ZN(n1052) );
NAND3_X1 U781 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1076) );
NAND2_X1 U782 ( .A1(n1055), .A2(n1081), .ZN(n1080) );
AND2_X1 U783 ( .A1(n1063), .A2(n1066), .ZN(n1055) );
NAND3_X1 U784 ( .A1(n1082), .A2(n1058), .A3(n1063), .ZN(n1079) );
NAND2_X1 U785 ( .A1(n1083), .A2(n1066), .ZN(n1078) );
NOR3_X1 U786 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1041) );
INV_X1 U787 ( .A(n1073), .ZN(n1084) );
NAND4_X1 U788 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1073) );
NOR4_X1 U789 ( .A1(n1057), .A2(n1067), .A3(n1089), .A4(n1090), .ZN(n1088) );
XNOR2_X1 U790 ( .A(n1091), .B(n1092), .ZN(n1089) );
NAND2_X1 U791 ( .A1(n1093), .A2(KEYINPUT8), .ZN(n1091) );
XOR2_X1 U792 ( .A(n1094), .B(KEYINPUT58), .Z(n1093) );
INV_X1 U793 ( .A(n1095), .ZN(n1067) );
NOR2_X1 U794 ( .A1(n1096), .A2(n1097), .ZN(n1087) );
XOR2_X1 U795 ( .A(n1098), .B(n1099), .Z(n1086) );
NAND2_X1 U796 ( .A1(KEYINPUT47), .A2(G475), .ZN(n1098) );
XOR2_X1 U797 ( .A(n1100), .B(n1101), .Z(n1085) );
NOR2_X1 U798 ( .A1(KEYINPUT61), .A2(n1102), .ZN(n1101) );
XOR2_X1 U799 ( .A(n1103), .B(n1104), .Z(G72) );
NOR2_X1 U800 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U801 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U802 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U803 ( .A(G140), .B(n1111), .ZN(n1107) );
NAND3_X1 U804 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1103) );
INV_X1 U805 ( .A(n1105), .ZN(n1114) );
OR2_X1 U806 ( .A1(n1074), .A2(G227), .ZN(n1113) );
NAND2_X1 U807 ( .A1(n1115), .A2(n1074), .ZN(n1112) );
NAND2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U809 ( .A(n1118), .B(KEYINPUT24), .Z(n1116) );
XOR2_X1 U810 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U811 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR3_X1 U812 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
INV_X1 U813 ( .A(n1126), .ZN(n1124) );
NOR2_X1 U814 ( .A1(G898), .A2(n1074), .ZN(n1123) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1074), .ZN(n1121) );
NAND2_X1 U816 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U817 ( .A(KEYINPUT52), .B(n1130), .ZN(n1129) );
NAND2_X1 U818 ( .A1(G953), .A2(n1131), .ZN(n1119) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1131) );
NOR2_X1 U820 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U821 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR3_X1 U822 ( .A1(n1136), .A2(KEYINPUT13), .A3(n1137), .ZN(n1135) );
NOR2_X1 U823 ( .A1(n1132), .A2(n1138), .ZN(G63) );
XOR2_X1 U824 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U825 ( .A1(n1102), .A2(n1136), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1132), .A2(n1141), .ZN(G60) );
XOR2_X1 U827 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U828 ( .A(KEYINPUT35), .B(n1144), .Z(n1143) );
AND2_X1 U829 ( .A1(G475), .A2(n1145), .ZN(n1142) );
NAND3_X1 U830 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(G6) );
OR2_X1 U831 ( .A1(n1130), .A2(G104), .ZN(n1148) );
NAND2_X1 U832 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
INV_X1 U833 ( .A(KEYINPUT17), .ZN(n1150) );
NAND2_X1 U834 ( .A1(G104), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U835 ( .A(KEYINPUT7), .B(n1130), .ZN(n1151) );
NAND2_X1 U836 ( .A1(KEYINPUT17), .A2(n1152), .ZN(n1146) );
NAND2_X1 U837 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND3_X1 U838 ( .A1(KEYINPUT7), .A2(G104), .A3(n1130), .ZN(n1154) );
OR2_X1 U839 ( .A1(n1130), .A2(KEYINPUT7), .ZN(n1153) );
NOR2_X1 U840 ( .A1(n1132), .A2(n1155), .ZN(G57) );
XOR2_X1 U841 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U842 ( .A1(n1158), .A2(KEYINPUT56), .ZN(n1157) );
XOR2_X1 U843 ( .A(n1159), .B(G101), .Z(n1156) );
NAND3_X1 U844 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1159) );
OR2_X1 U845 ( .A1(n1163), .A2(KEYINPUT14), .ZN(n1162) );
NAND4_X1 U846 ( .A1(n1163), .A2(KEYINPUT51), .A3(KEYINPUT14), .A4(n1164), .ZN(n1161) );
AND2_X1 U847 ( .A1(n1145), .A2(G472), .ZN(n1163) );
NAND2_X1 U848 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND3_X1 U849 ( .A1(n1145), .A2(G472), .A3(KEYINPUT51), .ZN(n1166) );
INV_X1 U850 ( .A(n1164), .ZN(n1165) );
XOR2_X1 U851 ( .A(n1167), .B(n1168), .Z(n1164) );
NOR2_X1 U852 ( .A1(n1132), .A2(n1169), .ZN(G54) );
XNOR2_X1 U853 ( .A(n1170), .B(n1171), .ZN(n1169) );
XOR2_X1 U854 ( .A(n1172), .B(n1173), .Z(n1171) );
AND2_X1 U855 ( .A1(G469), .A2(n1145), .ZN(n1173) );
INV_X1 U856 ( .A(n1136), .ZN(n1145) );
NAND3_X1 U857 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1172) );
OR2_X1 U858 ( .A1(n1177), .A2(KEYINPUT29), .ZN(n1175) );
NAND3_X1 U859 ( .A1(n1177), .A2(n1178), .A3(KEYINPUT29), .ZN(n1174) );
NOR2_X1 U860 ( .A1(n1132), .A2(n1179), .ZN(G51) );
XOR2_X1 U861 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U862 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR2_X1 U863 ( .A1(KEYINPUT43), .A2(n1184), .ZN(n1183) );
NOR2_X1 U864 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U865 ( .A(n1187), .B(KEYINPUT39), .Z(n1186) );
NAND2_X1 U866 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U867 ( .A1(n1094), .A2(n1136), .ZN(n1180) );
NAND2_X1 U868 ( .A1(G902), .A2(n1044), .ZN(n1136) );
NAND4_X1 U869 ( .A1(n1128), .A2(n1117), .A3(n1118), .A4(n1130), .ZN(n1044) );
NAND3_X1 U870 ( .A1(n1190), .A2(n1066), .A3(n1191), .ZN(n1130) );
AND2_X1 U871 ( .A1(n1192), .A2(n1193), .ZN(n1117) );
AND4_X1 U872 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR4_X1 U873 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1192) );
NOR3_X1 U874 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1201) );
XNOR2_X1 U875 ( .A(KEYINPUT42), .B(n1205), .ZN(n1202) );
INV_X1 U876 ( .A(n1206), .ZN(n1200) );
NOR2_X1 U877 ( .A1(n1207), .A2(n1208), .ZN(n1199) );
INV_X1 U878 ( .A(KEYINPUT59), .ZN(n1207) );
NOR3_X1 U879 ( .A1(KEYINPUT59), .A2(n1191), .A3(n1209), .ZN(n1198) );
AND2_X1 U880 ( .A1(n1210), .A2(n1211), .ZN(n1128) );
AND4_X1 U881 ( .A1(n1212), .A2(n1213), .A3(n1040), .A4(n1214), .ZN(n1211) );
NAND3_X1 U882 ( .A1(n1190), .A2(n1066), .A3(n1070), .ZN(n1040) );
NOR4_X1 U883 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1210) );
NOR2_X1 U884 ( .A1(KEYINPUT57), .A2(n1219), .ZN(n1218) );
NOR2_X1 U885 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
NOR2_X1 U886 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
AND3_X1 U887 ( .A1(n1082), .A2(n1224), .A3(n1190), .ZN(n1223) );
NOR4_X1 U888 ( .A1(n1205), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1222) );
INV_X1 U889 ( .A(KEYINPUT57), .ZN(n1227) );
NAND2_X1 U890 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
NOR3_X1 U891 ( .A1(n1224), .A2(n1230), .A3(n1228), .ZN(n1216) );
NOR4_X1 U892 ( .A1(n1231), .A2(n1205), .A3(n1232), .A4(n1221), .ZN(n1230) );
INV_X1 U893 ( .A(KEYINPUT48), .ZN(n1224) );
INV_X1 U894 ( .A(n1233), .ZN(n1215) );
NOR2_X1 U895 ( .A1(n1074), .A2(G952), .ZN(n1132) );
XNOR2_X1 U896 ( .A(G146), .B(n1206), .ZN(G48) );
NAND3_X1 U897 ( .A1(n1191), .A2(n1234), .A3(n1235), .ZN(n1206) );
XNOR2_X1 U898 ( .A(n1197), .B(n1236), .ZN(G45) );
NOR2_X1 U899 ( .A1(KEYINPUT44), .A2(n1237), .ZN(n1236) );
NAND4_X1 U900 ( .A1(n1238), .A2(n1234), .A3(n1239), .A4(n1240), .ZN(n1197) );
XOR2_X1 U901 ( .A(n1196), .B(n1241), .Z(G42) );
XOR2_X1 U902 ( .A(KEYINPUT19), .B(G140), .Z(n1241) );
NAND3_X1 U903 ( .A1(n1063), .A2(n1081), .A3(n1242), .ZN(n1196) );
XNOR2_X1 U904 ( .A(G137), .B(n1243), .ZN(G39) );
NAND2_X1 U905 ( .A1(n1244), .A2(n1235), .ZN(n1243) );
INV_X1 U906 ( .A(n1204), .ZN(n1244) );
NAND2_X1 U907 ( .A1(n1063), .A2(n1050), .ZN(n1204) );
XOR2_X1 U908 ( .A(G134), .B(n1245), .Z(G36) );
NOR2_X1 U909 ( .A1(KEYINPUT34), .A2(n1118), .ZN(n1245) );
NAND2_X1 U910 ( .A1(n1246), .A2(n1070), .ZN(n1118) );
NAND2_X1 U911 ( .A1(n1247), .A2(n1248), .ZN(G33) );
NAND2_X1 U912 ( .A1(KEYINPUT54), .A2(n1249), .ZN(n1248) );
XOR2_X1 U913 ( .A(n1208), .B(n1250), .Z(n1247) );
NOR2_X1 U914 ( .A1(KEYINPUT54), .A2(n1249), .ZN(n1250) );
INV_X1 U915 ( .A(G131), .ZN(n1249) );
NAND2_X1 U916 ( .A1(n1246), .A2(n1191), .ZN(n1208) );
INV_X1 U917 ( .A(n1209), .ZN(n1246) );
NAND2_X1 U918 ( .A1(n1063), .A2(n1238), .ZN(n1209) );
AND3_X1 U919 ( .A1(n1081), .A2(n1251), .A3(n1082), .ZN(n1238) );
AND2_X1 U920 ( .A1(n1065), .A2(n1095), .ZN(n1063) );
XNOR2_X1 U921 ( .A(n1252), .B(KEYINPUT4), .ZN(n1065) );
XNOR2_X1 U922 ( .A(G128), .B(n1195), .ZN(G30) );
NAND3_X1 U923 ( .A1(n1070), .A2(n1234), .A3(n1235), .ZN(n1195) );
NOR2_X1 U924 ( .A1(n1203), .A2(n1205), .ZN(n1235) );
NAND3_X1 U925 ( .A1(n1097), .A2(n1251), .A3(n1096), .ZN(n1203) );
XOR2_X1 U926 ( .A(n1253), .B(n1254), .Z(G3) );
XOR2_X1 U927 ( .A(KEYINPUT37), .B(G101), .Z(n1254) );
NAND3_X1 U928 ( .A1(n1190), .A2(n1255), .A3(n1082), .ZN(n1253) );
XNOR2_X1 U929 ( .A(KEYINPUT2), .B(n1221), .ZN(n1255) );
INV_X1 U930 ( .A(n1050), .ZN(n1221) );
XNOR2_X1 U931 ( .A(G125), .B(n1194), .ZN(G27) );
NAND2_X1 U932 ( .A1(n1242), .A2(n1083), .ZN(n1194) );
AND3_X1 U933 ( .A1(n1191), .A2(n1251), .A3(n1064), .ZN(n1242) );
NAND2_X1 U934 ( .A1(n1077), .A2(n1256), .ZN(n1251) );
NAND3_X1 U935 ( .A1(G902), .A2(n1257), .A3(n1105), .ZN(n1256) );
NOR2_X1 U936 ( .A1(G900), .A2(n1074), .ZN(n1105) );
XNOR2_X1 U937 ( .A(G122), .B(n1233), .ZN(G24) );
NAND4_X1 U938 ( .A1(n1258), .A2(n1066), .A3(n1239), .A4(n1240), .ZN(n1233) );
AND2_X1 U939 ( .A1(n1259), .A2(n1260), .ZN(n1066) );
XNOR2_X1 U940 ( .A(G119), .B(n1213), .ZN(G21) );
NAND4_X1 U941 ( .A1(n1050), .A2(n1258), .A3(n1096), .A4(n1097), .ZN(n1213) );
XNOR2_X1 U942 ( .A(G116), .B(n1212), .ZN(G18) );
NAND3_X1 U943 ( .A1(n1082), .A2(n1070), .A3(n1258), .ZN(n1212) );
NOR2_X1 U944 ( .A1(n1239), .A2(n1261), .ZN(n1070) );
INV_X1 U945 ( .A(n1240), .ZN(n1261) );
XNOR2_X1 U946 ( .A(G113), .B(n1214), .ZN(G15) );
NAND3_X1 U947 ( .A1(n1258), .A2(n1082), .A3(n1191), .ZN(n1214) );
INV_X1 U948 ( .A(n1072), .ZN(n1191) );
NAND2_X1 U949 ( .A1(n1262), .A2(n1239), .ZN(n1072) );
XNOR2_X1 U950 ( .A(n1240), .B(KEYINPUT25), .ZN(n1262) );
INV_X1 U951 ( .A(n1232), .ZN(n1082) );
NAND2_X1 U952 ( .A1(n1260), .A2(n1097), .ZN(n1232) );
INV_X1 U953 ( .A(n1096), .ZN(n1260) );
AND2_X1 U954 ( .A1(n1083), .A2(n1229), .ZN(n1258) );
AND2_X1 U955 ( .A1(n1058), .A2(n1234), .ZN(n1083) );
INV_X1 U956 ( .A(n1228), .ZN(n1234) );
AND2_X1 U957 ( .A1(n1056), .A2(n1263), .ZN(n1058) );
NAND2_X1 U958 ( .A1(n1264), .A2(n1265), .ZN(G12) );
NAND2_X1 U959 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U960 ( .A(KEYINPUT21), .B(n1268), .Z(n1264) );
NOR2_X1 U961 ( .A1(n1266), .A2(n1267), .ZN(n1268) );
INV_X1 U962 ( .A(n1219), .ZN(n1266) );
NAND3_X1 U963 ( .A1(n1050), .A2(n1190), .A3(n1064), .ZN(n1219) );
INV_X1 U964 ( .A(n1226), .ZN(n1064) );
NAND2_X1 U965 ( .A1(n1259), .A2(n1096), .ZN(n1226) );
XNOR2_X1 U966 ( .A(n1137), .B(n1269), .ZN(n1096) );
NOR2_X1 U967 ( .A1(G902), .A2(n1270), .ZN(n1269) );
XOR2_X1 U968 ( .A(n1134), .B(KEYINPUT28), .Z(n1270) );
NAND2_X1 U969 ( .A1(n1271), .A2(n1272), .ZN(n1134) );
NAND2_X1 U970 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U971 ( .A(n1275), .B(KEYINPUT1), .Z(n1271) );
OR2_X1 U972 ( .A1(n1274), .A2(n1273), .ZN(n1275) );
XOR2_X1 U973 ( .A(n1276), .B(n1277), .Z(n1273) );
AND4_X1 U974 ( .A1(n1278), .A2(n1279), .A3(G234), .A4(G221), .ZN(n1277) );
INV_X1 U975 ( .A(KEYINPUT45), .ZN(n1278) );
XNOR2_X1 U976 ( .A(G137), .B(KEYINPUT62), .ZN(n1276) );
XNOR2_X1 U977 ( .A(n1280), .B(n1281), .ZN(n1274) );
XOR2_X1 U978 ( .A(n1282), .B(n1177), .Z(n1281) );
XNOR2_X1 U979 ( .A(G119), .B(n1283), .ZN(n1280) );
XNOR2_X1 U980 ( .A(KEYINPUT16), .B(n1111), .ZN(n1283) );
INV_X1 U981 ( .A(G125), .ZN(n1111) );
NAND2_X1 U982 ( .A1(G217), .A2(n1284), .ZN(n1137) );
XNOR2_X1 U983 ( .A(n1097), .B(KEYINPUT63), .ZN(n1259) );
XNOR2_X1 U984 ( .A(n1285), .B(G472), .ZN(n1097) );
NAND2_X1 U985 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U986 ( .A(n1288), .B(n1289), .Z(n1286) );
XOR2_X1 U987 ( .A(n1290), .B(n1167), .Z(n1289) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1167) );
XNOR2_X1 U989 ( .A(G116), .B(n1293), .ZN(n1292) );
NAND2_X1 U990 ( .A1(n1294), .A2(KEYINPUT10), .ZN(n1293) );
XNOR2_X1 U991 ( .A(G113), .B(KEYINPUT30), .ZN(n1294) );
XNOR2_X1 U992 ( .A(n1109), .B(n1295), .ZN(n1291) );
NOR2_X1 U993 ( .A1(KEYINPUT23), .A2(n1296), .ZN(n1295) );
NAND2_X1 U994 ( .A1(KEYINPUT27), .A2(n1168), .ZN(n1290) );
XNOR2_X1 U995 ( .A(n1158), .B(n1297), .ZN(n1288) );
XNOR2_X1 U996 ( .A(G101), .B(KEYINPUT53), .ZN(n1297) );
AND2_X1 U997 ( .A1(G210), .A2(n1298), .ZN(n1158) );
NOR3_X1 U998 ( .A1(n1228), .A2(n1231), .A3(n1205), .ZN(n1190) );
INV_X1 U999 ( .A(n1081), .ZN(n1205) );
NOR2_X1 U1000 ( .A1(n1056), .A2(n1057), .ZN(n1081) );
INV_X1 U1001 ( .A(n1263), .ZN(n1057) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1284), .ZN(n1263) );
NAND2_X1 U1003 ( .A1(G234), .A2(n1287), .ZN(n1284) );
XOR2_X1 U1004 ( .A(n1090), .B(KEYINPUT6), .Z(n1056) );
XNOR2_X1 U1005 ( .A(n1299), .B(G469), .ZN(n1090) );
NAND2_X1 U1006 ( .A1(n1300), .A2(n1287), .ZN(n1299) );
XOR2_X1 U1007 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U1008 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND3_X1 U1009 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
INV_X1 U1010 ( .A(KEYINPUT22), .ZN(n1307) );
NAND2_X1 U1011 ( .A1(n1170), .A2(KEYINPUT22), .ZN(n1303) );
XOR2_X1 U1012 ( .A(n1306), .B(n1305), .Z(n1170) );
XNOR2_X1 U1013 ( .A(n1308), .B(n1309), .ZN(n1305) );
XOR2_X1 U1014 ( .A(n1310), .B(n1110), .Z(n1309) );
XNOR2_X1 U1015 ( .A(n1311), .B(n1312), .ZN(n1110) );
XNOR2_X1 U1016 ( .A(n1313), .B(n1314), .ZN(n1312) );
NOR2_X1 U1017 ( .A1(G143), .A2(KEYINPUT60), .ZN(n1314) );
NAND2_X1 U1018 ( .A1(KEYINPUT20), .A2(n1315), .ZN(n1311) );
XNOR2_X1 U1019 ( .A(KEYINPUT33), .B(n1316), .ZN(n1308) );
NOR2_X1 U1020 ( .A1(G104), .A2(KEYINPUT36), .ZN(n1316) );
XOR2_X1 U1021 ( .A(n1109), .B(KEYINPUT40), .Z(n1306) );
XOR2_X1 U1022 ( .A(G131), .B(n1317), .Z(n1109) );
XOR2_X1 U1023 ( .A(G137), .B(G134), .Z(n1317) );
NAND2_X1 U1024 ( .A1(n1176), .A2(n1318), .ZN(n1301) );
NAND2_X1 U1025 ( .A1(n1177), .A2(n1178), .ZN(n1318) );
OR2_X1 U1026 ( .A1(n1178), .A2(n1177), .ZN(n1176) );
XNOR2_X1 U1027 ( .A(n1267), .B(G140), .ZN(n1177) );
NAND2_X1 U1028 ( .A1(G227), .A2(n1279), .ZN(n1178) );
INV_X1 U1029 ( .A(n1229), .ZN(n1231) );
NAND2_X1 U1030 ( .A1(n1077), .A2(n1319), .ZN(n1229) );
NAND4_X1 U1031 ( .A1(G902), .A2(G953), .A3(n1257), .A4(n1320), .ZN(n1319) );
INV_X1 U1032 ( .A(G898), .ZN(n1320) );
NAND3_X1 U1033 ( .A1(n1257), .A2(n1074), .A3(G952), .ZN(n1077) );
INV_X1 U1034 ( .A(G953), .ZN(n1074) );
NAND2_X1 U1035 ( .A1(G237), .A2(G234), .ZN(n1257) );
NAND2_X1 U1036 ( .A1(n1252), .A2(n1095), .ZN(n1228) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1321), .ZN(n1095) );
XOR2_X1 U1038 ( .A(n1092), .B(n1094), .Z(n1252) );
NAND2_X1 U1039 ( .A1(G210), .A2(n1321), .ZN(n1094) );
NAND2_X1 U1040 ( .A1(n1322), .A2(n1287), .ZN(n1321) );
NAND2_X1 U1041 ( .A1(n1323), .A2(n1287), .ZN(n1092) );
XOR2_X1 U1042 ( .A(n1182), .B(n1324), .Z(n1323) );
NAND2_X1 U1043 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1044 ( .A1(n1327), .A2(n1188), .ZN(n1326) );
XNOR2_X1 U1045 ( .A(KEYINPUT41), .B(n1189), .ZN(n1327) );
INV_X1 U1046 ( .A(n1185), .ZN(n1325) );
NOR2_X1 U1047 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
NAND2_X1 U1048 ( .A1(G224), .A2(n1279), .ZN(n1189) );
XNOR2_X1 U1049 ( .A(n1168), .B(G125), .ZN(n1188) );
XNOR2_X1 U1050 ( .A(G143), .B(n1282), .ZN(n1168) );
XNOR2_X1 U1051 ( .A(n1315), .B(G146), .ZN(n1282) );
INV_X1 U1052 ( .A(G128), .ZN(n1315) );
NAND2_X1 U1053 ( .A1(n1328), .A2(n1126), .ZN(n1182) );
NAND2_X1 U1054 ( .A1(n1329), .A2(n1330), .ZN(n1126) );
XOR2_X1 U1055 ( .A(KEYINPUT9), .B(n1125), .Z(n1328) );
NOR2_X1 U1056 ( .A1(n1330), .A2(n1329), .ZN(n1125) );
XOR2_X1 U1057 ( .A(n1331), .B(n1332), .Z(n1329) );
XNOR2_X1 U1058 ( .A(n1296), .B(n1333), .ZN(n1332) );
XOR2_X1 U1059 ( .A(KEYINPUT55), .B(KEYINPUT30), .Z(n1333) );
INV_X1 U1060 ( .A(G119), .ZN(n1296) );
XOR2_X1 U1061 ( .A(n1334), .B(n1310), .Z(n1331) );
XOR2_X1 U1062 ( .A(G107), .B(G101), .Z(n1310) );
XNOR2_X1 U1063 ( .A(G116), .B(n1335), .ZN(n1334) );
NAND2_X1 U1064 ( .A1(n1336), .A2(n1337), .ZN(n1330) );
NAND2_X1 U1065 ( .A1(G122), .A2(n1267), .ZN(n1337) );
XOR2_X1 U1066 ( .A(KEYINPUT46), .B(n1338), .Z(n1336) );
NOR2_X1 U1067 ( .A1(G122), .A2(n1267), .ZN(n1338) );
INV_X1 U1068 ( .A(G110), .ZN(n1267) );
NOR2_X1 U1069 ( .A1(n1240), .A2(n1239), .ZN(n1050) );
XOR2_X1 U1070 ( .A(G475), .B(n1099), .Z(n1239) );
AND2_X1 U1071 ( .A1(n1144), .A2(n1339), .ZN(n1099) );
XNOR2_X1 U1072 ( .A(KEYINPUT38), .B(n1287), .ZN(n1339) );
INV_X1 U1073 ( .A(G902), .ZN(n1287) );
AND3_X1 U1074 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1144) );
NAND2_X1 U1075 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND2_X1 U1076 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XNOR2_X1 U1077 ( .A(n1347), .B(n1335), .ZN(n1343) );
NAND4_X1 U1078 ( .A1(n1345), .A2(n1346), .A3(n1348), .A4(n1349), .ZN(n1341) );
XNOR2_X1 U1079 ( .A(G122), .B(n1335), .ZN(n1348) );
XOR2_X1 U1080 ( .A(G113), .B(G104), .Z(n1335) );
INV_X1 U1081 ( .A(KEYINPUT11), .ZN(n1346) );
OR2_X1 U1082 ( .A1(n1345), .A2(n1349), .ZN(n1340) );
INV_X1 U1083 ( .A(KEYINPUT3), .ZN(n1349) );
XOR2_X1 U1084 ( .A(n1350), .B(n1351), .Z(n1345) );
XNOR2_X1 U1085 ( .A(n1237), .B(G131), .ZN(n1351) );
XOR2_X1 U1086 ( .A(n1352), .B(n1353), .Z(n1350) );
AND2_X1 U1087 ( .A1(n1298), .A2(G214), .ZN(n1353) );
AND2_X1 U1088 ( .A1(n1279), .A2(n1322), .ZN(n1298) );
INV_X1 U1089 ( .A(G237), .ZN(n1322) );
NAND2_X1 U1090 ( .A1(n1354), .A2(n1355), .ZN(n1352) );
NAND2_X1 U1091 ( .A1(n1356), .A2(n1313), .ZN(n1355) );
XOR2_X1 U1092 ( .A(KEYINPUT5), .B(n1357), .Z(n1354) );
NOR2_X1 U1093 ( .A1(n1313), .A2(n1356), .ZN(n1357) );
XNOR2_X1 U1094 ( .A(G125), .B(n1358), .ZN(n1356) );
NAND2_X1 U1095 ( .A1(KEYINPUT12), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1096 ( .A(KEYINPUT32), .B(G140), .Z(n1359) );
INV_X1 U1097 ( .A(G146), .ZN(n1313) );
XOR2_X1 U1098 ( .A(n1100), .B(n1102), .Z(n1240) );
INV_X1 U1099 ( .A(G478), .ZN(n1102) );
OR2_X1 U1100 ( .A1(n1140), .A2(G902), .ZN(n1100) );
XNOR2_X1 U1101 ( .A(n1360), .B(n1361), .ZN(n1140) );
NOR2_X1 U1102 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
XOR2_X1 U1103 ( .A(KEYINPUT15), .B(n1364), .Z(n1363) );
AND2_X1 U1104 ( .A1(n1365), .A2(G134), .ZN(n1364) );
NOR2_X1 U1105 ( .A1(G134), .A2(n1365), .ZN(n1362) );
XNOR2_X1 U1106 ( .A(G128), .B(n1237), .ZN(n1365) );
INV_X1 U1107 ( .A(G143), .ZN(n1237) );
XOR2_X1 U1108 ( .A(n1366), .B(n1367), .Z(n1360) );
NOR2_X1 U1109 ( .A1(KEYINPUT0), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1110 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1111 ( .A(n1347), .B(G116), .ZN(n1370) );
INV_X1 U1112 ( .A(G122), .ZN(n1347) );
NAND2_X1 U1113 ( .A1(KEYINPUT26), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1114 ( .A(KEYINPUT49), .B(G107), .Z(n1371) );
NAND3_X1 U1115 ( .A1(n1279), .A2(G217), .A3(G234), .ZN(n1366) );
XNOR2_X1 U1116 ( .A(G953), .B(KEYINPUT50), .ZN(n1279) );
endmodule


