//Key = 1000110110000110111001100011100001111001001111011001000000111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;

XNOR2_X1 U732 ( .A(G107), .B(n1026), .ZN(G9) );
NAND3_X1 U733 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
XNOR2_X1 U734 ( .A(n1030), .B(KEYINPUT32), .ZN(n1029) );
NAND4_X1 U735 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(G75) );
INV_X1 U736 ( .A(n1035), .ZN(n1034) );
NAND4_X1 U737 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1033) );
NOR4_X1 U738 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
XOR2_X1 U739 ( .A(n1044), .B(n1045), .Z(n1041) );
NOR2_X1 U740 ( .A1(n1046), .A2(KEYINPUT20), .ZN(n1045) );
XOR2_X1 U741 ( .A(n1047), .B(KEYINPUT5), .Z(n1038) );
NAND2_X1 U742 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U743 ( .A(KEYINPUT28), .B(n1050), .ZN(n1048) );
XOR2_X1 U744 ( .A(n1051), .B(KEYINPUT9), .Z(n1036) );
NAND2_X1 U745 ( .A1(G952), .A2(n1052), .ZN(n1032) );
NAND3_X1 U746 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U747 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NAND2_X1 U748 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND3_X1 U749 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U750 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND2_X1 U751 ( .A1(n1037), .A2(n1065), .ZN(n1064) );
OR2_X1 U752 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U753 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
NAND2_X1 U754 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U755 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U756 ( .A1(n1037), .A2(n1074), .A3(n1068), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1077), .ZN(n1076) );
OR2_X1 U759 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U760 ( .A(n1080), .ZN(n1062) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1081), .ZN(n1075) );
NAND2_X1 U762 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U763 ( .A1(n1040), .A2(n1084), .ZN(n1083) );
INV_X1 U764 ( .A(n1085), .ZN(n1056) );
NAND2_X1 U765 ( .A1(KEYINPUT2), .A2(n1086), .ZN(n1053) );
OR2_X1 U766 ( .A1(n1086), .A2(KEYINPUT2), .ZN(n1031) );
XOR2_X1 U767 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U768 ( .A1(n1089), .A2(n1086), .ZN(n1088) );
NOR2_X1 U769 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U770 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
NAND2_X1 U771 ( .A1(n1094), .A2(n1086), .ZN(n1093) );
XOR2_X1 U772 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U773 ( .A1(G900), .A2(n1096), .A3(G953), .ZN(n1092) );
XNOR2_X1 U774 ( .A(n1097), .B(n1098), .ZN(n1096) );
XOR2_X1 U775 ( .A(G131), .B(n1099), .Z(n1098) );
XOR2_X1 U776 ( .A(G137), .B(G134), .Z(n1099) );
XNOR2_X1 U777 ( .A(n1100), .B(n1101), .ZN(n1097) );
NAND2_X1 U778 ( .A1(KEYINPUT17), .A2(n1102), .ZN(n1100) );
NAND2_X1 U779 ( .A1(n1103), .A2(n1104), .ZN(G69) );
NAND2_X1 U780 ( .A1(n1105), .A2(G953), .ZN(n1104) );
XOR2_X1 U781 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U782 ( .A1(G898), .A2(G224), .ZN(n1106) );
NAND2_X1 U783 ( .A1(n1108), .A2(n1086), .ZN(n1103) );
NAND2_X1 U784 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U785 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U786 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
OR3_X1 U787 ( .A1(n1115), .A2(KEYINPUT56), .A3(KEYINPUT12), .ZN(n1114) );
INV_X1 U788 ( .A(n1116), .ZN(n1115) );
NAND2_X1 U789 ( .A1(n1107), .A2(KEYINPUT12), .ZN(n1113) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1117), .ZN(n1109) );
INV_X1 U791 ( .A(n1112), .ZN(n1117) );
NOR2_X1 U792 ( .A1(n1116), .A2(KEYINPUT56), .ZN(n1107) );
NAND3_X1 U793 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1116) );
XOR2_X1 U794 ( .A(KEYINPUT45), .B(n1121), .Z(n1120) );
NOR2_X1 U795 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U796 ( .A1(n1123), .A2(n1122), .ZN(n1119) );
NAND2_X1 U797 ( .A1(G953), .A2(n1124), .ZN(n1118) );
NOR2_X1 U798 ( .A1(n1035), .A2(n1125), .ZN(G66) );
XNOR2_X1 U799 ( .A(n1126), .B(n1127), .ZN(n1125) );
XNOR2_X1 U800 ( .A(KEYINPUT46), .B(n1128), .ZN(n1127) );
AND3_X1 U801 ( .A1(n1129), .A2(n1130), .A3(G217), .ZN(n1128) );
INV_X1 U802 ( .A(KEYINPUT52), .ZN(n1130) );
NOR2_X1 U803 ( .A1(n1035), .A2(n1131), .ZN(G63) );
XOR2_X1 U804 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U805 ( .A1(KEYINPUT1), .A2(n1134), .ZN(n1133) );
XOR2_X1 U806 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U807 ( .A1(n1129), .A2(G478), .ZN(n1132) );
NOR2_X1 U808 ( .A1(n1035), .A2(n1137), .ZN(G60) );
NOR2_X1 U809 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U810 ( .A(KEYINPUT30), .B(n1140), .Z(n1139) );
NOR2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
AND2_X1 U812 ( .A1(n1142), .A2(n1141), .ZN(n1138) );
NAND2_X1 U813 ( .A1(n1129), .A2(G475), .ZN(n1142) );
XNOR2_X1 U814 ( .A(G104), .B(n1143), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1035), .A2(n1144), .ZN(G57) );
XNOR2_X1 U816 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U818 ( .A(n1149), .B(KEYINPUT27), .Z(n1148) );
NAND3_X1 U819 ( .A1(n1129), .A2(G472), .A3(n1150), .ZN(n1149) );
NOR2_X1 U820 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
XNOR2_X1 U821 ( .A(n1152), .B(n1153), .ZN(n1150) );
XNOR2_X1 U822 ( .A(n1154), .B(n1155), .ZN(n1153) );
NAND2_X1 U823 ( .A1(KEYINPUT0), .A2(n1156), .ZN(n1154) );
AND2_X1 U824 ( .A1(G472), .A2(n1129), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1035), .A2(n1157), .ZN(G54) );
XOR2_X1 U826 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U827 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U828 ( .A1(n1162), .A2(KEYINPUT63), .ZN(n1160) );
XNOR2_X1 U829 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR2_X1 U830 ( .A1(G140), .A2(KEYINPUT37), .ZN(n1164) );
XOR2_X1 U831 ( .A(n1165), .B(KEYINPUT57), .Z(n1158) );
NAND2_X1 U832 ( .A1(n1129), .A2(G469), .ZN(n1165) );
NOR2_X1 U833 ( .A1(n1035), .A2(n1166), .ZN(G51) );
XOR2_X1 U834 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U835 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U836 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U837 ( .A1(KEYINPUT26), .A2(n1173), .ZN(n1171) );
XOR2_X1 U838 ( .A(n1174), .B(n1175), .Z(n1167) );
XNOR2_X1 U839 ( .A(KEYINPUT54), .B(KEYINPUT40), .ZN(n1175) );
NAND2_X1 U840 ( .A1(n1129), .A2(n1176), .ZN(n1174) );
XOR2_X1 U841 ( .A(KEYINPUT41), .B(G210), .Z(n1176) );
NOR2_X1 U842 ( .A1(n1177), .A2(n1055), .ZN(n1129) );
NOR2_X1 U843 ( .A1(n1112), .A2(n1095), .ZN(n1055) );
NAND4_X1 U844 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1095) );
AND3_X1 U845 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
NAND2_X1 U846 ( .A1(n1027), .A2(n1185), .ZN(n1180) );
NAND3_X1 U847 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
XNOR2_X1 U848 ( .A(n1189), .B(KEYINPUT10), .ZN(n1188) );
NAND4_X1 U849 ( .A1(n1190), .A2(n1067), .A3(n1191), .A4(n1192), .ZN(n1186) );
OR2_X1 U850 ( .A1(n1193), .A2(KEYINPUT11), .ZN(n1192) );
NAND2_X1 U851 ( .A1(KEYINPUT11), .A2(n1194), .ZN(n1191) );
NAND2_X1 U852 ( .A1(n1195), .A2(n1070), .ZN(n1194) );
NAND3_X1 U853 ( .A1(n1066), .A2(n1078), .A3(n1196), .ZN(n1178) );
NAND3_X1 U854 ( .A1(n1197), .A2(n1143), .A3(n1198), .ZN(n1112) );
NOR3_X1 U855 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
NAND4_X1 U856 ( .A1(n1066), .A2(n1202), .A3(n1203), .A4(n1060), .ZN(n1143) );
NAND2_X1 U857 ( .A1(n1027), .A2(n1204), .ZN(n1197) );
NAND4_X1 U858 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NAND4_X1 U859 ( .A1(n1209), .A2(n1078), .A3(n1068), .A4(n1203), .ZN(n1208) );
XNOR2_X1 U860 ( .A(n1030), .B(KEYINPUT29), .ZN(n1209) );
NAND2_X1 U861 ( .A1(n1028), .A2(n1210), .ZN(n1207) );
AND3_X1 U862 ( .A1(n1060), .A2(n1067), .A3(n1203), .ZN(n1028) );
XNOR2_X1 U863 ( .A(KEYINPUT13), .B(n1211), .ZN(n1206) );
XNOR2_X1 U864 ( .A(KEYINPUT61), .B(n1212), .ZN(n1205) );
NOR2_X1 U865 ( .A1(n1086), .A2(G952), .ZN(n1035) );
XNOR2_X1 U866 ( .A(G146), .B(n1213), .ZN(G48) );
NAND3_X1 U867 ( .A1(n1189), .A2(n1027), .A3(KEYINPUT59), .ZN(n1213) );
AND3_X1 U868 ( .A1(n1190), .A2(n1066), .A3(n1193), .ZN(n1189) );
XNOR2_X1 U869 ( .A(G143), .B(n1214), .ZN(G45) );
NAND2_X1 U870 ( .A1(n1215), .A2(n1027), .ZN(n1214) );
XOR2_X1 U871 ( .A(n1187), .B(KEYINPUT8), .Z(n1215) );
NAND4_X1 U872 ( .A1(n1193), .A2(n1078), .A3(n1042), .A4(n1216), .ZN(n1187) );
XNOR2_X1 U873 ( .A(G140), .B(n1179), .ZN(G42) );
NAND3_X1 U874 ( .A1(n1066), .A2(n1079), .A3(n1196), .ZN(n1179) );
XOR2_X1 U875 ( .A(n1182), .B(n1217), .Z(G39) );
NAND2_X1 U876 ( .A1(KEYINPUT43), .A2(G137), .ZN(n1217) );
NAND3_X1 U877 ( .A1(n1190), .A2(n1068), .A3(n1196), .ZN(n1182) );
XNOR2_X1 U878 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U879 ( .A1(n1078), .A2(n1067), .A3(n1196), .ZN(n1184) );
NOR2_X1 U880 ( .A1(n1218), .A2(n1080), .ZN(n1196) );
XOR2_X1 U881 ( .A(G131), .B(n1219), .Z(G33) );
NOR3_X1 U882 ( .A1(n1220), .A2(n1080), .A3(n1221), .ZN(n1219) );
XNOR2_X1 U883 ( .A(KEYINPUT47), .B(n1070), .ZN(n1221) );
NAND2_X1 U884 ( .A1(n1084), .A2(n1222), .ZN(n1080) );
NAND3_X1 U885 ( .A1(n1078), .A2(n1195), .A3(n1066), .ZN(n1220) );
XNOR2_X1 U886 ( .A(G128), .B(n1223), .ZN(G30) );
NAND4_X1 U887 ( .A1(n1224), .A2(n1193), .A3(n1190), .A4(n1067), .ZN(n1223) );
INV_X1 U888 ( .A(n1218), .ZN(n1193) );
NAND2_X1 U889 ( .A1(n1203), .A2(n1195), .ZN(n1218) );
XNOR2_X1 U890 ( .A(n1027), .B(KEYINPUT48), .ZN(n1224) );
XNOR2_X1 U891 ( .A(G101), .B(n1225), .ZN(G3) );
NAND3_X1 U892 ( .A1(n1226), .A2(n1078), .A3(n1227), .ZN(n1225) );
NOR3_X1 U893 ( .A1(n1228), .A2(n1030), .A3(n1070), .ZN(n1227) );
INV_X1 U894 ( .A(n1203), .ZN(n1070) );
XNOR2_X1 U895 ( .A(n1027), .B(KEYINPUT58), .ZN(n1226) );
XNOR2_X1 U896 ( .A(G125), .B(n1183), .ZN(G27) );
NAND4_X1 U897 ( .A1(n1066), .A2(n1079), .A3(n1229), .A4(n1037), .ZN(n1183) );
AND2_X1 U898 ( .A1(n1195), .A2(n1027), .ZN(n1229) );
NAND2_X1 U899 ( .A1(n1085), .A2(n1230), .ZN(n1195) );
NAND4_X1 U900 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1091), .ZN(n1230) );
INV_X1 U901 ( .A(G900), .ZN(n1091) );
XNOR2_X1 U902 ( .A(n1232), .B(n1233), .ZN(G24) );
NOR2_X1 U903 ( .A1(n1082), .A2(n1211), .ZN(n1233) );
NAND4_X1 U904 ( .A1(n1037), .A2(n1060), .A3(n1234), .A4(n1042), .ZN(n1211) );
NOR2_X1 U905 ( .A1(n1030), .A2(n1235), .ZN(n1234) );
NOR2_X1 U906 ( .A1(n1236), .A2(n1043), .ZN(n1060) );
XOR2_X1 U907 ( .A(n1237), .B(n1238), .Z(G21) );
XNOR2_X1 U908 ( .A(KEYINPUT24), .B(n1239), .ZN(n1238) );
NOR2_X1 U909 ( .A1(n1082), .A2(n1212), .ZN(n1237) );
NAND4_X1 U910 ( .A1(n1190), .A2(n1068), .A3(n1037), .A4(n1210), .ZN(n1212) );
AND2_X1 U911 ( .A1(n1043), .A2(n1236), .ZN(n1190) );
XOR2_X1 U912 ( .A(G116), .B(n1199), .Z(G18) );
AND2_X1 U913 ( .A1(n1240), .A2(n1067), .ZN(n1199) );
NOR2_X1 U914 ( .A1(n1042), .A2(n1235), .ZN(n1067) );
INV_X1 U915 ( .A(n1216), .ZN(n1235) );
XNOR2_X1 U916 ( .A(n1051), .B(KEYINPUT25), .ZN(n1216) );
XOR2_X1 U917 ( .A(n1201), .B(n1241), .Z(G15) );
XOR2_X1 U918 ( .A(KEYINPUT6), .B(G113), .Z(n1241) );
AND2_X1 U919 ( .A1(n1066), .A2(n1240), .ZN(n1201) );
AND3_X1 U920 ( .A1(n1202), .A2(n1037), .A3(n1078), .ZN(n1240) );
NOR2_X1 U921 ( .A1(n1236), .A2(n1242), .ZN(n1078) );
AND2_X1 U922 ( .A1(n1073), .A2(n1243), .ZN(n1037) );
AND2_X1 U923 ( .A1(n1051), .A2(n1042), .ZN(n1066) );
XOR2_X1 U924 ( .A(G110), .B(n1200), .Z(G12) );
AND4_X1 U925 ( .A1(n1068), .A2(n1202), .A3(n1079), .A4(n1203), .ZN(n1200) );
NOR2_X1 U926 ( .A1(n1073), .A2(n1072), .ZN(n1203) );
INV_X1 U927 ( .A(n1243), .ZN(n1072) );
NAND2_X1 U928 ( .A1(G221), .A2(n1244), .ZN(n1243) );
NAND2_X1 U929 ( .A1(G234), .A2(n1177), .ZN(n1244) );
XNOR2_X1 U930 ( .A(n1245), .B(n1246), .ZN(n1073) );
XOR2_X1 U931 ( .A(KEYINPUT42), .B(G469), .Z(n1246) );
NAND2_X1 U932 ( .A1(n1247), .A2(n1177), .ZN(n1245) );
XNOR2_X1 U933 ( .A(n1161), .B(n1248), .ZN(n1247) );
NOR2_X1 U934 ( .A1(KEYINPUT23), .A2(n1249), .ZN(n1248) );
XNOR2_X1 U935 ( .A(G140), .B(n1163), .ZN(n1249) );
XOR2_X1 U936 ( .A(G110), .B(n1250), .Z(n1163) );
NOR2_X1 U937 ( .A1(G953), .A2(n1090), .ZN(n1250) );
INV_X1 U938 ( .A(G227), .ZN(n1090) );
XOR2_X1 U939 ( .A(n1251), .B(n1102), .Z(n1161) );
XOR2_X1 U940 ( .A(n1252), .B(n1253), .Z(n1102) );
XNOR2_X1 U941 ( .A(n1254), .B(n1255), .ZN(n1251) );
INV_X1 U942 ( .A(n1155), .ZN(n1255) );
NAND3_X1 U943 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1254) );
NAND2_X1 U944 ( .A1(G101), .A2(n1259), .ZN(n1258) );
OR3_X1 U945 ( .A1(n1259), .A2(G101), .A3(KEYINPUT15), .ZN(n1257) );
OR2_X1 U946 ( .A1(KEYINPUT49), .A2(n1260), .ZN(n1259) );
NAND2_X1 U947 ( .A1(KEYINPUT15), .A2(n1260), .ZN(n1256) );
XNOR2_X1 U948 ( .A(G104), .B(G107), .ZN(n1260) );
AND2_X1 U949 ( .A1(n1242), .A2(n1236), .ZN(n1079) );
NAND2_X1 U950 ( .A1(n1050), .A2(n1049), .ZN(n1236) );
NAND3_X1 U951 ( .A1(n1261), .A2(n1177), .A3(n1262), .ZN(n1049) );
INV_X1 U952 ( .A(n1126), .ZN(n1262) );
NAND2_X1 U953 ( .A1(G217), .A2(n1263), .ZN(n1261) );
NAND2_X1 U954 ( .A1(G217), .A2(n1264), .ZN(n1050) );
NAND2_X1 U955 ( .A1(n1265), .A2(n1177), .ZN(n1264) );
NAND2_X1 U956 ( .A1(n1126), .A2(n1263), .ZN(n1265) );
XNOR2_X1 U957 ( .A(n1266), .B(n1267), .ZN(n1126) );
XOR2_X1 U958 ( .A(G137), .B(n1268), .Z(n1267) );
NOR2_X1 U959 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U960 ( .A(n1271), .B(KEYINPUT14), .Z(n1270) );
NAND2_X1 U961 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U962 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
AND3_X1 U963 ( .A1(n1276), .A2(n1274), .A3(n1275), .ZN(n1269) );
NAND2_X1 U964 ( .A1(G146), .A2(n1277), .ZN(n1275) );
NAND2_X1 U965 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
INV_X1 U966 ( .A(KEYINPUT53), .ZN(n1279) );
NAND2_X1 U967 ( .A1(n1101), .A2(KEYINPUT33), .ZN(n1278) );
INV_X1 U968 ( .A(n1280), .ZN(n1101) );
NAND2_X1 U969 ( .A1(n1280), .A2(n1281), .ZN(n1274) );
NAND2_X1 U970 ( .A1(KEYINPUT33), .A2(n1282), .ZN(n1281) );
OR2_X1 U971 ( .A1(KEYINPUT53), .A2(G146), .ZN(n1282) );
XOR2_X1 U972 ( .A(G125), .B(G140), .Z(n1280) );
INV_X1 U973 ( .A(n1272), .ZN(n1276) );
XNOR2_X1 U974 ( .A(G110), .B(n1283), .ZN(n1272) );
XNOR2_X1 U975 ( .A(n1252), .B(G119), .ZN(n1283) );
NAND2_X1 U976 ( .A1(n1284), .A2(G221), .ZN(n1266) );
INV_X1 U977 ( .A(n1043), .ZN(n1242) );
XNOR2_X1 U978 ( .A(n1285), .B(G472), .ZN(n1043) );
NAND2_X1 U979 ( .A1(n1286), .A2(n1177), .ZN(n1285) );
XNOR2_X1 U980 ( .A(n1287), .B(n1288), .ZN(n1286) );
INV_X1 U981 ( .A(n1145), .ZN(n1288) );
XOR2_X1 U982 ( .A(n1289), .B(n1290), .Z(n1145) );
INV_X1 U983 ( .A(G101), .ZN(n1290) );
NAND3_X1 U984 ( .A1(n1291), .A2(n1292), .A3(G210), .ZN(n1289) );
XNOR2_X1 U985 ( .A(KEYINPUT36), .B(n1086), .ZN(n1291) );
NAND2_X1 U986 ( .A1(n1293), .A2(KEYINPUT22), .ZN(n1287) );
XOR2_X1 U987 ( .A(n1156), .B(n1294), .Z(n1293) );
XNOR2_X1 U988 ( .A(n1295), .B(n1155), .ZN(n1294) );
XNOR2_X1 U989 ( .A(n1296), .B(G131), .ZN(n1155) );
NAND3_X1 U990 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1296) );
NAND2_X1 U991 ( .A1(G137), .A2(n1300), .ZN(n1299) );
OR3_X1 U992 ( .A1(n1300), .A2(G137), .A3(KEYINPUT38), .ZN(n1298) );
OR2_X1 U993 ( .A1(G134), .A2(KEYINPUT55), .ZN(n1300) );
NAND2_X1 U994 ( .A1(KEYINPUT38), .A2(G134), .ZN(n1297) );
NAND2_X1 U995 ( .A1(KEYINPUT16), .A2(n1152), .ZN(n1295) );
XOR2_X1 U996 ( .A(n1301), .B(n1302), .Z(n1156) );
XNOR2_X1 U997 ( .A(KEYINPUT18), .B(n1239), .ZN(n1302) );
XOR2_X1 U998 ( .A(n1303), .B(G113), .Z(n1301) );
NAND2_X1 U999 ( .A1(KEYINPUT7), .A2(n1304), .ZN(n1303) );
NOR2_X1 U1000 ( .A1(n1082), .A2(n1030), .ZN(n1202) );
INV_X1 U1001 ( .A(n1210), .ZN(n1030) );
NAND2_X1 U1002 ( .A1(n1085), .A2(n1305), .ZN(n1210) );
NAND4_X1 U1003 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1124), .ZN(n1305) );
INV_X1 U1004 ( .A(G898), .ZN(n1124) );
NAND3_X1 U1005 ( .A1(n1231), .A2(n1086), .A3(G952), .ZN(n1085) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1231) );
INV_X1 U1007 ( .A(n1027), .ZN(n1082) );
NOR2_X1 U1008 ( .A1(n1084), .A2(n1040), .ZN(n1027) );
INV_X1 U1009 ( .A(n1222), .ZN(n1040) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1306), .ZN(n1222) );
XNOR2_X1 U1011 ( .A(n1044), .B(n1307), .ZN(n1084) );
NOR2_X1 U1012 ( .A1(n1046), .A2(KEYINPUT50), .ZN(n1307) );
AND2_X1 U1013 ( .A1(n1308), .A2(n1177), .ZN(n1046) );
XNOR2_X1 U1014 ( .A(n1169), .B(n1309), .ZN(n1308) );
XNOR2_X1 U1015 ( .A(n1173), .B(n1172), .ZN(n1309) );
XNOR2_X1 U1016 ( .A(n1152), .B(G125), .ZN(n1172) );
XNOR2_X1 U1017 ( .A(n1310), .B(n1253), .ZN(n1152) );
NAND2_X1 U1018 ( .A1(KEYINPUT60), .A2(n1252), .ZN(n1310) );
AND2_X1 U1019 ( .A1(G224), .A2(n1086), .ZN(n1173) );
XNOR2_X1 U1020 ( .A(n1311), .B(n1123), .ZN(n1169) );
XNOR2_X1 U1021 ( .A(n1312), .B(n1313), .ZN(n1123) );
XNOR2_X1 U1022 ( .A(n1304), .B(n1314), .ZN(n1313) );
XOR2_X1 U1023 ( .A(n1315), .B(n1316), .Z(n1312) );
NOR2_X1 U1024 ( .A1(KEYINPUT3), .A2(n1239), .ZN(n1316) );
INV_X1 U1025 ( .A(G119), .ZN(n1239) );
XNOR2_X1 U1026 ( .A(G101), .B(G107), .ZN(n1315) );
NAND2_X1 U1027 ( .A1(KEYINPUT51), .A2(n1317), .ZN(n1311) );
INV_X1 U1028 ( .A(n1122), .ZN(n1317) );
NAND2_X1 U1029 ( .A1(n1318), .A2(n1319), .ZN(n1122) );
NAND2_X1 U1030 ( .A1(G110), .A2(n1232), .ZN(n1319) );
XOR2_X1 U1031 ( .A(KEYINPUT34), .B(n1320), .Z(n1318) );
NOR2_X1 U1032 ( .A1(G110), .A2(n1232), .ZN(n1320) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1306), .ZN(n1044) );
NAND2_X1 U1034 ( .A1(n1292), .A2(n1177), .ZN(n1306) );
INV_X1 U1035 ( .A(n1228), .ZN(n1068) );
NAND2_X1 U1036 ( .A1(n1321), .A2(n1051), .ZN(n1228) );
XOR2_X1 U1037 ( .A(n1322), .B(G478), .Z(n1051) );
NAND2_X1 U1038 ( .A1(n1323), .A2(n1177), .ZN(n1322) );
XNOR2_X1 U1039 ( .A(n1135), .B(n1136), .ZN(n1323) );
XOR2_X1 U1040 ( .A(G107), .B(n1324), .Z(n1136) );
XNOR2_X1 U1041 ( .A(G143), .B(n1252), .ZN(n1324) );
INV_X1 U1042 ( .A(G128), .ZN(n1252) );
XNOR2_X1 U1043 ( .A(n1325), .B(n1326), .ZN(n1135) );
XOR2_X1 U1044 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1045 ( .A1(n1284), .A2(G217), .ZN(n1328) );
NOR2_X1 U1046 ( .A1(n1263), .A2(G953), .ZN(n1284) );
INV_X1 U1047 ( .A(G234), .ZN(n1263) );
NAND2_X1 U1048 ( .A1(n1329), .A2(n1330), .ZN(n1327) );
NAND2_X1 U1049 ( .A1(n1331), .A2(n1304), .ZN(n1330) );
XOR2_X1 U1050 ( .A(KEYINPUT21), .B(n1332), .Z(n1329) );
NOR2_X1 U1051 ( .A1(n1304), .A2(n1331), .ZN(n1332) );
XNOR2_X1 U1052 ( .A(KEYINPUT19), .B(G122), .ZN(n1331) );
XNOR2_X1 U1053 ( .A(G116), .B(KEYINPUT44), .ZN(n1304) );
NAND2_X1 U1054 ( .A1(KEYINPUT35), .A2(G134), .ZN(n1325) );
XNOR2_X1 U1055 ( .A(n1042), .B(KEYINPUT62), .ZN(n1321) );
XNOR2_X1 U1056 ( .A(n1333), .B(G475), .ZN(n1042) );
NAND2_X1 U1057 ( .A1(n1141), .A2(n1177), .ZN(n1333) );
INV_X1 U1058 ( .A(G902), .ZN(n1177) );
XOR2_X1 U1059 ( .A(n1334), .B(n1335), .Z(n1141) );
XOR2_X1 U1060 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1061 ( .A(G131), .B(n1232), .ZN(n1337) );
INV_X1 U1062 ( .A(G122), .ZN(n1232) );
NOR3_X1 U1063 ( .A1(n1338), .A2(KEYINPUT31), .A3(n1339), .ZN(n1336) );
NOR2_X1 U1064 ( .A1(G140), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1065 ( .A(KEYINPUT4), .B(n1341), .ZN(n1340) );
XOR2_X1 U1066 ( .A(n1342), .B(KEYINPUT39), .Z(n1338) );
NAND2_X1 U1067 ( .A1(G140), .A2(n1341), .ZN(n1342) );
INV_X1 U1068 ( .A(G125), .ZN(n1341) );
XOR2_X1 U1069 ( .A(n1343), .B(n1314), .Z(n1334) );
XOR2_X1 U1070 ( .A(G104), .B(G113), .Z(n1314) );
XOR2_X1 U1071 ( .A(n1344), .B(n1253), .Z(n1343) );
XOR2_X1 U1072 ( .A(G143), .B(G146), .Z(n1253) );
NAND3_X1 U1073 ( .A1(n1292), .A2(n1086), .A3(G214), .ZN(n1344) );
INV_X1 U1074 ( .A(G953), .ZN(n1086) );
INV_X1 U1075 ( .A(G237), .ZN(n1292) );
endmodule


