//Key = 1100010001101010110010110111011000101110001010000011011100110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;

XNOR2_X1 U767 ( .A(n1069), .B(n1070), .ZN(G9) );
NAND2_X1 U768 ( .A1(KEYINPUT0), .A2(G107), .ZN(n1070) );
NOR2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(G75) );
NOR4_X1 U770 ( .A1(G953), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR4_X1 U774 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1081) );
NOR2_X1 U775 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1085) );
XOR2_X1 U777 ( .A(KEYINPUT38), .B(n1091), .Z(n1090) );
INV_X1 U778 ( .A(n1092), .ZN(n1089) );
NOR3_X1 U779 ( .A1(n1093), .A2(KEYINPUT20), .A3(n1094), .ZN(n1084) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1096), .ZN(n1083) );
NOR3_X1 U781 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1095) );
AND3_X1 U782 ( .A1(KEYINPUT25), .A2(n1100), .A3(n1101), .ZN(n1099) );
NOR2_X1 U783 ( .A1(KEYINPUT25), .A2(n1088), .ZN(n1098) );
AND2_X1 U784 ( .A1(n1102), .A2(KEYINPUT20), .ZN(n1097) );
NOR3_X1 U785 ( .A1(n1088), .A2(n1103), .A3(n1096), .ZN(n1078) );
INV_X1 U786 ( .A(n1093), .ZN(n1096) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1082), .ZN(n1105) );
INV_X1 U789 ( .A(n1107), .ZN(n1082) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
AND2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1080), .ZN(n1104) );
INV_X1 U793 ( .A(n1113), .ZN(n1080) );
NOR2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR3_X1 U796 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1071) );
AND4_X1 U797 ( .A1(n1111), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1073) );
NOR4_X1 U798 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U800 ( .A(n1127), .B(KEYINPUT3), .Z(n1126) );
XOR2_X1 U801 ( .A(n1128), .B(KEYINPUT7), .Z(n1122) );
NAND2_X1 U802 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U803 ( .A(n1131), .B(KEYINPUT12), .Z(n1121) );
NOR3_X1 U804 ( .A1(n1132), .A2(n1133), .A3(n1101), .ZN(n1119) );
NAND2_X1 U805 ( .A1(n1134), .A2(n1135), .ZN(n1118) );
XOR2_X1 U806 ( .A(n1136), .B(n1137), .Z(G72) );
NAND2_X1 U807 ( .A1(G953), .A2(n1138), .ZN(n1137) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1138) );
NAND2_X1 U809 ( .A1(KEYINPUT16), .A2(n1139), .ZN(n1136) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U811 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
INV_X1 U812 ( .A(n1144), .ZN(n1143) );
XOR2_X1 U813 ( .A(n1145), .B(n1146), .Z(n1142) );
XOR2_X1 U814 ( .A(G125), .B(n1147), .Z(n1146) );
XOR2_X1 U815 ( .A(n1148), .B(n1149), .Z(n1145) );
NAND2_X1 U816 ( .A1(n1150), .A2(n1151), .ZN(n1140) );
NAND3_X1 U817 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
NAND2_X1 U818 ( .A1(n1155), .A2(n1156), .ZN(G69) );
NAND2_X1 U819 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U820 ( .A(n1159), .ZN(n1157) );
NAND2_X1 U821 ( .A1(n1159), .A2(n1160), .ZN(n1155) );
NAND2_X1 U822 ( .A1(n1161), .A2(n1158), .ZN(n1160) );
NAND2_X1 U823 ( .A1(G953), .A2(n1162), .ZN(n1158) );
XOR2_X1 U824 ( .A(n1163), .B(n1164), .Z(n1159) );
NOR2_X1 U825 ( .A1(n1165), .A2(G953), .ZN(n1164) );
NOR2_X1 U826 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U827 ( .A1(n1168), .A2(n1161), .ZN(n1163) );
INV_X1 U828 ( .A(n1169), .ZN(n1161) );
XOR2_X1 U829 ( .A(n1170), .B(n1171), .Z(n1168) );
XOR2_X1 U830 ( .A(n1172), .B(n1173), .Z(n1170) );
NOR2_X1 U831 ( .A1(KEYINPUT60), .A2(n1174), .ZN(n1173) );
NOR2_X1 U832 ( .A1(n1175), .A2(n1176), .ZN(G66) );
XOR2_X1 U833 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U834 ( .A1(n1179), .A2(G217), .ZN(n1177) );
NOR3_X1 U835 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G63) );
NOR3_X1 U836 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
AND2_X1 U837 ( .A1(n1183), .A2(n1175), .ZN(n1181) );
INV_X1 U838 ( .A(KEYINPUT21), .ZN(n1183) );
NOR3_X1 U839 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1180) );
NOR3_X1 U840 ( .A1(n1189), .A2(n1127), .A3(n1190), .ZN(n1188) );
NOR2_X1 U841 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
AND2_X1 U842 ( .A1(n1075), .A2(G478), .ZN(n1191) );
NOR2_X1 U843 ( .A1(n1175), .A2(n1193), .ZN(G60) );
XNOR2_X1 U844 ( .A(n1194), .B(n1195), .ZN(n1193) );
NAND3_X1 U845 ( .A1(n1179), .A2(G475), .A3(KEYINPUT50), .ZN(n1194) );
XNOR2_X1 U846 ( .A(G104), .B(n1196), .ZN(G6) );
NOR2_X1 U847 ( .A1(n1175), .A2(n1197), .ZN(G57) );
NOR2_X1 U848 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U849 ( .A(n1200), .B(KEYINPUT62), .Z(n1199) );
NAND2_X1 U850 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NOR2_X1 U851 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
AND2_X1 U852 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND2_X1 U853 ( .A1(n1205), .A2(G101), .ZN(n1204) );
NAND2_X1 U854 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
XOR2_X1 U855 ( .A(n1208), .B(KEYINPUT6), .Z(n1206) );
XOR2_X1 U856 ( .A(n1209), .B(n1210), .Z(n1201) );
XOR2_X1 U857 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U858 ( .A1(n1179), .A2(G472), .ZN(n1211) );
INV_X1 U859 ( .A(n1190), .ZN(n1179) );
XNOR2_X1 U860 ( .A(n1213), .B(n1214), .ZN(n1209) );
NAND2_X1 U861 ( .A1(KEYINPUT58), .A2(n1215), .ZN(n1214) );
NAND2_X1 U862 ( .A1(KEYINPUT14), .A2(n1216), .ZN(n1213) );
NOR3_X1 U863 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(G54) );
AND2_X1 U864 ( .A1(n1175), .A2(KEYINPUT23), .ZN(n1219) );
NOR3_X1 U865 ( .A1(KEYINPUT23), .A2(n1184), .A3(n1185), .ZN(n1218) );
XOR2_X1 U866 ( .A(n1220), .B(n1221), .Z(n1217) );
XNOR2_X1 U867 ( .A(n1222), .B(n1223), .ZN(n1221) );
NOR3_X1 U868 ( .A1(n1190), .A2(KEYINPUT32), .A3(n1224), .ZN(n1223) );
INV_X1 U869 ( .A(G469), .ZN(n1224) );
NAND2_X1 U870 ( .A1(n1225), .A2(KEYINPUT5), .ZN(n1222) );
XOR2_X1 U871 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U872 ( .A1(G110), .A2(KEYINPUT46), .ZN(n1227) );
XNOR2_X1 U873 ( .A(G140), .B(n1228), .ZN(n1226) );
NOR2_X1 U874 ( .A1(n1175), .A2(n1229), .ZN(G51) );
XNOR2_X1 U875 ( .A(n1230), .B(n1231), .ZN(n1229) );
XOR2_X1 U876 ( .A(n1232), .B(n1233), .Z(n1230) );
NOR3_X1 U877 ( .A1(n1190), .A2(KEYINPUT19), .A3(n1234), .ZN(n1233) );
NAND2_X1 U878 ( .A1(G902), .A2(n1075), .ZN(n1190) );
NAND4_X1 U879 ( .A1(n1152), .A2(n1235), .A3(n1154), .A4(n1236), .ZN(n1075) );
NOR2_X1 U880 ( .A1(n1167), .A2(n1237), .ZN(n1236) );
XOR2_X1 U881 ( .A(KEYINPUT11), .B(n1166), .Z(n1237) );
NAND4_X1 U882 ( .A1(n1196), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1167) );
NOR4_X1 U883 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1069), .ZN(n1240) );
AND3_X1 U884 ( .A1(n1092), .A2(n1113), .A3(n1244), .ZN(n1069) );
NAND2_X1 U885 ( .A1(n1245), .A2(n1102), .ZN(n1239) );
XOR2_X1 U886 ( .A(n1246), .B(KEYINPUT37), .Z(n1245) );
NAND3_X1 U887 ( .A1(n1244), .A2(n1113), .A3(n1247), .ZN(n1196) );
AND4_X1 U888 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1154) );
NAND2_X1 U889 ( .A1(n1252), .A2(n1092), .ZN(n1248) );
XNOR2_X1 U890 ( .A(KEYINPUT53), .B(n1153), .ZN(n1235) );
AND3_X1 U891 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1152) );
NAND2_X1 U892 ( .A1(n1252), .A2(n1247), .ZN(n1255) );
NAND2_X1 U893 ( .A1(n1102), .A2(n1256), .ZN(n1253) );
XNOR2_X1 U894 ( .A(KEYINPUT35), .B(n1257), .ZN(n1256) );
NAND3_X1 U895 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1232) );
NAND2_X1 U896 ( .A1(KEYINPUT10), .A2(n1261), .ZN(n1259) );
NAND2_X1 U897 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U898 ( .A1(n1264), .A2(n1265), .ZN(n1258) );
INV_X1 U899 ( .A(KEYINPUT10), .ZN(n1265) );
XOR2_X1 U900 ( .A(n1266), .B(n1267), .Z(n1264) );
NAND2_X1 U901 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
NOR2_X1 U902 ( .A1(n1185), .A2(n1270), .ZN(n1175) );
INV_X1 U903 ( .A(n1184), .ZN(n1270) );
XOR2_X1 U904 ( .A(G953), .B(KEYINPUT45), .Z(n1184) );
XOR2_X1 U905 ( .A(G952), .B(KEYINPUT49), .Z(n1185) );
XOR2_X1 U906 ( .A(n1254), .B(n1271), .Z(G48) );
NOR2_X1 U907 ( .A1(G146), .A2(KEYINPUT18), .ZN(n1271) );
NAND4_X1 U908 ( .A1(n1272), .A2(n1247), .A3(n1273), .A4(n1115), .ZN(n1254) );
XOR2_X1 U909 ( .A(n1274), .B(n1275), .Z(G45) );
NOR2_X1 U910 ( .A1(KEYINPUT57), .A2(n1276), .ZN(n1275) );
NOR2_X1 U911 ( .A1(n1094), .A2(n1257), .ZN(n1276) );
NAND4_X1 U912 ( .A1(n1277), .A2(n1109), .A3(n1115), .A4(n1278), .ZN(n1257) );
XOR2_X1 U913 ( .A(n1279), .B(KEYINPUT41), .Z(n1274) );
XNOR2_X1 U914 ( .A(G140), .B(n1153), .ZN(G42) );
NAND4_X1 U915 ( .A1(n1280), .A2(n1247), .A3(n1111), .A4(n1110), .ZN(n1153) );
XOR2_X1 U916 ( .A(n1281), .B(n1249), .Z(G39) );
NAND4_X1 U917 ( .A1(n1273), .A2(n1280), .A3(n1093), .A4(n1110), .ZN(n1249) );
XNOR2_X1 U918 ( .A(G134), .B(n1282), .ZN(G36) );
NAND3_X1 U919 ( .A1(n1252), .A2(n1092), .A3(KEYINPUT54), .ZN(n1282) );
XNOR2_X1 U920 ( .A(G131), .B(n1283), .ZN(G33) );
NAND2_X1 U921 ( .A1(n1252), .A2(n1284), .ZN(n1283) );
XOR2_X1 U922 ( .A(KEYINPUT13), .B(n1247), .Z(n1284) );
AND2_X1 U923 ( .A1(n1280), .A2(n1109), .ZN(n1252) );
AND3_X1 U924 ( .A1(n1115), .A2(n1278), .A3(n1091), .ZN(n1280) );
INV_X1 U925 ( .A(n1088), .ZN(n1091) );
NAND2_X1 U926 ( .A1(n1100), .A2(n1285), .ZN(n1088) );
XOR2_X1 U927 ( .A(n1286), .B(n1250), .Z(G30) );
NAND4_X1 U928 ( .A1(n1273), .A2(n1272), .A3(n1287), .A4(n1092), .ZN(n1250) );
XOR2_X1 U929 ( .A(n1207), .B(n1238), .Z(G3) );
NAND3_X1 U930 ( .A1(n1093), .A2(n1244), .A3(n1109), .ZN(n1238) );
INV_X1 U931 ( .A(G101), .ZN(n1207) );
XOR2_X1 U932 ( .A(n1269), .B(n1251), .Z(G27) );
NAND4_X1 U933 ( .A1(n1272), .A2(n1247), .A3(n1107), .A4(n1111), .ZN(n1251) );
AND3_X1 U934 ( .A1(n1278), .A2(n1110), .A3(n1102), .ZN(n1272) );
NAND2_X1 U935 ( .A1(n1077), .A2(n1288), .ZN(n1278) );
NAND3_X1 U936 ( .A1(G902), .A2(n1289), .A3(n1144), .ZN(n1288) );
NOR2_X1 U937 ( .A1(n1151), .A2(G900), .ZN(n1144) );
XOR2_X1 U938 ( .A(G122), .B(n1290), .Z(G24) );
NOR2_X1 U939 ( .A1(n1094), .A2(n1246), .ZN(n1290) );
NAND4_X1 U940 ( .A1(n1277), .A2(n1113), .A3(n1107), .A4(n1291), .ZN(n1246) );
NOR2_X1 U941 ( .A1(n1110), .A2(n1273), .ZN(n1113) );
AND2_X1 U942 ( .A1(n1292), .A2(n1123), .ZN(n1277) );
XOR2_X1 U943 ( .A(KEYINPUT42), .B(n1293), .Z(n1292) );
INV_X1 U944 ( .A(n1102), .ZN(n1094) );
XOR2_X1 U945 ( .A(G119), .B(n1243), .Z(G21) );
AND4_X1 U946 ( .A1(n1273), .A2(n1294), .A3(n1093), .A4(n1110), .ZN(n1243) );
XOR2_X1 U947 ( .A(n1242), .B(n1295), .Z(G18) );
NOR2_X1 U948 ( .A1(KEYINPUT33), .A2(n1296), .ZN(n1295) );
AND3_X1 U949 ( .A1(n1294), .A2(n1092), .A3(n1109), .ZN(n1242) );
NOR2_X1 U950 ( .A1(n1293), .A2(n1123), .ZN(n1092) );
XOR2_X1 U951 ( .A(G113), .B(n1166), .Z(G15) );
AND3_X1 U952 ( .A1(n1109), .A2(n1294), .A3(n1247), .ZN(n1166) );
INV_X1 U953 ( .A(n1087), .ZN(n1247) );
NAND2_X1 U954 ( .A1(n1123), .A2(n1293), .ZN(n1087) );
INV_X1 U955 ( .A(n1297), .ZN(n1293) );
AND3_X1 U956 ( .A1(n1107), .A2(n1291), .A3(n1102), .ZN(n1294) );
NAND2_X1 U957 ( .A1(n1298), .A2(n1299), .ZN(n1107) );
OR3_X1 U958 ( .A1(n1116), .A2(n1132), .A3(KEYINPUT39), .ZN(n1299) );
INV_X1 U959 ( .A(n1131), .ZN(n1116) );
NAND2_X1 U960 ( .A1(KEYINPUT39), .A2(n1115), .ZN(n1298) );
NOR2_X1 U961 ( .A1(n1111), .A2(n1110), .ZN(n1109) );
XOR2_X1 U962 ( .A(n1241), .B(n1300), .Z(G12) );
NOR2_X1 U963 ( .A1(KEYINPUT8), .A2(n1301), .ZN(n1300) );
AND4_X1 U964 ( .A1(n1093), .A2(n1244), .A3(n1111), .A4(n1110), .ZN(n1241) );
NAND2_X1 U965 ( .A1(n1302), .A2(n1130), .ZN(n1110) );
NAND3_X1 U966 ( .A1(n1303), .A2(n1304), .A3(n1178), .ZN(n1130) );
NAND2_X1 U967 ( .A1(G217), .A2(n1305), .ZN(n1303) );
XNOR2_X1 U968 ( .A(KEYINPUT9), .B(n1129), .ZN(n1302) );
NAND3_X1 U969 ( .A1(n1306), .A2(n1307), .A3(G217), .ZN(n1129) );
NAND2_X1 U970 ( .A1(n1178), .A2(n1304), .ZN(n1306) );
XOR2_X1 U971 ( .A(n1308), .B(n1309), .Z(n1178) );
XNOR2_X1 U972 ( .A(n1149), .B(n1310), .ZN(n1309) );
XOR2_X1 U973 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U974 ( .A(G137), .B(G140), .Z(n1149) );
XOR2_X1 U975 ( .A(n1313), .B(n1314), .Z(n1308) );
XOR2_X1 U976 ( .A(n1301), .B(n1315), .Z(n1314) );
NAND3_X1 U977 ( .A1(n1316), .A2(n1151), .A3(G221), .ZN(n1315) );
NAND2_X1 U978 ( .A1(KEYINPUT27), .A2(G125), .ZN(n1313) );
INV_X1 U979 ( .A(n1273), .ZN(n1111) );
XOR2_X1 U980 ( .A(n1317), .B(n1318), .Z(n1273) );
XOR2_X1 U981 ( .A(KEYINPUT30), .B(G472), .Z(n1318) );
NAND2_X1 U982 ( .A1(n1319), .A2(n1304), .ZN(n1317) );
XOR2_X1 U983 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U984 ( .A(n1205), .B(n1215), .Z(n1321) );
NAND2_X1 U985 ( .A1(n1322), .A2(n1323), .ZN(n1215) );
NAND2_X1 U986 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
INV_X1 U987 ( .A(KEYINPUT55), .ZN(n1325) );
NAND2_X1 U988 ( .A1(KEYINPUT55), .A2(n1326), .ZN(n1322) );
INV_X1 U989 ( .A(n1208), .ZN(n1205) );
NAND2_X1 U990 ( .A1(n1327), .A2(G210), .ZN(n1208) );
XOR2_X1 U991 ( .A(n1328), .B(G101), .Z(n1320) );
NAND2_X1 U992 ( .A1(n1329), .A2(KEYINPUT44), .ZN(n1328) );
XOR2_X1 U993 ( .A(n1216), .B(n1212), .Z(n1329) );
AND3_X1 U994 ( .A1(n1287), .A2(n1291), .A3(n1102), .ZN(n1244) );
NOR2_X1 U995 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
NOR2_X1 U996 ( .A1(n1330), .A2(n1133), .ZN(n1100) );
NOR2_X1 U997 ( .A1(n1135), .A2(n1134), .ZN(n1133) );
AND2_X1 U998 ( .A1(n1331), .A2(n1135), .ZN(n1330) );
NAND2_X1 U999 ( .A1(n1332), .A2(n1304), .ZN(n1135) );
XOR2_X1 U1000 ( .A(n1333), .B(n1334), .Z(n1332) );
AND3_X1 U1001 ( .A1(n1263), .A2(n1260), .A3(n1262), .ZN(n1334) );
NAND2_X1 U1002 ( .A1(n1335), .A2(n1269), .ZN(n1262) );
XOR2_X1 U1003 ( .A(n1267), .B(n1268), .Z(n1335) );
OR3_X1 U1004 ( .A1(n1268), .A2(n1267), .A3(n1269), .ZN(n1260) );
INV_X1 U1005 ( .A(G125), .ZN(n1269) );
NAND3_X1 U1006 ( .A1(G125), .A2(n1268), .A3(n1267), .ZN(n1263) );
NOR2_X1 U1007 ( .A1(n1162), .A2(G953), .ZN(n1267) );
INV_X1 U1008 ( .A(G224), .ZN(n1162) );
INV_X1 U1009 ( .A(n1212), .ZN(n1268) );
XOR2_X1 U1010 ( .A(n1336), .B(n1337), .Z(n1212) );
NOR2_X1 U1011 ( .A1(KEYINPUT56), .A2(n1286), .ZN(n1337) );
XOR2_X1 U1012 ( .A(G146), .B(n1279), .Z(n1336) );
NAND2_X1 U1013 ( .A1(KEYINPUT51), .A2(n1231), .ZN(n1333) );
XNOR2_X1 U1014 ( .A(n1338), .B(n1172), .ZN(n1231) );
XOR2_X1 U1015 ( .A(n1301), .B(G122), .Z(n1172) );
NAND2_X1 U1016 ( .A1(n1339), .A2(KEYINPUT26), .ZN(n1338) );
XOR2_X1 U1017 ( .A(n1174), .B(n1171), .Z(n1339) );
XOR2_X1 U1018 ( .A(G101), .B(n1340), .Z(n1171) );
NOR2_X1 U1019 ( .A1(KEYINPUT31), .A2(n1341), .ZN(n1340) );
INV_X1 U1020 ( .A(n1326), .ZN(n1174) );
NOR2_X1 U1021 ( .A1(n1324), .A2(n1342), .ZN(n1326) );
AND2_X1 U1022 ( .A1(n1343), .A2(G113), .ZN(n1342) );
NOR2_X1 U1023 ( .A1(n1343), .A2(G113), .ZN(n1324) );
XOR2_X1 U1024 ( .A(n1296), .B(n1311), .Z(n1343) );
XOR2_X1 U1025 ( .A(G119), .B(KEYINPUT22), .Z(n1311) );
INV_X1 U1026 ( .A(G116), .ZN(n1296) );
XOR2_X1 U1027 ( .A(KEYINPUT4), .B(n1134), .Z(n1331) );
INV_X1 U1028 ( .A(n1234), .ZN(n1134) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1344), .ZN(n1234) );
INV_X1 U1030 ( .A(n1285), .ZN(n1101) );
NAND2_X1 U1031 ( .A1(n1345), .A2(n1344), .ZN(n1285) );
NAND2_X1 U1032 ( .A1(n1346), .A2(n1304), .ZN(n1344) );
INV_X1 U1033 ( .A(G237), .ZN(n1346) );
XOR2_X1 U1034 ( .A(KEYINPUT2), .B(G214), .Z(n1345) );
NAND2_X1 U1035 ( .A1(n1077), .A2(n1347), .ZN(n1291) );
NAND3_X1 U1036 ( .A1(n1169), .A2(n1289), .A3(G902), .ZN(n1347) );
NOR2_X1 U1037 ( .A1(G898), .A2(n1151), .ZN(n1169) );
NAND3_X1 U1038 ( .A1(n1289), .A2(n1151), .A3(G952), .ZN(n1077) );
NAND2_X1 U1039 ( .A1(G237), .A2(G234), .ZN(n1289) );
XNOR2_X1 U1040 ( .A(n1115), .B(KEYINPUT59), .ZN(n1287) );
NOR2_X1 U1041 ( .A1(n1131), .A2(n1132), .ZN(n1115) );
INV_X1 U1042 ( .A(n1117), .ZN(n1132) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1307), .ZN(n1117) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1304), .ZN(n1307) );
XOR2_X1 U1045 ( .A(n1348), .B(G469), .Z(n1131) );
NAND2_X1 U1046 ( .A1(n1349), .A2(n1304), .ZN(n1348) );
XOR2_X1 U1047 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1048 ( .A(n1220), .B(n1228), .Z(n1351) );
AND2_X1 U1049 ( .A1(G227), .A2(n1151), .ZN(n1228) );
XOR2_X1 U1050 ( .A(n1352), .B(n1353), .Z(n1220) );
XOR2_X1 U1051 ( .A(n1216), .B(n1354), .Z(n1353) );
XOR2_X1 U1052 ( .A(KEYINPUT48), .B(G101), .Z(n1354) );
XOR2_X1 U1053 ( .A(n1147), .B(n1355), .Z(n1216) );
NOR2_X1 U1054 ( .A1(KEYINPUT52), .A2(n1281), .ZN(n1355) );
INV_X1 U1055 ( .A(G137), .ZN(n1281) );
XOR2_X1 U1056 ( .A(G134), .B(G131), .Z(n1147) );
XNOR2_X1 U1057 ( .A(n1148), .B(n1341), .ZN(n1352) );
XNOR2_X1 U1058 ( .A(G104), .B(G107), .ZN(n1341) );
NAND2_X1 U1059 ( .A1(n1356), .A2(n1357), .ZN(n1148) );
NAND2_X1 U1060 ( .A1(n1312), .A2(n1279), .ZN(n1357) );
INV_X1 U1061 ( .A(G143), .ZN(n1279) );
NAND2_X1 U1062 ( .A1(n1358), .A2(G143), .ZN(n1356) );
XNOR2_X1 U1063 ( .A(KEYINPUT61), .B(n1312), .ZN(n1358) );
XOR2_X1 U1064 ( .A(n1286), .B(G146), .Z(n1312) );
INV_X1 U1065 ( .A(G128), .ZN(n1286) );
XOR2_X1 U1066 ( .A(n1301), .B(G140), .Z(n1350) );
INV_X1 U1067 ( .A(G110), .ZN(n1301) );
NOR2_X1 U1068 ( .A1(n1123), .A2(n1297), .ZN(n1093) );
XOR2_X1 U1069 ( .A(n1359), .B(n1186), .Z(n1297) );
INV_X1 U1070 ( .A(n1125), .ZN(n1186) );
NAND2_X1 U1071 ( .A1(n1189), .A2(n1304), .ZN(n1125) );
INV_X1 U1072 ( .A(G902), .ZN(n1304) );
INV_X1 U1073 ( .A(n1192), .ZN(n1189) );
XOR2_X1 U1074 ( .A(n1360), .B(n1361), .Z(n1192) );
XOR2_X1 U1075 ( .A(G128), .B(n1362), .Z(n1361) );
XOR2_X1 U1076 ( .A(G143), .B(G134), .Z(n1362) );
XOR2_X1 U1077 ( .A(n1363), .B(n1364), .Z(n1360) );
AND3_X1 U1078 ( .A1(G217), .A2(n1151), .A3(n1316), .ZN(n1364) );
XNOR2_X1 U1079 ( .A(n1305), .B(KEYINPUT40), .ZN(n1316) );
INV_X1 U1080 ( .A(G234), .ZN(n1305) );
INV_X1 U1081 ( .A(G953), .ZN(n1151) );
NAND2_X1 U1082 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
NAND2_X1 U1083 ( .A1(G107), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1084 ( .A(KEYINPUT36), .B(n1368), .Z(n1365) );
NOR2_X1 U1085 ( .A1(G107), .A2(n1367), .ZN(n1368) );
XOR2_X1 U1086 ( .A(G122), .B(G116), .Z(n1367) );
NAND2_X1 U1087 ( .A1(KEYINPUT29), .A2(n1127), .ZN(n1359) );
INV_X1 U1088 ( .A(G478), .ZN(n1127) );
XNOR2_X1 U1089 ( .A(n1369), .B(n1370), .ZN(n1123) );
NOR2_X1 U1090 ( .A1(n1195), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1091 ( .A(KEYINPUT47), .B(G902), .Z(n1371) );
NAND2_X1 U1092 ( .A1(n1372), .A2(n1373), .ZN(n1195) );
NAND2_X1 U1093 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1094 ( .A1(KEYINPUT34), .A2(n1376), .ZN(n1375) );
NAND2_X1 U1095 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
NAND2_X1 U1096 ( .A1(n1379), .A2(n1380), .ZN(n1372) );
NAND2_X1 U1097 ( .A1(n1378), .A2(n1381), .ZN(n1380) );
NAND2_X1 U1098 ( .A1(KEYINPUT34), .A2(n1382), .ZN(n1381) );
INV_X1 U1099 ( .A(n1374), .ZN(n1382) );
XOR2_X1 U1100 ( .A(n1383), .B(n1384), .Z(n1374) );
XOR2_X1 U1101 ( .A(KEYINPUT28), .B(G122), .Z(n1384) );
XNOR2_X1 U1102 ( .A(G104), .B(G113), .ZN(n1383) );
INV_X1 U1103 ( .A(KEYINPUT43), .ZN(n1378) );
INV_X1 U1104 ( .A(n1377), .ZN(n1379) );
NAND2_X1 U1105 ( .A1(n1385), .A2(n1386), .ZN(n1377) );
OR2_X1 U1106 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XOR2_X1 U1107 ( .A(n1389), .B(KEYINPUT24), .Z(n1385) );
NAND2_X1 U1108 ( .A1(n1388), .A2(n1387), .ZN(n1389) );
NAND2_X1 U1109 ( .A1(n1390), .A2(n1391), .ZN(n1387) );
OR2_X1 U1110 ( .A1(n1392), .A2(G131), .ZN(n1391) );
XOR2_X1 U1111 ( .A(n1393), .B(KEYINPUT15), .Z(n1390) );
NAND2_X1 U1112 ( .A1(G131), .A2(n1392), .ZN(n1393) );
XNOR2_X1 U1113 ( .A(n1394), .B(n1395), .ZN(n1392) );
XOR2_X1 U1114 ( .A(KEYINPUT17), .B(G143), .Z(n1395) );
NAND2_X1 U1115 ( .A1(n1327), .A2(G214), .ZN(n1394) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1327) );
XNOR2_X1 U1117 ( .A(n1396), .B(G146), .ZN(n1388) );
NAND2_X1 U1118 ( .A1(KEYINPUT1), .A2(n1397), .ZN(n1396) );
XOR2_X1 U1119 ( .A(G140), .B(G125), .Z(n1397) );
XNOR2_X1 U1120 ( .A(G475), .B(KEYINPUT63), .ZN(n1369) );
endmodule


