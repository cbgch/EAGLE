//Key = 0110000110010110011001011011110011110110100101011101001110011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329;

XNOR2_X1 U726 ( .A(n1005), .B(n1006), .ZN(G9) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U728 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1008) );
NOR2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR3_X1 U730 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1013) );
NOR3_X1 U731 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
INV_X1 U732 ( .A(KEYINPUT34), .ZN(n1018) );
NOR3_X1 U733 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1016) );
NOR2_X1 U734 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NAND3_X1 U735 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1021) );
NAND4_X1 U736 ( .A1(n1029), .A2(n1030), .A3(n1024), .A4(n1031), .ZN(n1027) );
OR2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1029) );
NAND2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1026) );
XOR2_X1 U739 ( .A(KEYINPUT42), .B(n1036), .Z(n1015) );
NOR2_X1 U740 ( .A1(n1037), .A2(n1020), .ZN(n1036) );
NOR2_X1 U741 ( .A1(KEYINPUT34), .A2(n1038), .ZN(n1011) );
NOR2_X1 U742 ( .A1(n1039), .A2(n1020), .ZN(n1038) );
INV_X1 U743 ( .A(n1040), .ZN(n1039) );
NAND4_X1 U744 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1009) );
NAND3_X1 U745 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1042) );
NAND2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1041) );
XNOR2_X1 U747 ( .A(n1045), .B(KEYINPUT26), .ZN(n1048) );
NOR2_X1 U748 ( .A1(n1020), .A2(n1023), .ZN(n1045) );
NAND3_X1 U749 ( .A1(n1025), .A2(n1024), .A3(n1028), .ZN(n1020) );
INV_X1 U750 ( .A(n1050), .ZN(n1028) );
NOR3_X1 U751 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1007) );
INV_X1 U752 ( .A(n1043), .ZN(n1051) );
NAND4_X1 U753 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1043) );
NOR3_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U756 ( .A1(G469), .A2(KEYINPUT46), .ZN(n1060) );
NOR2_X1 U757 ( .A1(n1061), .A2(n1062), .ZN(n1057) );
NAND3_X1 U758 ( .A1(n1063), .A2(n1064), .A3(n1032), .ZN(n1056) );
NOR3_X1 U759 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1054) );
NOR3_X1 U760 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
AND2_X1 U761 ( .A1(n1068), .A2(n1070), .ZN(n1066) );
INV_X1 U762 ( .A(KEYINPUT59), .ZN(n1068) );
XNOR2_X1 U763 ( .A(n1071), .B(n1072), .ZN(n1065) );
XOR2_X1 U764 ( .A(n1073), .B(n1074), .Z(n1053) );
NOR2_X1 U765 ( .A1(G478), .A2(KEYINPUT6), .ZN(n1074) );
XOR2_X1 U766 ( .A(n1075), .B(n1076), .Z(G72) );
XOR2_X1 U767 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U768 ( .A1(n1079), .A2(n1044), .ZN(n1078) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U770 ( .A1(n1082), .A2(n1083), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1084), .A2(G953), .ZN(n1083) );
XNOR2_X1 U772 ( .A(G900), .B(KEYINPUT44), .ZN(n1084) );
XNOR2_X1 U773 ( .A(n1085), .B(n1086), .ZN(n1082) );
XNOR2_X1 U774 ( .A(n1087), .B(n1088), .ZN(n1086) );
INV_X1 U775 ( .A(G125), .ZN(n1088) );
NAND2_X1 U776 ( .A1(KEYINPUT29), .A2(n1089), .ZN(n1087) );
NAND2_X1 U777 ( .A1(n1044), .A2(n1090), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(G69) );
XOR2_X1 U780 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U782 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND2_X1 U783 ( .A1(KEYINPUT13), .A2(n1101), .ZN(n1095) );
NAND2_X1 U784 ( .A1(G953), .A2(n1102), .ZN(n1101) );
NAND2_X1 U785 ( .A1(G224), .A2(G898), .ZN(n1102) );
NAND2_X1 U786 ( .A1(KEYINPUT8), .A2(n1103), .ZN(n1093) );
NAND2_X1 U787 ( .A1(n1104), .A2(n1044), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U789 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1070), .A2(n1109), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1110), .ZN(G63) );
NOR3_X1 U792 ( .A1(n1073), .A2(n1111), .A3(n1112), .ZN(n1110) );
AND3_X1 U793 ( .A1(n1113), .A2(G902), .A3(n1114), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR3_X1 U795 ( .A1(KEYINPUT36), .A2(n1115), .A3(n1116), .ZN(n1114) );
XNOR2_X1 U796 ( .A(KEYINPUT41), .B(n1010), .ZN(n1116) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1117), .ZN(G60) );
NOR3_X1 U798 ( .A1(n1072), .A2(n1118), .A3(n1119), .ZN(n1117) );
NOR3_X1 U799 ( .A1(n1120), .A2(n1071), .A3(n1109), .ZN(n1119) );
NOR2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
AND2_X1 U801 ( .A1(n1010), .A2(G475), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(G6) );
XNOR2_X1 U803 ( .A(G104), .B(KEYINPUT62), .ZN(n1124) );
NAND4_X1 U804 ( .A1(n1125), .A2(n1024), .A3(n1126), .A4(n1127), .ZN(n1123) );
NAND2_X1 U805 ( .A1(KEYINPUT27), .A2(n1128), .ZN(n1127) );
NAND2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
INV_X1 U807 ( .A(KEYINPUT27), .ZN(n1130) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U809 ( .A1(n1105), .A2(n1133), .ZN(G57) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U812 ( .A(KEYINPUT57), .B(n1138), .Z(n1137) );
NOR2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U814 ( .A(KEYINPUT10), .B(n1141), .ZN(n1140) );
NOR2_X1 U815 ( .A1(n1142), .A2(n1141), .ZN(n1136) );
OR2_X1 U816 ( .A1(n1109), .A2(n1062), .ZN(n1141) );
XNOR2_X1 U817 ( .A(n1139), .B(n1143), .ZN(n1142) );
XOR2_X1 U818 ( .A(KEYINPUT25), .B(KEYINPUT19), .Z(n1143) );
XOR2_X1 U819 ( .A(n1144), .B(n1085), .Z(n1139) );
XNOR2_X1 U820 ( .A(n1145), .B(n1146), .ZN(n1085) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1134) );
INV_X1 U822 ( .A(n1149), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1105), .A2(n1150), .ZN(G54) );
XOR2_X1 U824 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U827 ( .A1(KEYINPUT56), .A2(n1157), .ZN(n1155) );
XOR2_X1 U828 ( .A(n1158), .B(n1159), .Z(n1151) );
XOR2_X1 U829 ( .A(KEYINPUT47), .B(n1160), .Z(n1159) );
NOR2_X1 U830 ( .A1(n1161), .A2(n1109), .ZN(n1160) );
NAND2_X1 U831 ( .A1(G902), .A2(n1010), .ZN(n1109) );
NAND2_X1 U832 ( .A1(KEYINPUT35), .A2(n1162), .ZN(n1158) );
XNOR2_X1 U833 ( .A(n1089), .B(n1163), .ZN(n1162) );
XOR2_X1 U834 ( .A(KEYINPUT53), .B(G110), .Z(n1163) );
NOR2_X1 U835 ( .A1(n1105), .A2(n1164), .ZN(G51) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U838 ( .A1(KEYINPUT14), .A2(n1169), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(KEYINPUT60), .Z(n1165) );
NAND4_X1 U840 ( .A1(G210), .A2(n1010), .A3(n1171), .A4(n1172), .ZN(n1170) );
NAND2_X1 U841 ( .A1(KEYINPUT4), .A2(G902), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND2_X1 U843 ( .A1(KEYINPUT4), .A2(G237), .ZN(n1173) );
NAND3_X1 U844 ( .A1(n1175), .A2(n1091), .A3(n1176), .ZN(n1010) );
XOR2_X1 U845 ( .A(n1092), .B(KEYINPUT31), .Z(n1176) );
AND4_X1 U846 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1091) );
AND4_X1 U847 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
NAND3_X1 U848 ( .A1(n1185), .A2(n1049), .A3(n1186), .ZN(n1179) );
INV_X1 U849 ( .A(n1104), .ZN(n1175) );
NAND4_X1 U850 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1104) );
NOR3_X1 U851 ( .A1(n1191), .A2(n1006), .A3(n1192), .ZN(n1190) );
NOR4_X1 U852 ( .A1(n1030), .A2(n1035), .A3(n1019), .A4(n1193), .ZN(n1006) );
NAND2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1189) );
NAND2_X1 U854 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND4_X1 U855 ( .A1(n1198), .A2(n1035), .A3(n1199), .A4(n1200), .ZN(n1197) );
NAND2_X1 U856 ( .A1(n1201), .A2(n1034), .ZN(n1200) );
NAND2_X1 U857 ( .A1(n1202), .A2(n1030), .ZN(n1199) );
INV_X1 U858 ( .A(n1125), .ZN(n1196) );
NOR3_X1 U859 ( .A1(n1030), .A2(n1035), .A3(n1037), .ZN(n1125) );
NOR2_X1 U860 ( .A1(n1044), .A2(G952), .ZN(n1105) );
XNOR2_X1 U861 ( .A(G146), .B(n1177), .ZN(G48) );
NAND3_X1 U862 ( .A1(n1203), .A2(n1049), .A3(n1204), .ZN(n1177) );
XNOR2_X1 U863 ( .A(G143), .B(n1092), .ZN(G45) );
NAND4_X1 U864 ( .A1(n1205), .A2(n1049), .A3(n1201), .A4(n1206), .ZN(n1092) );
NAND2_X1 U865 ( .A1(n1207), .A2(n1208), .ZN(G42) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U867 ( .A1(G140), .A2(n1211), .ZN(n1210) );
OR2_X1 U868 ( .A1(KEYINPUT16), .A2(KEYINPUT49), .ZN(n1211) );
NAND3_X1 U869 ( .A1(n1212), .A2(n1213), .A3(KEYINPUT49), .ZN(n1207) );
OR2_X1 U870 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1213) );
NAND2_X1 U871 ( .A1(G140), .A2(n1214), .ZN(n1212) );
OR2_X1 U872 ( .A1(n1209), .A2(KEYINPUT16), .ZN(n1214) );
INV_X1 U873 ( .A(n1178), .ZN(n1209) );
NAND3_X1 U874 ( .A1(n1052), .A2(n1215), .A3(n1186), .ZN(n1178) );
XNOR2_X1 U875 ( .A(G137), .B(n1184), .ZN(G39) );
NAND3_X1 U876 ( .A1(n1216), .A2(n1052), .A3(n1204), .ZN(n1184) );
XOR2_X1 U877 ( .A(n1183), .B(n1217), .Z(G36) );
XOR2_X1 U878 ( .A(KEYINPUT40), .B(G134), .Z(n1217) );
NAND2_X1 U879 ( .A1(n1040), .A2(n1205), .ZN(n1183) );
NOR2_X1 U880 ( .A1(n1014), .A2(n1019), .ZN(n1040) );
INV_X1 U881 ( .A(n1218), .ZN(n1019) );
INV_X1 U882 ( .A(n1052), .ZN(n1014) );
XNOR2_X1 U883 ( .A(G131), .B(n1182), .ZN(G33) );
NAND3_X1 U884 ( .A1(n1203), .A2(n1052), .A3(n1205), .ZN(n1182) );
AND4_X1 U885 ( .A1(n1215), .A2(n1024), .A3(n1219), .A4(n1035), .ZN(n1205) );
NOR2_X1 U886 ( .A1(n1220), .A2(n1047), .ZN(n1052) );
XOR2_X1 U887 ( .A(n1181), .B(n1221), .Z(G30) );
NAND2_X1 U888 ( .A1(KEYINPUT38), .A2(G128), .ZN(n1221) );
NAND3_X1 U889 ( .A1(n1218), .A2(n1049), .A3(n1204), .ZN(n1181) );
AND4_X1 U890 ( .A1(n1215), .A2(n1219), .A3(n1222), .A4(n1035), .ZN(n1204) );
XNOR2_X1 U891 ( .A(G101), .B(n1223), .ZN(G3) );
NAND4_X1 U892 ( .A1(KEYINPUT24), .A2(n1216), .A3(n1224), .A4(n1215), .ZN(n1223) );
NOR2_X1 U893 ( .A1(n1031), .A2(n1193), .ZN(n1224) );
XNOR2_X1 U894 ( .A(G125), .B(n1225), .ZN(G27) );
NAND3_X1 U895 ( .A1(n1185), .A2(n1226), .A3(n1186), .ZN(n1225) );
AND4_X1 U896 ( .A1(n1203), .A2(n1031), .A3(n1219), .A4(n1222), .ZN(n1186) );
NAND2_X1 U897 ( .A1(n1050), .A2(n1227), .ZN(n1219) );
NAND4_X1 U898 ( .A1(G902), .A2(G953), .A3(n1228), .A4(n1081), .ZN(n1227) );
INV_X1 U899 ( .A(G900), .ZN(n1081) );
XNOR2_X1 U900 ( .A(KEYINPUT3), .B(n1131), .ZN(n1226) );
XOR2_X1 U901 ( .A(n1187), .B(n1229), .Z(G24) );
NOR2_X1 U902 ( .A1(G122), .A2(KEYINPUT39), .ZN(n1229) );
NAND4_X1 U903 ( .A1(n1025), .A2(n1194), .A3(n1201), .A4(n1206), .ZN(n1187) );
NOR2_X1 U904 ( .A1(n1034), .A2(n1035), .ZN(n1025) );
XNOR2_X1 U905 ( .A(G119), .B(n1188), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1230), .A2(n1035), .A3(n1185), .ZN(n1188) );
XNOR2_X1 U907 ( .A(G116), .B(n1231), .ZN(G18) );
NAND4_X1 U908 ( .A1(n1024), .A2(n1035), .A3(n1218), .A4(n1232), .ZN(n1231) );
NOR3_X1 U909 ( .A1(n1034), .A2(n1233), .A3(n1234), .ZN(n1232) );
NOR2_X1 U910 ( .A1(KEYINPUT21), .A2(n1235), .ZN(n1234) );
AND2_X1 U911 ( .A1(n1132), .A2(n1131), .ZN(n1235) );
INV_X1 U912 ( .A(n1049), .ZN(n1131) );
AND2_X1 U913 ( .A1(n1128), .A2(KEYINPUT21), .ZN(n1233) );
NOR2_X1 U914 ( .A1(n1206), .A2(n1202), .ZN(n1218) );
XOR2_X1 U915 ( .A(G113), .B(n1236), .Z(G15) );
NOR2_X1 U916 ( .A1(KEYINPUT20), .A2(n1237), .ZN(n1236) );
INV_X1 U917 ( .A(n1191), .ZN(n1237) );
NOR4_X1 U918 ( .A1(n1037), .A2(n1034), .A3(n1193), .A4(n1031), .ZN(n1191) );
INV_X1 U919 ( .A(n1194), .ZN(n1193) );
NOR2_X1 U920 ( .A1(n1128), .A2(n1222), .ZN(n1194) );
INV_X1 U921 ( .A(n1185), .ZN(n1034) );
NOR2_X1 U922 ( .A1(n1033), .A2(n1238), .ZN(n1185) );
INV_X1 U923 ( .A(n1032), .ZN(n1238) );
INV_X1 U924 ( .A(n1203), .ZN(n1037) );
NOR2_X1 U925 ( .A1(n1201), .A2(n1198), .ZN(n1203) );
INV_X1 U926 ( .A(n1206), .ZN(n1198) );
XOR2_X1 U927 ( .A(G110), .B(n1192), .Z(G12) );
AND3_X1 U928 ( .A1(n1215), .A2(n1031), .A3(n1230), .ZN(n1192) );
NOR3_X1 U929 ( .A1(n1128), .A2(n1024), .A3(n1023), .ZN(n1230) );
INV_X1 U930 ( .A(n1216), .ZN(n1023) );
NOR2_X1 U931 ( .A1(n1201), .A2(n1206), .ZN(n1216) );
XNOR2_X1 U932 ( .A(n1239), .B(n1240), .ZN(n1206) );
XOR2_X1 U933 ( .A(KEYINPUT37), .B(n1072), .Z(n1240) );
NOR2_X1 U934 ( .A1(n1122), .A2(G902), .ZN(n1072) );
INV_X1 U935 ( .A(n1120), .ZN(n1122) );
XOR2_X1 U936 ( .A(n1241), .B(n1242), .Z(n1120) );
XOR2_X1 U937 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U938 ( .A(G122), .B(G113), .Z(n1244) );
XNOR2_X1 U939 ( .A(n1245), .B(G125), .ZN(n1243) );
INV_X1 U940 ( .A(G131), .ZN(n1245) );
XOR2_X1 U941 ( .A(n1246), .B(n1247), .Z(n1241) );
XNOR2_X1 U942 ( .A(n1089), .B(n1248), .ZN(n1247) );
XNOR2_X1 U943 ( .A(n1249), .B(n1250), .ZN(n1246) );
NAND4_X1 U944 ( .A1(KEYINPUT48), .A2(G214), .A3(n1251), .A4(n1044), .ZN(n1250) );
NAND2_X1 U945 ( .A1(KEYINPUT2), .A2(n1252), .ZN(n1249) );
XOR2_X1 U946 ( .A(KEYINPUT18), .B(G104), .Z(n1252) );
NAND2_X1 U947 ( .A1(KEYINPUT33), .A2(n1071), .ZN(n1239) );
INV_X1 U948 ( .A(G475), .ZN(n1071) );
INV_X1 U949 ( .A(n1202), .ZN(n1201) );
XOR2_X1 U950 ( .A(n1073), .B(n1115), .Z(n1202) );
INV_X1 U951 ( .A(G478), .ZN(n1115) );
NOR2_X1 U952 ( .A1(n1113), .A2(G902), .ZN(n1073) );
AND2_X1 U953 ( .A1(n1253), .A2(n1254), .ZN(n1113) );
NAND3_X1 U954 ( .A1(n1255), .A2(n1256), .A3(G217), .ZN(n1254) );
XNOR2_X1 U955 ( .A(KEYINPUT22), .B(n1257), .ZN(n1256) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1258), .ZN(n1253) );
NAND2_X1 U957 ( .A1(G217), .A2(n1255), .ZN(n1258) );
XOR2_X1 U958 ( .A(n1259), .B(n1260), .Z(n1257) );
XOR2_X1 U959 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U960 ( .A(n1263), .B(n1264), .ZN(n1262) );
NOR2_X1 U961 ( .A1(G134), .A2(KEYINPUT30), .ZN(n1264) );
NAND2_X1 U962 ( .A1(KEYINPUT51), .A2(G128), .ZN(n1263) );
XNOR2_X1 U963 ( .A(G116), .B(n1265), .ZN(n1259) );
XOR2_X1 U964 ( .A(KEYINPUT12), .B(G143), .Z(n1265) );
INV_X1 U965 ( .A(n1222), .ZN(n1024) );
NAND3_X1 U966 ( .A1(n1266), .A2(n1267), .A3(n1063), .ZN(n1222) );
NAND2_X1 U967 ( .A1(n1069), .A2(n1070), .ZN(n1063) );
OR3_X1 U968 ( .A1(n1070), .A2(n1069), .A3(KEYINPUT9), .ZN(n1267) );
NOR2_X1 U969 ( .A1(n1108), .A2(G902), .ZN(n1069) );
XNOR2_X1 U970 ( .A(n1268), .B(n1269), .ZN(n1108) );
XOR2_X1 U971 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND2_X1 U972 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U973 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
INV_X1 U974 ( .A(G128), .ZN(n1275) );
XOR2_X1 U975 ( .A(KEYINPUT52), .B(G119), .Z(n1274) );
NAND2_X1 U976 ( .A1(n1276), .A2(G128), .ZN(n1272) );
XOR2_X1 U977 ( .A(KEYINPUT54), .B(G119), .Z(n1276) );
NAND2_X1 U978 ( .A1(n1277), .A2(n1278), .ZN(n1270) );
NAND3_X1 U979 ( .A1(G137), .A2(G221), .A3(n1255), .ZN(n1278) );
NAND2_X1 U980 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
NAND2_X1 U981 ( .A1(n1255), .A2(G221), .ZN(n1280) );
AND2_X1 U982 ( .A1(G234), .A2(n1044), .ZN(n1255) );
XOR2_X1 U983 ( .A(KEYINPUT17), .B(G137), .Z(n1279) );
XOR2_X1 U984 ( .A(n1281), .B(G110), .Z(n1268) );
NAND2_X1 U985 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U986 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U987 ( .A(KEYINPUT23), .B(n1286), .Z(n1282) );
NOR2_X1 U988 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
XNOR2_X1 U989 ( .A(n1089), .B(n1287), .ZN(n1284) );
NOR2_X1 U990 ( .A1(G125), .A2(KEYINPUT15), .ZN(n1287) );
NAND2_X1 U991 ( .A1(KEYINPUT9), .A2(n1070), .ZN(n1266) );
NAND2_X1 U992 ( .A1(G217), .A2(n1288), .ZN(n1070) );
NAND2_X1 U993 ( .A1(n1049), .A2(n1132), .ZN(n1128) );
NAND2_X1 U994 ( .A1(n1289), .A2(n1050), .ZN(n1132) );
NAND3_X1 U995 ( .A1(n1228), .A2(n1044), .A3(G952), .ZN(n1050) );
NAND3_X1 U996 ( .A1(n1097), .A2(n1228), .A3(G902), .ZN(n1289) );
NAND2_X1 U997 ( .A1(G237), .A2(G234), .ZN(n1228) );
AND2_X1 U998 ( .A1(n1290), .A2(G953), .ZN(n1097) );
XNOR2_X1 U999 ( .A(G898), .B(KEYINPUT5), .ZN(n1290) );
NOR2_X1 U1000 ( .A1(n1046), .A2(n1047), .ZN(n1049) );
AND2_X1 U1001 ( .A1(G214), .A2(n1291), .ZN(n1047) );
NAND2_X1 U1002 ( .A1(n1251), .A2(n1174), .ZN(n1291) );
INV_X1 U1003 ( .A(n1220), .ZN(n1046) );
NAND2_X1 U1004 ( .A1(n1292), .A2(n1293), .ZN(n1220) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1294), .ZN(n1293) );
NAND2_X1 U1006 ( .A1(n1174), .A2(n1295), .ZN(n1294) );
OR2_X1 U1007 ( .A1(n1251), .A2(n1296), .ZN(n1295) );
NAND3_X1 U1008 ( .A1(n1297), .A2(n1174), .A3(n1296), .ZN(n1292) );
XOR2_X1 U1009 ( .A(n1169), .B(n1168), .Z(n1296) );
XNOR2_X1 U1010 ( .A(n1298), .B(n1157), .ZN(n1168) );
XNOR2_X1 U1011 ( .A(G125), .B(n1299), .ZN(n1298) );
AND2_X1 U1012 ( .A1(n1044), .A2(G224), .ZN(n1299) );
XNOR2_X1 U1013 ( .A(n1300), .B(n1301), .ZN(n1169) );
INV_X1 U1014 ( .A(n1099), .ZN(n1301) );
XNOR2_X1 U1015 ( .A(n1302), .B(n1303), .ZN(n1099) );
XOR2_X1 U1016 ( .A(G110), .B(G104), .Z(n1303) );
XOR2_X1 U1017 ( .A(n1304), .B(n1261), .Z(n1302) );
XNOR2_X1 U1018 ( .A(n1005), .B(G122), .ZN(n1261) );
NAND2_X1 U1019 ( .A1(KEYINPUT7), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1020 ( .A1(KEYINPUT32), .A2(n1100), .ZN(n1300) );
INV_X1 U1021 ( .A(n1144), .ZN(n1100) );
NAND2_X1 U1022 ( .A1(G237), .A2(G210), .ZN(n1297) );
INV_X1 U1023 ( .A(n1035), .ZN(n1031) );
NAND3_X1 U1024 ( .A1(n1306), .A2(n1307), .A3(n1064), .ZN(n1035) );
NAND2_X1 U1025 ( .A1(n1061), .A2(n1062), .ZN(n1064) );
INV_X1 U1026 ( .A(G472), .ZN(n1062) );
INV_X1 U1027 ( .A(n1308), .ZN(n1061) );
OR2_X1 U1028 ( .A1(G472), .A2(KEYINPUT43), .ZN(n1307) );
NAND3_X1 U1029 ( .A1(G472), .A2(n1308), .A3(KEYINPUT43), .ZN(n1306) );
NAND2_X1 U1030 ( .A1(n1309), .A2(n1174), .ZN(n1308) );
XOR2_X1 U1031 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1032 ( .A(n1312), .B(n1313), .Z(n1311) );
XNOR2_X1 U1033 ( .A(KEYINPUT11), .B(n1314), .ZN(n1313) );
NOR3_X1 U1034 ( .A1(n1315), .A2(KEYINPUT58), .A3(n1149), .ZN(n1314) );
NOR2_X1 U1035 ( .A1(n1316), .A2(n1317), .ZN(n1149) );
XOR2_X1 U1036 ( .A(n1147), .B(KEYINPUT55), .Z(n1315) );
NAND2_X1 U1037 ( .A1(n1317), .A2(n1316), .ZN(n1147) );
NAND3_X1 U1038 ( .A1(n1251), .A2(n1044), .A3(G210), .ZN(n1316) );
INV_X1 U1039 ( .A(G953), .ZN(n1044) );
INV_X1 U1040 ( .A(G237), .ZN(n1251) );
NAND2_X1 U1041 ( .A1(KEYINPUT45), .A2(n1145), .ZN(n1312) );
XNOR2_X1 U1042 ( .A(n1157), .B(n1144), .ZN(n1310) );
XOR2_X1 U1043 ( .A(G113), .B(n1318), .Z(n1144) );
XOR2_X1 U1044 ( .A(G119), .B(G116), .Z(n1318) );
INV_X1 U1045 ( .A(n1030), .ZN(n1215) );
NAND2_X1 U1046 ( .A1(n1033), .A2(n1032), .ZN(n1030) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1288), .ZN(n1032) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1174), .ZN(n1288) );
XOR2_X1 U1049 ( .A(n1059), .B(n1161), .Z(n1033) );
INV_X1 U1050 ( .A(G469), .ZN(n1161) );
NAND2_X1 U1051 ( .A1(n1319), .A2(n1174), .ZN(n1059) );
INV_X1 U1052 ( .A(G902), .ZN(n1174) );
XOR2_X1 U1053 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1054 ( .A(n1156), .B(n1153), .ZN(n1321) );
XOR2_X1 U1055 ( .A(n1145), .B(n1322), .Z(n1153) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1080), .ZN(n1322) );
INV_X1 U1057 ( .A(G227), .ZN(n1080) );
XOR2_X1 U1058 ( .A(G131), .B(n1323), .Z(n1145) );
XOR2_X1 U1059 ( .A(G137), .B(G134), .Z(n1323) );
XOR2_X1 U1060 ( .A(n1324), .B(n1325), .Z(n1156) );
XOR2_X1 U1061 ( .A(KEYINPUT61), .B(G104), .Z(n1325) );
XNOR2_X1 U1062 ( .A(n1326), .B(n1305), .ZN(n1324) );
XOR2_X1 U1063 ( .A(n1317), .B(KEYINPUT1), .Z(n1305) );
INV_X1 U1064 ( .A(G101), .ZN(n1317) );
NAND2_X1 U1065 ( .A1(KEYINPUT28), .A2(n1005), .ZN(n1326) );
INV_X1 U1066 ( .A(G107), .ZN(n1005) );
XOR2_X1 U1067 ( .A(n1089), .B(n1327), .Z(n1320) );
XNOR2_X1 U1068 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1069 ( .A1(KEYINPUT63), .A2(n1146), .ZN(n1329) );
INV_X1 U1070 ( .A(n1157), .ZN(n1146) );
XOR2_X1 U1071 ( .A(G128), .B(n1248), .Z(n1157) );
XNOR2_X1 U1072 ( .A(G143), .B(n1285), .ZN(n1248) );
INV_X1 U1073 ( .A(G146), .ZN(n1285) );
NOR2_X1 U1074 ( .A1(G110), .A2(KEYINPUT50), .ZN(n1328) );
XNOR2_X1 U1075 ( .A(G140), .B(KEYINPUT0), .ZN(n1089) );
endmodule


