//Key = 0110001101111101100011111111100110011010010010010011100011011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;

XOR2_X1 U762 ( .A(n1060), .B(n1061), .Z(G9) );
NAND4_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(G75) );
NAND3_X1 U764 ( .A1(KEYINPUT45), .A2(n1066), .A3(n1067), .ZN(n1065) );
NAND2_X1 U765 ( .A1(G952), .A2(n1068), .ZN(n1064) );
NAND4_X1 U766 ( .A1(n1066), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1068) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND4_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
NAND2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1078), .A2(n1086), .ZN(n1085) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
OR3_X1 U775 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
XOR2_X1 U777 ( .A(n1091), .B(KEYINPUT38), .Z(n1092) );
NAND2_X1 U778 ( .A1(n1077), .A2(n1094), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U780 ( .A1(n1078), .A2(n1097), .ZN(n1096) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U783 ( .A1(n1076), .A2(n1102), .ZN(n1095) );
NAND2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U786 ( .A(KEYINPUT44), .B(n1107), .Z(n1103) );
INV_X1 U787 ( .A(n1108), .ZN(n1072) );
XOR2_X1 U788 ( .A(KEYINPUT62), .B(n1109), .Z(n1070) );
NAND4_X1 U789 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1063) );
NOR4_X1 U790 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1113) );
XOR2_X1 U791 ( .A(KEYINPUT4), .B(n1118), .Z(n1117) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1119), .ZN(n1112) );
XNOR2_X1 U793 ( .A(n1120), .B(n1121), .ZN(n1119) );
NAND2_X1 U794 ( .A1(KEYINPUT57), .A2(n1122), .ZN(n1120) );
XOR2_X1 U795 ( .A(n1101), .B(n1123), .Z(n1111) );
XNOR2_X1 U796 ( .A(KEYINPUT7), .B(KEYINPUT43), .ZN(n1123) );
XOR2_X1 U797 ( .A(KEYINPUT20), .B(n1124), .Z(n1110) );
OR2_X1 U798 ( .A1(n1066), .A2(KEYINPUT45), .ZN(n1062) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(G72) );
NAND2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U801 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U802 ( .A1(KEYINPUT42), .A2(n1131), .ZN(n1130) );
NAND3_X1 U803 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1125) );
INV_X1 U804 ( .A(KEYINPUT42), .ZN(n1134) );
NAND2_X1 U805 ( .A1(n1135), .A2(n1131), .ZN(n1133) );
INV_X1 U806 ( .A(KEYINPUT17), .ZN(n1131) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1136), .ZN(n1132) );
OR2_X1 U808 ( .A1(n1127), .A2(KEYINPUT17), .ZN(n1136) );
XNOR2_X1 U809 ( .A(n1137), .B(n1138), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1069), .A2(n1139), .ZN(n1138) );
XOR2_X1 U811 ( .A(n1140), .B(KEYINPUT41), .Z(n1139) );
NAND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1137) );
NAND2_X1 U813 ( .A1(G953), .A2(n1143), .ZN(n1142) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(n1141) );
XNOR2_X1 U815 ( .A(n1146), .B(n1147), .ZN(n1145) );
NAND2_X1 U816 ( .A1(KEYINPUT36), .A2(n1148), .ZN(n1146) );
INV_X1 U817 ( .A(n1135), .ZN(n1129) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1135) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1150) );
XOR2_X1 U820 ( .A(n1140), .B(KEYINPUT52), .Z(n1149) );
NAND3_X1 U821 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(G69) );
OR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND3_X1 U823 ( .A1(n1155), .A2(n1154), .A3(G953), .ZN(n1152) );
NAND2_X1 U824 ( .A1(G898), .A2(G224), .ZN(n1155) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1140), .ZN(n1151) );
NAND2_X1 U826 ( .A1(n1154), .A2(n1157), .ZN(n1156) );
OR2_X1 U827 ( .A1(n1158), .A2(n1109), .ZN(n1157) );
NAND3_X1 U828 ( .A1(n1159), .A2(n1160), .A3(n1158), .ZN(n1154) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1158) );
XOR2_X1 U830 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U831 ( .A1(KEYINPUT40), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U832 ( .A(n1166), .B(KEYINPUT29), .ZN(n1165) );
NAND2_X1 U833 ( .A1(G953), .A2(n1167), .ZN(n1160) );
XOR2_X1 U834 ( .A(KEYINPUT51), .B(n1168), .Z(n1159) );
NOR2_X1 U835 ( .A1(n1109), .A2(G953), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(G66) );
XOR2_X1 U837 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U838 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NOR2_X1 U839 ( .A1(n1169), .A2(n1175), .ZN(G63) );
XOR2_X1 U840 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND3_X1 U841 ( .A1(n1178), .A2(n1179), .A3(G478), .ZN(n1177) );
XOR2_X1 U842 ( .A(KEYINPUT8), .B(G902), .Z(n1178) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1180), .ZN(G60) );
XNOR2_X1 U844 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U845 ( .A1(n1183), .A2(n1174), .ZN(n1182) );
INV_X1 U846 ( .A(G475), .ZN(n1183) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(G6) );
NOR2_X1 U848 ( .A1(KEYINPUT30), .A2(n1186), .ZN(n1185) );
NOR4_X1 U849 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1080), .ZN(n1184) );
INV_X1 U850 ( .A(n1078), .ZN(n1189) );
NOR2_X1 U851 ( .A1(KEYINPUT59), .A2(n1190), .ZN(n1188) );
NOR3_X1 U852 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
NOR2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1187) );
INV_X1 U854 ( .A(KEYINPUT59), .ZN(n1195) );
NOR2_X1 U855 ( .A1(n1169), .A2(n1196), .ZN(G57) );
XOR2_X1 U856 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U857 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U858 ( .A1(n1201), .A2(n1174), .ZN(n1200) );
INV_X1 U859 ( .A(G472), .ZN(n1201) );
NAND2_X1 U860 ( .A1(n1202), .A2(n1203), .ZN(n1197) );
NAND2_X1 U861 ( .A1(KEYINPUT15), .A2(n1204), .ZN(n1203) );
NAND2_X1 U862 ( .A1(KEYINPUT61), .A2(n1205), .ZN(n1202) );
INV_X1 U863 ( .A(n1204), .ZN(n1205) );
XOR2_X1 U864 ( .A(n1206), .B(G101), .Z(n1204) );
NAND2_X1 U865 ( .A1(KEYINPUT12), .A2(n1207), .ZN(n1206) );
INV_X1 U866 ( .A(n1208), .ZN(n1207) );
NOR2_X1 U867 ( .A1(n1169), .A2(n1209), .ZN(G54) );
XOR2_X1 U868 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U869 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U870 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U871 ( .A1(n1122), .A2(n1174), .ZN(n1215) );
INV_X1 U872 ( .A(G469), .ZN(n1122) );
NOR2_X1 U873 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
XOR2_X1 U874 ( .A(n1218), .B(KEYINPUT10), .Z(n1217) );
NAND2_X1 U875 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U876 ( .A(n1221), .B(KEYINPUT16), .Z(n1219) );
NOR2_X1 U877 ( .A1(n1220), .A2(n1222), .ZN(n1216) );
NOR2_X1 U878 ( .A1(n1223), .A2(n1224), .ZN(n1212) );
XOR2_X1 U879 ( .A(n1225), .B(KEYINPUT13), .Z(n1224) );
NAND2_X1 U880 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NOR2_X1 U881 ( .A1(n1227), .A2(n1226), .ZN(n1223) );
XOR2_X1 U882 ( .A(n1228), .B(n1229), .Z(n1210) );
NOR2_X1 U883 ( .A1(n1169), .A2(n1230), .ZN(G51) );
XOR2_X1 U884 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U885 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U886 ( .A1(n1235), .A2(n1174), .ZN(n1234) );
NAND2_X1 U887 ( .A1(G902), .A2(n1179), .ZN(n1174) );
NAND2_X1 U888 ( .A1(n1069), .A2(n1109), .ZN(n1179) );
AND4_X1 U889 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1109) );
AND4_X1 U890 ( .A1(n1061), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1239) );
NAND3_X1 U891 ( .A1(n1078), .A2(n1243), .A3(n1194), .ZN(n1061) );
NAND2_X1 U892 ( .A1(n1194), .A2(n1244), .ZN(n1236) );
NAND2_X1 U893 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U894 ( .A1(n1082), .A2(n1107), .ZN(n1246) );
NAND2_X1 U895 ( .A1(n1247), .A2(n1078), .ZN(n1245) );
AND4_X1 U896 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1069) );
NOR4_X1 U897 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1251) );
NOR3_X1 U898 ( .A1(n1256), .A2(n1257), .A3(n1091), .ZN(n1255) );
XOR2_X1 U899 ( .A(KEYINPUT11), .B(n1247), .Z(n1256) );
AND2_X1 U900 ( .A1(n1258), .A2(n1259), .ZN(n1250) );
NOR2_X1 U901 ( .A1(n1260), .A2(n1261), .ZN(n1233) );
AND2_X1 U902 ( .A1(n1262), .A2(n1067), .ZN(n1169) );
INV_X1 U903 ( .A(G952), .ZN(n1067) );
XOR2_X1 U904 ( .A(KEYINPUT3), .B(G953), .Z(n1262) );
XNOR2_X1 U905 ( .A(G146), .B(n1248), .ZN(G48) );
NAND3_X1 U906 ( .A1(n1247), .A2(n1192), .A3(n1263), .ZN(n1248) );
XNOR2_X1 U907 ( .A(G143), .B(n1249), .ZN(G45) );
OR4_X1 U908 ( .A1(n1257), .A2(n1098), .A3(n1264), .A4(n1265), .ZN(n1249) );
NAND2_X1 U909 ( .A1(n1266), .A2(n1267), .ZN(G42) );
NAND2_X1 U910 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U911 ( .A(G140), .ZN(n1269) );
NAND2_X1 U912 ( .A1(n1259), .A2(n1270), .ZN(n1268) );
NAND2_X1 U913 ( .A1(KEYINPUT49), .A2(KEYINPUT27), .ZN(n1270) );
NAND3_X1 U914 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1266) );
INV_X1 U915 ( .A(KEYINPUT49), .ZN(n1273) );
NAND2_X1 U916 ( .A1(n1259), .A2(n1274), .ZN(n1272) );
INV_X1 U917 ( .A(KEYINPUT27), .ZN(n1274) );
NAND2_X1 U918 ( .A1(KEYINPUT27), .A2(n1275), .ZN(n1271) );
NAND2_X1 U919 ( .A1(G140), .A2(n1259), .ZN(n1275) );
NAND3_X1 U920 ( .A1(n1276), .A2(n1093), .A3(n1076), .ZN(n1259) );
NAND2_X1 U921 ( .A1(n1277), .A2(n1278), .ZN(G39) );
OR2_X1 U922 ( .A1(n1258), .A2(G137), .ZN(n1278) );
XOR2_X1 U923 ( .A(n1279), .B(KEYINPUT34), .Z(n1277) );
NAND2_X1 U924 ( .A1(G137), .A2(n1258), .ZN(n1279) );
NAND3_X1 U925 ( .A1(n1076), .A2(n1263), .A3(n1082), .ZN(n1258) );
XOR2_X1 U926 ( .A(G134), .B(n1254), .Z(G36) );
NOR3_X1 U927 ( .A1(n1257), .A2(n1081), .A3(n1091), .ZN(n1254) );
XOR2_X1 U928 ( .A(G131), .B(n1280), .Z(G33) );
NOR3_X1 U929 ( .A1(n1281), .A2(n1080), .A3(n1257), .ZN(n1280) );
NAND3_X1 U930 ( .A1(n1093), .A2(n1282), .A3(n1107), .ZN(n1257) );
XOR2_X1 U931 ( .A(KEYINPUT22), .B(n1076), .Z(n1281) );
INV_X1 U932 ( .A(n1091), .ZN(n1076) );
NAND2_X1 U933 ( .A1(n1101), .A2(n1283), .ZN(n1091) );
XOR2_X1 U934 ( .A(G128), .B(n1253), .Z(G30) );
AND3_X1 U935 ( .A1(n1243), .A2(n1192), .A3(n1263), .ZN(n1253) );
AND4_X1 U936 ( .A1(n1093), .A2(n1114), .A3(n1106), .A4(n1282), .ZN(n1263) );
INV_X1 U937 ( .A(n1191), .ZN(n1093) );
XOR2_X1 U938 ( .A(n1284), .B(n1285), .Z(G3) );
NAND3_X1 U939 ( .A1(n1107), .A2(n1194), .A3(n1286), .ZN(n1285) );
XNOR2_X1 U940 ( .A(n1082), .B(KEYINPUT47), .ZN(n1286) );
XOR2_X1 U941 ( .A(G125), .B(n1252), .Z(G27) );
AND3_X1 U942 ( .A1(n1276), .A2(n1192), .A3(n1077), .ZN(n1252) );
AND4_X1 U943 ( .A1(n1105), .A2(n1247), .A3(n1106), .A4(n1282), .ZN(n1276) );
NAND2_X1 U944 ( .A1(n1108), .A2(n1287), .ZN(n1282) );
NAND4_X1 U945 ( .A1(G953), .A2(G902), .A3(n1288), .A4(n1143), .ZN(n1287) );
INV_X1 U946 ( .A(G900), .ZN(n1143) );
XNOR2_X1 U947 ( .A(G122), .B(n1237), .ZN(G24) );
NAND4_X1 U948 ( .A1(n1289), .A2(n1078), .A3(n1116), .A4(n1124), .ZN(n1237) );
NOR2_X1 U949 ( .A1(n1106), .A2(n1114), .ZN(n1078) );
XNOR2_X1 U950 ( .A(G119), .B(n1242), .ZN(G21) );
NAND4_X1 U951 ( .A1(n1289), .A2(n1082), .A3(n1114), .A4(n1106), .ZN(n1242) );
INV_X1 U952 ( .A(n1105), .ZN(n1114) );
XOR2_X1 U953 ( .A(n1290), .B(n1241), .Z(G18) );
NAND3_X1 U954 ( .A1(n1107), .A2(n1243), .A3(n1289), .ZN(n1241) );
AND3_X1 U955 ( .A1(n1192), .A2(n1291), .A3(n1077), .ZN(n1289) );
INV_X1 U956 ( .A(n1081), .ZN(n1243) );
NAND2_X1 U957 ( .A1(n1265), .A2(n1116), .ZN(n1081) );
XOR2_X1 U958 ( .A(n1292), .B(G113), .Z(G15) );
NAND2_X1 U959 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR2_X1 U960 ( .A1(n1238), .A2(KEYINPUT54), .ZN(n1294) );
OR2_X1 U961 ( .A1(n1295), .A2(n1098), .ZN(n1238) );
NAND3_X1 U962 ( .A1(n1192), .A2(n1295), .A3(KEYINPUT54), .ZN(n1293) );
NAND4_X1 U963 ( .A1(n1107), .A2(n1077), .A3(n1247), .A4(n1291), .ZN(n1295) );
INV_X1 U964 ( .A(n1080), .ZN(n1247) );
NAND2_X1 U965 ( .A1(n1264), .A2(n1124), .ZN(n1080) );
NOR2_X1 U966 ( .A1(n1089), .A2(n1118), .ZN(n1077) );
INV_X1 U967 ( .A(n1090), .ZN(n1118) );
NOR2_X1 U968 ( .A1(n1106), .A2(n1105), .ZN(n1107) );
XOR2_X1 U969 ( .A(n1240), .B(n1296), .Z(G12) );
NAND2_X1 U970 ( .A1(KEYINPUT56), .A2(n1297), .ZN(n1296) );
XOR2_X1 U971 ( .A(KEYINPUT55), .B(G110), .Z(n1297) );
NAND4_X1 U972 ( .A1(n1082), .A2(n1194), .A3(n1105), .A4(n1106), .ZN(n1240) );
XOR2_X1 U973 ( .A(n1115), .B(KEYINPUT37), .Z(n1106) );
XOR2_X1 U974 ( .A(n1298), .B(n1173), .Z(n1115) );
NAND2_X1 U975 ( .A1(G217), .A2(n1299), .ZN(n1173) );
OR2_X1 U976 ( .A1(n1172), .A2(G902), .ZN(n1298) );
XNOR2_X1 U977 ( .A(n1300), .B(n1301), .ZN(n1172) );
XOR2_X1 U978 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U979 ( .A(G128), .B(G110), .Z(n1303) );
XOR2_X1 U980 ( .A(KEYINPUT1), .B(G137), .Z(n1302) );
XOR2_X1 U981 ( .A(n1304), .B(n1305), .Z(n1300) );
XOR2_X1 U982 ( .A(n1306), .B(n1307), .Z(n1305) );
NAND2_X1 U983 ( .A1(KEYINPUT25), .A2(n1308), .ZN(n1306) );
NAND2_X1 U984 ( .A1(n1309), .A2(G221), .ZN(n1308) );
NAND2_X1 U985 ( .A1(n1310), .A2(n1311), .ZN(n1304) );
NAND3_X1 U986 ( .A1(G146), .A2(n1147), .A3(n1312), .ZN(n1311) );
OR2_X1 U987 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
INV_X1 U988 ( .A(KEYINPUT35), .ZN(n1312) );
XOR2_X1 U989 ( .A(n1314), .B(G472), .Z(n1105) );
NAND2_X1 U990 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U991 ( .A(n1199), .B(n1317), .Z(n1315) );
XOR2_X1 U992 ( .A(n1284), .B(n1208), .Z(n1317) );
NAND3_X1 U993 ( .A1(n1318), .A2(n1140), .A3(G210), .ZN(n1208) );
XOR2_X1 U994 ( .A(KEYINPUT21), .B(G237), .Z(n1318) );
XOR2_X1 U995 ( .A(n1319), .B(n1320), .Z(n1199) );
XOR2_X1 U996 ( .A(KEYINPUT58), .B(KEYINPUT28), .Z(n1320) );
XNOR2_X1 U997 ( .A(n1321), .B(n1322), .ZN(n1319) );
NOR2_X1 U998 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NOR2_X1 U999 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NOR2_X1 U1000 ( .A1(n1327), .A2(n1328), .ZN(n1325) );
INV_X1 U1001 ( .A(KEYINPUT6), .ZN(n1328) );
NOR2_X1 U1002 ( .A1(KEYINPUT39), .A2(n1329), .ZN(n1327) );
NOR2_X1 U1003 ( .A1(G113), .A2(n1330), .ZN(n1323) );
NOR2_X1 U1004 ( .A1(n1331), .A2(KEYINPUT39), .ZN(n1330) );
AND2_X1 U1005 ( .A1(n1326), .A2(KEYINPUT6), .ZN(n1331) );
XNOR2_X1 U1006 ( .A(n1332), .B(n1333), .ZN(n1326) );
NOR2_X1 U1007 ( .A1(KEYINPUT0), .A2(n1307), .ZN(n1333) );
XOR2_X1 U1008 ( .A(n1290), .B(KEYINPUT14), .Z(n1332) );
NOR3_X1 U1009 ( .A1(n1191), .A2(n1193), .A3(n1098), .ZN(n1194) );
INV_X1 U1010 ( .A(n1192), .ZN(n1098) );
NOR2_X1 U1011 ( .A1(n1101), .A2(n1100), .ZN(n1192) );
INV_X1 U1012 ( .A(n1283), .ZN(n1100) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1334), .ZN(n1283) );
XNOR2_X1 U1014 ( .A(n1335), .B(n1235), .ZN(n1101) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1334), .ZN(n1235) );
NAND2_X1 U1016 ( .A1(n1336), .A2(n1316), .ZN(n1334) );
NAND2_X1 U1017 ( .A1(n1337), .A2(n1316), .ZN(n1335) );
XNOR2_X1 U1018 ( .A(n1231), .B(n1338), .ZN(n1337) );
NOR2_X1 U1019 ( .A1(n1261), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U1020 ( .A(n1260), .B(KEYINPUT60), .ZN(n1339) );
AND3_X1 U1021 ( .A1(n1340), .A2(n1140), .A3(G224), .ZN(n1260) );
NOR2_X1 U1022 ( .A1(n1340), .A2(n1341), .ZN(n1261) );
AND2_X1 U1023 ( .A1(G224), .A2(n1140), .ZN(n1341) );
XNOR2_X1 U1024 ( .A(n1342), .B(n1222), .ZN(n1340) );
INV_X1 U1025 ( .A(n1221), .ZN(n1222) );
XNOR2_X1 U1026 ( .A(G125), .B(KEYINPUT28), .ZN(n1342) );
XOR2_X1 U1027 ( .A(n1164), .B(n1343), .Z(n1231) );
XNOR2_X1 U1028 ( .A(n1344), .B(n1345), .ZN(n1343) );
NOR2_X1 U1029 ( .A1(KEYINPUT63), .A2(n1161), .ZN(n1345) );
XNOR2_X1 U1030 ( .A(G110), .B(n1346), .ZN(n1161) );
XOR2_X1 U1031 ( .A(KEYINPUT9), .B(G122), .Z(n1346) );
NAND2_X1 U1032 ( .A1(KEYINPUT24), .A2(n1166), .ZN(n1344) );
XNOR2_X1 U1033 ( .A(n1347), .B(KEYINPUT19), .ZN(n1166) );
NAND4_X1 U1034 ( .A1(n1348), .A2(n1349), .A3(n1350), .A4(n1351), .ZN(n1347) );
NAND3_X1 U1035 ( .A1(G101), .A2(n1352), .A3(n1186), .ZN(n1351) );
NAND3_X1 U1036 ( .A1(n1353), .A2(n1284), .A3(G104), .ZN(n1350) );
NAND2_X1 U1037 ( .A1(KEYINPUT32), .A2(n1060), .ZN(n1353) );
OR2_X1 U1038 ( .A1(n1354), .A2(n1352), .ZN(n1348) );
INV_X1 U1039 ( .A(KEYINPUT32), .ZN(n1352) );
XNOR2_X1 U1040 ( .A(n1355), .B(G113), .ZN(n1164) );
NAND2_X1 U1041 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1042 ( .A1(G116), .A2(n1307), .ZN(n1357) );
XOR2_X1 U1043 ( .A(KEYINPUT31), .B(n1358), .Z(n1356) );
NOR2_X1 U1044 ( .A1(G116), .A2(n1307), .ZN(n1358) );
XNOR2_X1 U1045 ( .A(G119), .B(KEYINPUT33), .ZN(n1307) );
INV_X1 U1046 ( .A(n1291), .ZN(n1193) );
NAND2_X1 U1047 ( .A1(n1108), .A2(n1359), .ZN(n1291) );
NAND4_X1 U1048 ( .A1(G953), .A2(G902), .A3(n1288), .A4(n1167), .ZN(n1359) );
INV_X1 U1049 ( .A(G898), .ZN(n1167) );
NAND3_X1 U1050 ( .A1(n1066), .A2(n1288), .A3(G952), .ZN(n1108) );
NAND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1288) );
XNOR2_X1 U1052 ( .A(G953), .B(KEYINPUT18), .ZN(n1066) );
NAND2_X1 U1053 ( .A1(n1089), .A2(n1090), .ZN(n1191) );
NAND2_X1 U1054 ( .A1(G221), .A2(n1299), .ZN(n1090) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1316), .ZN(n1299) );
XNOR2_X1 U1056 ( .A(n1121), .B(G469), .ZN(n1089) );
NAND2_X1 U1057 ( .A1(n1360), .A2(n1316), .ZN(n1121) );
XOR2_X1 U1058 ( .A(n1321), .B(n1361), .Z(n1360) );
XNOR2_X1 U1059 ( .A(n1220), .B(n1362), .ZN(n1361) );
NAND2_X1 U1060 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1061 ( .A1(n1227), .A2(n1365), .ZN(n1364) );
NAND2_X1 U1062 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NAND2_X1 U1063 ( .A1(KEYINPUT46), .A2(KEYINPUT26), .ZN(n1367) );
INV_X1 U1064 ( .A(n1368), .ZN(n1227) );
NAND3_X1 U1065 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1363) );
INV_X1 U1066 ( .A(KEYINPUT46), .ZN(n1371) );
NAND2_X1 U1067 ( .A1(KEYINPUT26), .A2(n1372), .ZN(n1370) );
NAND2_X1 U1068 ( .A1(n1366), .A2(n1368), .ZN(n1372) );
NAND2_X1 U1069 ( .A1(G227), .A2(n1140), .ZN(n1368) );
INV_X1 U1070 ( .A(n1226), .ZN(n1366) );
OR2_X1 U1071 ( .A1(n1226), .A2(KEYINPUT26), .ZN(n1369) );
XNOR2_X1 U1072 ( .A(G110), .B(n1373), .ZN(n1226) );
XOR2_X1 U1073 ( .A(KEYINPUT5), .B(G140), .Z(n1373) );
AND3_X1 U1074 ( .A1(n1354), .A2(n1349), .A3(n1374), .ZN(n1220) );
NAND3_X1 U1075 ( .A1(G107), .A2(n1284), .A3(G104), .ZN(n1374) );
INV_X1 U1076 ( .A(G101), .ZN(n1284) );
NAND3_X1 U1077 ( .A1(G101), .A2(n1186), .A3(G107), .ZN(n1349) );
NAND2_X1 U1078 ( .A1(n1375), .A2(n1060), .ZN(n1354) );
INV_X1 U1079 ( .A(G107), .ZN(n1060) );
XOR2_X1 U1080 ( .A(n1186), .B(G101), .Z(n1375) );
INV_X1 U1081 ( .A(G104), .ZN(n1186) );
XOR2_X1 U1082 ( .A(n1229), .B(n1144), .Z(n1321) );
XOR2_X1 U1083 ( .A(n1228), .B(n1221), .Z(n1144) );
XNOR2_X1 U1084 ( .A(G146), .B(n1376), .ZN(n1221) );
XNOR2_X1 U1085 ( .A(G134), .B(G137), .ZN(n1228) );
XNOR2_X1 U1086 ( .A(n1148), .B(KEYINPUT50), .ZN(n1229) );
INV_X1 U1087 ( .A(G131), .ZN(n1148) );
NOR2_X1 U1088 ( .A1(n1116), .A2(n1124), .ZN(n1082) );
INV_X1 U1089 ( .A(n1265), .ZN(n1124) );
XOR2_X1 U1090 ( .A(n1377), .B(G475), .Z(n1265) );
NAND2_X1 U1091 ( .A1(n1181), .A2(n1316), .ZN(n1377) );
XNOR2_X1 U1092 ( .A(n1378), .B(n1379), .ZN(n1181) );
XOR2_X1 U1093 ( .A(G104), .B(n1380), .Z(n1379) );
NOR2_X1 U1094 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
XOR2_X1 U1095 ( .A(n1383), .B(KEYINPUT23), .Z(n1382) );
NAND2_X1 U1096 ( .A1(n1384), .A2(n1313), .ZN(n1383) );
XOR2_X1 U1097 ( .A(n1385), .B(KEYINPUT53), .Z(n1384) );
NOR2_X1 U1098 ( .A1(n1313), .A2(n1385), .ZN(n1381) );
XOR2_X1 U1099 ( .A(n1386), .B(n1387), .Z(n1385) );
XOR2_X1 U1100 ( .A(G143), .B(G131), .Z(n1387) );
NAND3_X1 U1101 ( .A1(n1336), .A2(n1140), .A3(G214), .ZN(n1386) );
INV_X1 U1102 ( .A(G237), .ZN(n1336) );
XNOR2_X1 U1103 ( .A(G146), .B(n1147), .ZN(n1313) );
XOR2_X1 U1104 ( .A(G125), .B(G140), .Z(n1147) );
XOR2_X1 U1105 ( .A(n1329), .B(G122), .Z(n1378) );
INV_X1 U1106 ( .A(G113), .ZN(n1329) );
INV_X1 U1107 ( .A(n1264), .ZN(n1116) );
XOR2_X1 U1108 ( .A(n1388), .B(G478), .Z(n1264) );
NAND2_X1 U1109 ( .A1(n1316), .A2(n1176), .ZN(n1388) );
NAND2_X1 U1110 ( .A1(n1389), .A2(n1390), .ZN(n1176) );
NAND3_X1 U1111 ( .A1(G217), .A2(n1391), .A3(n1309), .ZN(n1390) );
INV_X1 U1112 ( .A(n1392), .ZN(n1391) );
XOR2_X1 U1113 ( .A(n1393), .B(KEYINPUT48), .Z(n1389) );
NAND2_X1 U1114 ( .A1(n1392), .A2(n1394), .ZN(n1393) );
NAND2_X1 U1115 ( .A1(n1309), .A2(G217), .ZN(n1394) );
AND2_X1 U1116 ( .A1(G234), .A2(n1140), .ZN(n1309) );
INV_X1 U1117 ( .A(G953), .ZN(n1140) );
XOR2_X1 U1118 ( .A(n1395), .B(n1396), .Z(n1392) );
XOR2_X1 U1119 ( .A(G107), .B(n1397), .Z(n1396) );
XOR2_X1 U1120 ( .A(G134), .B(G122), .Z(n1397) );
XOR2_X1 U1121 ( .A(n1398), .B(n1376), .Z(n1395) );
XOR2_X1 U1122 ( .A(G128), .B(G143), .Z(n1376) );
NAND2_X1 U1123 ( .A1(KEYINPUT2), .A2(n1290), .ZN(n1398) );
INV_X1 U1124 ( .A(G116), .ZN(n1290) );
INV_X1 U1125 ( .A(G902), .ZN(n1316) );
endmodule


