//Key = 0111001010010100011010010010001101000010010001001111100010001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286;

XOR2_X1 U710 ( .A(G107), .B(n978), .Z(G9) );
NOR4_X1 U711 ( .A1(n979), .A2(n980), .A3(KEYINPUT9), .A4(n981), .ZN(n978) );
NOR2_X1 U712 ( .A1(KEYINPUT26), .A2(n982), .ZN(n980) );
NOR3_X1 U713 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
AND2_X1 U714 ( .A1(n986), .A2(KEYINPUT26), .ZN(n979) );
NOR2_X1 U715 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U716 ( .A1(n989), .A2(n990), .A3(n991), .A4(n992), .ZN(n988) );
NOR2_X1 U717 ( .A1(n983), .A2(n993), .ZN(n992) );
NOR3_X1 U718 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n991) );
NOR2_X1 U719 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U720 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NOR2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1001) );
XNOR2_X1 U725 ( .A(n1009), .B(KEYINPUT37), .ZN(n1007) );
NOR2_X1 U726 ( .A1(n1010), .A2(n1004), .ZN(n997) );
NOR2_X1 U727 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U728 ( .A1(n1008), .A2(n1013), .ZN(n1011) );
NAND4_X1 U729 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n989) );
NAND4_X1 U730 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1015) );
NOR3_X1 U731 ( .A1(n1022), .A2(n996), .A3(n1023), .ZN(n1021) );
XNOR2_X1 U732 ( .A(KEYINPUT60), .B(n994), .ZN(n1022) );
XOR2_X1 U733 ( .A(KEYINPUT25), .B(n1024), .Z(n1019) );
NAND3_X1 U734 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1014) );
XOR2_X1 U735 ( .A(n993), .B(KEYINPUT38), .Z(n1027) );
OR4_X1 U736 ( .A1(n994), .A2(n1004), .A3(n1000), .A4(n1008), .ZN(n993) );
NAND2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n994) );
INV_X1 U738 ( .A(KEYINPUT4), .ZN(n1029) );
AND3_X1 U739 ( .A1(n1016), .A2(n1017), .A3(n1030), .ZN(n987) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1016) );
NOR4_X1 U741 ( .A1(n1026), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1032) );
XNOR2_X1 U742 ( .A(n1036), .B(n1037), .ZN(n1034) );
NOR2_X1 U743 ( .A1(G475), .A2(KEYINPUT44), .ZN(n1037) );
NOR4_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1031) );
XNOR2_X1 U745 ( .A(n1042), .B(n1043), .ZN(n1041) );
XNOR2_X1 U746 ( .A(G469), .B(KEYINPUT59), .ZN(n1043) );
XOR2_X1 U747 ( .A(n1044), .B(n1045), .Z(n1040) );
XNOR2_X1 U748 ( .A(KEYINPUT62), .B(n1046), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1047), .A2(KEYINPUT12), .ZN(n1044) );
INV_X1 U750 ( .A(n1048), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(G72) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1054), .A3(G953), .ZN(n1052) );
NAND3_X1 U754 ( .A1(n1055), .A2(n1054), .A3(n1056), .ZN(n1049) );
INV_X1 U755 ( .A(n1051), .ZN(n1056) );
XNOR2_X1 U756 ( .A(n1057), .B(n1058), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1059), .A2(G953), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
XOR2_X1 U759 ( .A(n1062), .B(n1063), .Z(n1060) );
XOR2_X1 U760 ( .A(n1064), .B(n1065), .Z(n1063) );
XNOR2_X1 U761 ( .A(n1066), .B(n1067), .ZN(n1064) );
XOR2_X1 U762 ( .A(n1068), .B(n1069), .Z(n1062) );
XOR2_X1 U763 ( .A(KEYINPUT27), .B(G134), .Z(n1069) );
NAND2_X1 U764 ( .A1(KEYINPUT6), .A2(G137), .ZN(n1068) );
INV_X1 U765 ( .A(KEYINPUT28), .ZN(n1054) );
NAND2_X1 U766 ( .A1(n1061), .A2(n1070), .ZN(n1055) );
NAND2_X1 U767 ( .A1(G953), .A2(n1053), .ZN(n1070) );
INV_X1 U768 ( .A(n1071), .ZN(n1061) );
XOR2_X1 U769 ( .A(n1072), .B(n1073), .Z(G69) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1017), .ZN(n1073) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1017), .ZN(n1078) );
XNOR2_X1 U774 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U776 ( .A1(G898), .A2(n1080), .A3(G953), .ZN(n1077) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(G66) );
XOR2_X1 U778 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U779 ( .A1(n1048), .A2(n1088), .ZN(n1087) );
NAND2_X1 U780 ( .A1(KEYINPUT63), .A2(n1089), .ZN(n1086) );
NOR2_X1 U781 ( .A1(n1084), .A2(n1090), .ZN(G63) );
XOR2_X1 U782 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U783 ( .A(n1093), .B(KEYINPUT23), .Z(n1091) );
NAND2_X1 U784 ( .A1(n1094), .A2(G478), .ZN(n1093) );
NOR2_X1 U785 ( .A1(n1084), .A2(n1095), .ZN(G60) );
NOR3_X1 U786 ( .A1(n1036), .A2(n1096), .A3(n1097), .ZN(n1095) );
AND3_X1 U787 ( .A1(n1098), .A2(G475), .A3(n1094), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1098), .ZN(n1096) );
AND2_X1 U789 ( .A1(n990), .A2(G475), .ZN(n1099) );
XNOR2_X1 U790 ( .A(G104), .B(n1100), .ZN(G6) );
NOR2_X1 U791 ( .A1(n1084), .A2(n1101), .ZN(G57) );
XOR2_X1 U792 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U793 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U794 ( .A(n1106), .B(n1107), .ZN(n1102) );
XOR2_X1 U795 ( .A(n1108), .B(n1109), .Z(n1107) );
AND2_X1 U796 ( .A1(G472), .A2(n1094), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1084), .A2(n1110), .ZN(G54) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U799 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U800 ( .A1(n1115), .A2(KEYINPUT56), .ZN(n1113) );
XNOR2_X1 U801 ( .A(n1116), .B(n1117), .ZN(n1115) );
XNOR2_X1 U802 ( .A(KEYINPUT20), .B(n1118), .ZN(n1117) );
XOR2_X1 U803 ( .A(n1119), .B(n1120), .Z(n1111) );
NOR3_X1 U804 ( .A1(n1088), .A2(KEYINPUT29), .A3(n1121), .ZN(n1120) );
INV_X1 U805 ( .A(G469), .ZN(n1121) );
XNOR2_X1 U806 ( .A(KEYINPUT8), .B(n1122), .ZN(n1119) );
NOR2_X1 U807 ( .A1(KEYINPUT57), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U808 ( .A(G110), .B(n1124), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1084), .A2(n1125), .ZN(G51) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U811 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1128) );
XOR2_X1 U814 ( .A(KEYINPUT50), .B(n1131), .Z(n1132) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(n1126) );
NOR2_X1 U816 ( .A1(KEYINPUT15), .A2(n1136), .ZN(n1135) );
INV_X1 U817 ( .A(n1080), .ZN(n1136) );
NAND2_X1 U818 ( .A1(n1094), .A2(n1137), .ZN(n1134) );
INV_X1 U819 ( .A(n1088), .ZN(n1094) );
NAND2_X1 U820 ( .A1(G902), .A2(n990), .ZN(n1088) );
NAND3_X1 U821 ( .A1(n1059), .A2(n1138), .A3(n1139), .ZN(n990) );
INV_X1 U822 ( .A(n1083), .ZN(n1139) );
NAND4_X1 U823 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1083) );
AND4_X1 U824 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
NAND2_X1 U825 ( .A1(n1012), .A2(n1148), .ZN(n1147) );
INV_X1 U826 ( .A(n981), .ZN(n1012) );
NAND2_X1 U827 ( .A1(n1018), .A2(n1149), .ZN(n981) );
INV_X1 U828 ( .A(n1008), .ZN(n1018) );
NAND2_X1 U829 ( .A1(n1150), .A2(n1151), .ZN(n1142) );
XOR2_X1 U830 ( .A(n1152), .B(KEYINPUT31), .Z(n1150) );
NAND2_X1 U831 ( .A1(KEYINPUT11), .A2(n1153), .ZN(n1141) );
NAND3_X1 U832 ( .A1(n1154), .A2(n985), .A3(n1006), .ZN(n1140) );
NAND2_X1 U833 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
INV_X1 U834 ( .A(n1157), .ZN(n1156) );
OR4_X1 U835 ( .A1(n1000), .A2(n984), .A3(n1151), .A4(KEYINPUT11), .ZN(n1155) );
INV_X1 U836 ( .A(n1158), .ZN(n984) );
XNOR2_X1 U837 ( .A(KEYINPUT41), .B(n1100), .ZN(n1138) );
INV_X1 U838 ( .A(n1082), .ZN(n1100) );
NOR3_X1 U839 ( .A1(n986), .A2(n1008), .A3(n1013), .ZN(n1082) );
AND4_X1 U840 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1059) );
NOR4_X1 U841 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NOR3_X1 U842 ( .A1(n1167), .A2(n1168), .A3(n983), .ZN(n1166) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1170), .ZN(n1161) );
AND2_X1 U844 ( .A1(n1171), .A2(n1030), .ZN(n1084) );
INV_X1 U845 ( .A(G952), .ZN(n1030) );
XNOR2_X1 U846 ( .A(G953), .B(KEYINPUT52), .ZN(n1171) );
XNOR2_X1 U847 ( .A(n1172), .B(n1165), .ZN(G48) );
AND2_X1 U848 ( .A1(n1173), .A2(n1174), .ZN(n1165) );
XOR2_X1 U849 ( .A(G143), .B(n1175), .Z(G45) );
NOR3_X1 U850 ( .A1(n1167), .A2(n1168), .A3(n1176), .ZN(n1175) );
XNOR2_X1 U851 ( .A(n1151), .B(KEYINPUT55), .ZN(n1176) );
XOR2_X1 U852 ( .A(G140), .B(n1169), .Z(G42) );
AND3_X1 U853 ( .A1(n1173), .A2(n1005), .A3(n1177), .ZN(n1169) );
XOR2_X1 U854 ( .A(G137), .B(n1164), .Z(G39) );
AND3_X1 U855 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1164) );
NOR3_X1 U856 ( .A1(n1000), .A2(n1180), .A3(n1181), .ZN(n1179) );
INV_X1 U857 ( .A(n1020), .ZN(n1000) );
XOR2_X1 U858 ( .A(G134), .B(n1163), .Z(G36) );
NOR3_X1 U859 ( .A1(n1182), .A2(n996), .A3(n1167), .ZN(n1163) );
NAND3_X1 U860 ( .A1(n1006), .A2(n1039), .A3(n1178), .ZN(n1167) );
XNOR2_X1 U861 ( .A(G131), .B(n1159), .ZN(G33) );
NAND3_X1 U862 ( .A1(n1173), .A2(n1006), .A3(n1177), .ZN(n1159) );
INV_X1 U863 ( .A(n996), .ZN(n1177) );
NAND2_X1 U864 ( .A1(n1025), .A2(n1183), .ZN(n996) );
XNOR2_X1 U865 ( .A(n1038), .B(KEYINPUT16), .ZN(n1025) );
AND2_X1 U866 ( .A1(n1178), .A2(n1184), .ZN(n1173) );
AND2_X1 U867 ( .A1(n1009), .A2(n1185), .ZN(n1178) );
XNOR2_X1 U868 ( .A(G128), .B(n1160), .ZN(G30) );
NAND4_X1 U869 ( .A1(n1174), .A2(n1149), .A3(n1158), .A4(n1185), .ZN(n1160) );
XOR2_X1 U870 ( .A(n1153), .B(n1186), .Z(G3) );
NOR2_X1 U871 ( .A1(KEYINPUT34), .A2(n1187), .ZN(n1186) );
AND3_X1 U872 ( .A1(n1148), .A2(n1020), .A3(n1006), .ZN(n1153) );
XNOR2_X1 U873 ( .A(G125), .B(n1188), .ZN(G27) );
NOR2_X1 U874 ( .A1(n1170), .A2(KEYINPUT36), .ZN(n1188) );
AND3_X1 U875 ( .A1(n1005), .A2(n1185), .A3(n1157), .ZN(n1170) );
NOR3_X1 U876 ( .A1(n1004), .A2(n983), .A3(n1013), .ZN(n1157) );
INV_X1 U877 ( .A(n1184), .ZN(n1013) );
NAND2_X1 U878 ( .A1(n1189), .A2(n1190), .ZN(n1185) );
NAND3_X1 U879 ( .A1(G902), .A2(n1028), .A3(n1071), .ZN(n1190) );
NOR2_X1 U880 ( .A1(G900), .A2(n1017), .ZN(n1071) );
XOR2_X1 U881 ( .A(n1191), .B(n1192), .Z(G24) );
NOR2_X1 U882 ( .A1(KEYINPUT46), .A2(n1193), .ZN(n1192) );
NOR2_X1 U883 ( .A1(n983), .A2(n1152), .ZN(n1191) );
NAND4_X1 U884 ( .A1(n1182), .A2(n985), .A3(n1039), .A4(n1194), .ZN(n1152) );
NOR2_X1 U885 ( .A1(n1008), .A2(n1004), .ZN(n1194) );
NAND2_X1 U886 ( .A1(n1180), .A2(n1195), .ZN(n1008) );
XNOR2_X1 U887 ( .A(G119), .B(n1146), .ZN(G21) );
NAND4_X1 U888 ( .A1(n1174), .A2(n1196), .A3(n1020), .A4(n985), .ZN(n1146) );
NOR3_X1 U889 ( .A1(n1181), .A2(n1180), .A3(n983), .ZN(n1174) );
INV_X1 U890 ( .A(n1151), .ZN(n983) );
NAND2_X1 U891 ( .A1(n1197), .A2(n1198), .ZN(G18) );
NAND2_X1 U892 ( .A1(G116), .A2(n1145), .ZN(n1198) );
XOR2_X1 U893 ( .A(KEYINPUT2), .B(n1199), .Z(n1197) );
NOR2_X1 U894 ( .A1(G116), .A2(n1145), .ZN(n1199) );
NAND3_X1 U895 ( .A1(n1200), .A2(n1149), .A3(n1196), .ZN(n1145) );
NOR2_X1 U896 ( .A1(n1182), .A2(n1201), .ZN(n1149) );
INV_X1 U897 ( .A(n1039), .ZN(n1201) );
XNOR2_X1 U898 ( .A(G113), .B(n1202), .ZN(G15) );
NAND3_X1 U899 ( .A1(n1184), .A2(n1200), .A3(n1203), .ZN(n1202) );
XNOR2_X1 U900 ( .A(n1196), .B(KEYINPUT49), .ZN(n1203) );
INV_X1 U901 ( .A(n1004), .ZN(n1196) );
NAND2_X1 U902 ( .A1(n1024), .A2(n1023), .ZN(n1004) );
AND3_X1 U903 ( .A1(n1151), .A2(n985), .A3(n1006), .ZN(n1200) );
AND2_X1 U904 ( .A1(n1195), .A2(n1035), .ZN(n1006) );
NOR2_X1 U905 ( .A1(n1039), .A2(n1168), .ZN(n1184) );
XNOR2_X1 U906 ( .A(G110), .B(n1144), .ZN(G12) );
NAND3_X1 U907 ( .A1(n1020), .A2(n1005), .A3(n1148), .ZN(n1144) );
INV_X1 U908 ( .A(n986), .ZN(n1148) );
NAND3_X1 U909 ( .A1(n1158), .A2(n985), .A3(n1151), .ZN(n986) );
NOR2_X1 U910 ( .A1(n1204), .A2(n1026), .ZN(n1151) );
INV_X1 U911 ( .A(n1183), .ZN(n1026) );
NAND2_X1 U912 ( .A1(G214), .A2(n1205), .ZN(n1183) );
INV_X1 U913 ( .A(n1038), .ZN(n1204) );
XNOR2_X1 U914 ( .A(n1206), .B(n1137), .ZN(n1038) );
AND2_X1 U915 ( .A1(G210), .A2(n1205), .ZN(n1137) );
NAND2_X1 U916 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U917 ( .A(G237), .ZN(n1207) );
NAND2_X1 U918 ( .A1(n1209), .A2(n1208), .ZN(n1206) );
XOR2_X1 U919 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U920 ( .A(KEYINPUT53), .B(n1130), .ZN(n1211) );
XNOR2_X1 U921 ( .A(n1080), .B(n1131), .ZN(n1210) );
XOR2_X1 U922 ( .A(G125), .B(n1212), .Z(n1131) );
NOR2_X1 U923 ( .A1(G953), .A2(n1075), .ZN(n1212) );
INV_X1 U924 ( .A(G224), .ZN(n1075) );
XNOR2_X1 U925 ( .A(n1213), .B(n1214), .ZN(n1080) );
XNOR2_X1 U926 ( .A(n1193), .B(n1215), .ZN(n1214) );
NOR2_X1 U927 ( .A1(KEYINPUT5), .A2(n1118), .ZN(n1215) );
XNOR2_X1 U928 ( .A(n1216), .B(n1106), .ZN(n1213) );
NAND2_X1 U929 ( .A1(n1189), .A2(n1217), .ZN(n985) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1028), .A4(n1076), .ZN(n1217) );
INV_X1 U931 ( .A(G898), .ZN(n1076) );
NAND3_X1 U932 ( .A1(n1028), .A2(n1017), .A3(G952), .ZN(n1189) );
NAND2_X1 U933 ( .A1(n1218), .A2(G234), .ZN(n1028) );
XNOR2_X1 U934 ( .A(G237), .B(KEYINPUT13), .ZN(n1218) );
XOR2_X1 U935 ( .A(n1009), .B(KEYINPUT14), .Z(n1158) );
NOR2_X1 U936 ( .A1(n1024), .A2(n1033), .ZN(n1009) );
INV_X1 U937 ( .A(n1023), .ZN(n1033) );
NAND2_X1 U938 ( .A1(G221), .A2(n1219), .ZN(n1023) );
XNOR2_X1 U939 ( .A(n1220), .B(n1221), .ZN(n1024) );
NOR2_X1 U940 ( .A1(KEYINPUT39), .A2(n1042), .ZN(n1221) );
AND2_X1 U941 ( .A1(n1222), .A2(n1208), .ZN(n1042) );
XOR2_X1 U942 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U943 ( .A(n1124), .B(n1216), .ZN(n1224) );
XOR2_X1 U944 ( .A(G110), .B(n1116), .Z(n1216) );
XOR2_X1 U945 ( .A(G104), .B(G107), .Z(n1116) );
XNOR2_X1 U946 ( .A(G140), .B(n1225), .ZN(n1124) );
NOR2_X1 U947 ( .A1(G953), .A2(n1053), .ZN(n1225) );
INV_X1 U948 ( .A(G227), .ZN(n1053) );
XOR2_X1 U949 ( .A(n1118), .B(n1114), .Z(n1223) );
XOR2_X1 U950 ( .A(n1067), .B(n1109), .Z(n1114) );
XOR2_X1 U951 ( .A(n1226), .B(n1066), .Z(n1109) );
XNOR2_X1 U952 ( .A(G128), .B(n1227), .ZN(n1066) );
XOR2_X1 U953 ( .A(n1228), .B(KEYINPUT10), .Z(n1067) );
XNOR2_X1 U954 ( .A(G101), .B(KEYINPUT17), .ZN(n1118) );
XNOR2_X1 U955 ( .A(G469), .B(KEYINPUT0), .ZN(n1220) );
AND2_X1 U956 ( .A1(n1229), .A2(n1180), .ZN(n1005) );
INV_X1 U957 ( .A(n1035), .ZN(n1180) );
XNOR2_X1 U958 ( .A(n1230), .B(G472), .ZN(n1035) );
NAND2_X1 U959 ( .A1(n1231), .A2(n1208), .ZN(n1230) );
XOR2_X1 U960 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U961 ( .A(n1226), .B(n1234), .Z(n1233) );
XOR2_X1 U962 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U963 ( .A1(KEYINPUT21), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U964 ( .A(KEYINPUT33), .B(n1238), .ZN(n1237) );
INV_X1 U965 ( .A(n1106), .ZN(n1238) );
XNOR2_X1 U966 ( .A(n1239), .B(n1240), .ZN(n1106) );
XOR2_X1 U967 ( .A(KEYINPUT22), .B(G119), .Z(n1240) );
XNOR2_X1 U968 ( .A(G113), .B(G116), .ZN(n1239) );
NOR2_X1 U969 ( .A1(n1133), .A2(n1241), .ZN(n1235) );
XOR2_X1 U970 ( .A(KEYINPUT54), .B(KEYINPUT42), .Z(n1241) );
INV_X1 U971 ( .A(n1130), .ZN(n1133) );
XOR2_X1 U972 ( .A(G128), .B(n1105), .Z(n1130) );
NAND2_X1 U973 ( .A1(n1242), .A2(n1243), .ZN(n1105) );
OR2_X1 U974 ( .A1(n1228), .A2(KEYINPUT43), .ZN(n1243) );
NAND3_X1 U975 ( .A1(G143), .A2(n1172), .A3(KEYINPUT43), .ZN(n1242) );
XOR2_X1 U976 ( .A(KEYINPUT7), .B(n1244), .Z(n1226) );
NOR2_X1 U977 ( .A1(KEYINPUT32), .A2(n1245), .ZN(n1244) );
XOR2_X1 U978 ( .A(G137), .B(G134), .Z(n1245) );
XNOR2_X1 U979 ( .A(n1104), .B(n1227), .ZN(n1232) );
INV_X1 U980 ( .A(n1246), .ZN(n1227) );
XNOR2_X1 U981 ( .A(n1247), .B(n1187), .ZN(n1104) );
INV_X1 U982 ( .A(G101), .ZN(n1187) );
NAND2_X1 U983 ( .A1(G210), .A2(n1248), .ZN(n1247) );
XOR2_X1 U984 ( .A(n1181), .B(KEYINPUT51), .Z(n1229) );
XOR2_X1 U985 ( .A(n1195), .B(KEYINPUT40), .Z(n1181) );
XNOR2_X1 U986 ( .A(n1046), .B(n1048), .ZN(n1195) );
NAND2_X1 U987 ( .A1(G217), .A2(n1219), .ZN(n1048) );
NAND2_X1 U988 ( .A1(G234), .A2(n1208), .ZN(n1219) );
NAND2_X1 U989 ( .A1(n1089), .A2(n1208), .ZN(n1046) );
INV_X1 U990 ( .A(G902), .ZN(n1208) );
XOR2_X1 U991 ( .A(n1249), .B(n1250), .Z(n1089) );
NOR2_X1 U992 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U993 ( .A(n1253), .B(KEYINPUT48), .Z(n1252) );
NAND2_X1 U994 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U995 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
XNOR2_X1 U996 ( .A(n1256), .B(n1065), .ZN(n1255) );
XOR2_X1 U997 ( .A(G125), .B(G140), .Z(n1065) );
XNOR2_X1 U998 ( .A(G146), .B(KEYINPUT45), .ZN(n1256) );
XOR2_X1 U999 ( .A(n1257), .B(G110), .Z(n1254) );
NAND2_X1 U1000 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
OR2_X1 U1001 ( .A1(n1260), .A2(G119), .ZN(n1259) );
XOR2_X1 U1002 ( .A(n1261), .B(KEYINPUT47), .Z(n1258) );
NAND2_X1 U1003 ( .A1(G119), .A2(n1260), .ZN(n1261) );
NAND2_X1 U1004 ( .A1(KEYINPUT1), .A2(n1262), .ZN(n1249) );
XNOR2_X1 U1005 ( .A(G137), .B(n1263), .ZN(n1262) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1264), .ZN(n1263) );
NOR2_X1 U1007 ( .A1(n1039), .A2(n1182), .ZN(n1020) );
INV_X1 U1008 ( .A(n1168), .ZN(n1182) );
XNOR2_X1 U1009 ( .A(n1036), .B(G475), .ZN(n1168) );
NOR2_X1 U1010 ( .A1(n1098), .A2(G902), .ZN(n1036) );
XNOR2_X1 U1011 ( .A(n1265), .B(n1266), .ZN(n1098) );
XOR2_X1 U1012 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U1013 ( .A(n1269), .B(n1270), .ZN(n1268) );
NOR2_X1 U1014 ( .A1(KEYINPUT58), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U1015 ( .A(n1272), .B(n1273), .ZN(n1271) );
XNOR2_X1 U1016 ( .A(n1193), .B(G113), .ZN(n1273) );
INV_X1 U1017 ( .A(G104), .ZN(n1272) );
NOR2_X1 U1018 ( .A1(KEYINPUT35), .A2(n1274), .ZN(n1269) );
XNOR2_X1 U1019 ( .A(G125), .B(KEYINPUT18), .ZN(n1274) );
XNOR2_X1 U1020 ( .A(G140), .B(KEYINPUT19), .ZN(n1267) );
XOR2_X1 U1021 ( .A(n1275), .B(n1228), .Z(n1265) );
XNOR2_X1 U1022 ( .A(G143), .B(n1172), .ZN(n1228) );
INV_X1 U1023 ( .A(G146), .ZN(n1172) );
XNOR2_X1 U1024 ( .A(n1246), .B(n1276), .ZN(n1275) );
AND2_X1 U1025 ( .A1(n1248), .A2(G214), .ZN(n1276) );
AND2_X1 U1026 ( .A1(n1277), .A2(n1017), .ZN(n1248) );
XNOR2_X1 U1027 ( .A(G237), .B(KEYINPUT24), .ZN(n1277) );
XOR2_X1 U1028 ( .A(G131), .B(KEYINPUT30), .Z(n1246) );
XNOR2_X1 U1029 ( .A(n1278), .B(G478), .ZN(n1039) );
OR2_X1 U1030 ( .A1(n1092), .A2(G902), .ZN(n1278) );
XNOR2_X1 U1031 ( .A(n1279), .B(n1280), .ZN(n1092) );
XOR2_X1 U1032 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U1033 ( .A1(n1283), .A2(KEYINPUT61), .ZN(n1282) );
XNOR2_X1 U1034 ( .A(G107), .B(n1284), .ZN(n1283) );
XNOR2_X1 U1035 ( .A(n1193), .B(G116), .ZN(n1284) );
INV_X1 U1036 ( .A(G122), .ZN(n1193) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1264), .ZN(n1281) );
AND2_X1 U1038 ( .A1(G234), .A2(n1017), .ZN(n1264) );
INV_X1 U1039 ( .A(G953), .ZN(n1017) );
XOR2_X1 U1040 ( .A(n1285), .B(G134), .Z(n1279) );
NAND2_X1 U1041 ( .A1(KEYINPUT3), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U1042 ( .A(G143), .B(n1260), .ZN(n1286) );
INV_X1 U1043 ( .A(G128), .ZN(n1260) );
endmodule


