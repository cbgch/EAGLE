//Key = 1010100010011110000100001110100000011100001011111001100011000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354;

XNOR2_X1 U743 ( .A(G107), .B(n1023), .ZN(G9) );
NOR2_X1 U744 ( .A1(n1024), .A2(n1025), .ZN(G75) );
XOR2_X1 U745 ( .A(n1026), .B(KEYINPUT2), .Z(n1025) );
NAND3_X1 U746 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NOR3_X1 U747 ( .A1(n1030), .A2(n1027), .A3(n1031), .ZN(n1024) );
INV_X1 U748 ( .A(G952), .ZN(n1027) );
NAND3_X1 U749 ( .A1(n1029), .A2(n1028), .A3(n1032), .ZN(n1030) );
NAND2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U751 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND4_X1 U752 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NAND2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1043), .ZN(n1035) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND3_X1 U757 ( .A1(n1038), .A2(n1044), .A3(n1037), .ZN(n1048) );
OR3_X1 U758 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1039), .A2(n1052), .ZN(n1047) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1038), .A2(n1055), .ZN(n1054) );
OR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1037), .A2(n1058), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U766 ( .A(n1063), .ZN(n1059) );
INV_X1 U767 ( .A(n1064), .ZN(n1033) );
NAND4_X1 U768 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1029) );
NOR4_X1 U769 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
XNOR2_X1 U770 ( .A(n1073), .B(n1074), .ZN(n1072) );
XOR2_X1 U771 ( .A(KEYINPUT8), .B(n1075), .Z(n1074) );
AND2_X1 U772 ( .A1(n1076), .A2(G478), .ZN(n1071) );
XNOR2_X1 U773 ( .A(n1077), .B(n1078), .ZN(n1070) );
NAND2_X1 U774 ( .A1(KEYINPUT13), .A2(n1079), .ZN(n1077) );
XOR2_X1 U775 ( .A(KEYINPUT44), .B(G475), .Z(n1079) );
NAND3_X1 U776 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1069) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
OR2_X1 U779 ( .A1(n1087), .A2(KEYINPUT51), .ZN(n1086) );
NAND2_X1 U780 ( .A1(KEYINPUT51), .A2(n1088), .ZN(n1085) );
INV_X1 U781 ( .A(n1089), .ZN(n1088) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1089), .ZN(n1080) );
NOR2_X1 U783 ( .A1(n1087), .A2(KEYINPUT39), .ZN(n1089) );
NOR3_X1 U784 ( .A1(n1051), .A2(n1091), .A3(n1092), .ZN(n1067) );
NAND2_X1 U785 ( .A1(G469), .A2(n1093), .ZN(n1065) );
XOR2_X1 U786 ( .A(n1094), .B(n1095), .Z(G72) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U789 ( .A(KEYINPUT30), .B(n1100), .Z(n1099) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1098) );
NAND3_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1101) );
NAND2_X1 U792 ( .A1(KEYINPUT5), .A2(n1106), .ZN(n1105) );
OR3_X1 U793 ( .A1(n1106), .A2(KEYINPUT5), .A3(n1107), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1103) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U796 ( .A(KEYINPUT5), .ZN(n1110) );
XNOR2_X1 U797 ( .A(n1106), .B(KEYINPUT21), .ZN(n1109) );
XNOR2_X1 U798 ( .A(n1111), .B(G131), .ZN(n1107) );
NOR2_X1 U799 ( .A1(G953), .A2(n1112), .ZN(n1096) );
NOR3_X1 U800 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
XOR2_X1 U801 ( .A(KEYINPUT17), .B(n1116), .Z(n1115) );
XOR2_X1 U802 ( .A(KEYINPUT38), .B(n1117), .Z(n1113) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1028), .ZN(n1094) );
AND2_X1 U804 ( .A1(G227), .A2(G900), .ZN(n1118) );
NAND2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(G69) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
OR2_X1 U807 ( .A1(n1028), .A2(G224), .ZN(n1122) );
NAND3_X1 U808 ( .A1(n1123), .A2(n1124), .A3(G953), .ZN(n1119) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1124) );
XOR2_X1 U810 ( .A(KEYINPUT56), .B(n1121), .Z(n1123) );
XNOR2_X1 U811 ( .A(n1125), .B(n1126), .ZN(n1121) );
NOR3_X1 U812 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NOR2_X1 U813 ( .A1(G898), .A2(n1028), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1028), .A2(n1132), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U817 ( .A(KEYINPUT53), .B(n1135), .Z(n1134) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1133) );
NOR2_X1 U819 ( .A1(n1138), .A2(KEYINPUT27), .ZN(n1137) );
NAND2_X1 U820 ( .A1(n1139), .A2(n1075), .ZN(n1136) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1140), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1141), .B(n1142), .ZN(n1140) );
NOR3_X1 U823 ( .A1(n1143), .A2(KEYINPUT59), .A3(n1144), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1135), .A2(n1145), .ZN(G60) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U826 ( .A(KEYINPUT19), .B(n1148), .Z(n1147) );
AND2_X1 U827 ( .A1(G475), .A2(n1139), .ZN(n1148) );
XOR2_X1 U828 ( .A(n1149), .B(n1150), .Z(G6) );
XOR2_X1 U829 ( .A(KEYINPUT28), .B(G104), .Z(n1150) );
NAND4_X1 U830 ( .A1(n1056), .A2(n1151), .A3(n1152), .A4(n1063), .ZN(n1149) );
NOR2_X1 U831 ( .A1(KEYINPUT54), .A2(n1153), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(G57) );
XOR2_X1 U833 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U834 ( .A(n1158), .B(n1159), .ZN(n1157) );
XOR2_X1 U835 ( .A(n1160), .B(n1161), .Z(n1156) );
AND2_X1 U836 ( .A1(G472), .A2(n1139), .ZN(n1160) );
NOR2_X1 U837 ( .A1(G952), .A2(n1162), .ZN(n1154) );
XNOR2_X1 U838 ( .A(KEYINPUT11), .B(n1028), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1135), .A2(n1163), .ZN(G54) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U843 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
NOR2_X1 U845 ( .A1(KEYINPUT6), .A2(n1174), .ZN(n1168) );
INV_X1 U846 ( .A(n1106), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1175), .A2(n1143), .ZN(n1166) );
XNOR2_X1 U848 ( .A(n1176), .B(n1177), .ZN(n1164) );
NOR2_X1 U849 ( .A1(n1135), .A2(n1178), .ZN(G51) );
XOR2_X1 U850 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U851 ( .A1(KEYINPUT46), .A2(n1181), .ZN(n1179) );
NAND2_X1 U852 ( .A1(n1139), .A2(n1090), .ZN(n1181) );
INV_X1 U853 ( .A(n1143), .ZN(n1139) );
NAND2_X1 U854 ( .A1(G902), .A2(n1031), .ZN(n1143) );
OR4_X1 U855 ( .A1(n1132), .A2(n1114), .A3(n1117), .A4(n1116), .ZN(n1031) );
NAND4_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1114) );
NOR3_X1 U857 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
NAND4_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1057), .ZN(n1184) );
XNOR2_X1 U859 ( .A(KEYINPUT52), .B(n1063), .ZN(n1189) );
NAND4_X1 U860 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1132) );
AND4_X1 U861 ( .A1(n1023), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1195) );
NAND4_X1 U862 ( .A1(n1151), .A2(n1057), .A3(n1063), .A4(n1039), .ZN(n1023) );
NAND3_X1 U863 ( .A1(n1039), .A2(n1199), .A3(n1151), .ZN(n1194) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND3_X1 U865 ( .A1(n1202), .A2(n1203), .A3(n1038), .ZN(n1201) );
NAND2_X1 U866 ( .A1(n1056), .A2(n1063), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1028), .A2(G952), .ZN(n1135) );
XNOR2_X1 U868 ( .A(G146), .B(n1182), .ZN(G48) );
NAND4_X1 U869 ( .A1(n1190), .A2(n1191), .A3(n1056), .A4(n1063), .ZN(n1182) );
XNOR2_X1 U870 ( .A(G143), .B(n1183), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1190), .A2(n1050), .A3(n1204), .A4(n1063), .ZN(n1183) );
NOR2_X1 U872 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XNOR2_X1 U873 ( .A(n1207), .B(n1117), .ZN(G42) );
AND3_X1 U874 ( .A1(n1208), .A2(n1049), .A3(n1056), .ZN(n1117) );
XOR2_X1 U875 ( .A(G137), .B(n1186), .Z(G39) );
AND3_X1 U876 ( .A1(n1208), .A2(n1037), .A3(n1191), .ZN(n1186) );
XOR2_X1 U877 ( .A(n1188), .B(n1209), .Z(G36) );
NOR2_X1 U878 ( .A1(KEYINPUT16), .A2(n1210), .ZN(n1209) );
AND3_X1 U879 ( .A1(n1208), .A2(n1057), .A3(n1050), .ZN(n1188) );
XOR2_X1 U880 ( .A(G131), .B(n1116), .Z(G33) );
AND3_X1 U881 ( .A1(n1050), .A2(n1208), .A3(n1056), .ZN(n1116) );
AND4_X1 U882 ( .A1(n1063), .A2(n1043), .A3(n1211), .A4(n1046), .ZN(n1208) );
XOR2_X1 U883 ( .A(n1212), .B(n1213), .Z(G30) );
NOR2_X1 U884 ( .A1(n1214), .A2(n1041), .ZN(n1213) );
INV_X1 U885 ( .A(n1215), .ZN(n1041) );
XOR2_X1 U886 ( .A(n1216), .B(KEYINPUT22), .Z(n1214) );
NAND4_X1 U887 ( .A1(n1191), .A2(n1057), .A3(n1063), .A4(n1211), .ZN(n1216) );
NOR2_X1 U888 ( .A1(KEYINPUT1), .A2(n1217), .ZN(n1212) );
XNOR2_X1 U889 ( .A(G101), .B(n1192), .ZN(G3) );
NAND2_X1 U890 ( .A1(n1218), .A2(n1050), .ZN(n1192) );
XOR2_X1 U891 ( .A(G125), .B(n1187), .Z(G27) );
AND4_X1 U892 ( .A1(n1190), .A2(n1056), .A3(n1038), .A4(n1049), .ZN(n1187) );
AND2_X1 U893 ( .A1(n1215), .A2(n1211), .ZN(n1190) );
NAND2_X1 U894 ( .A1(n1064), .A2(n1219), .ZN(n1211) );
NAND3_X1 U895 ( .A1(G902), .A2(n1220), .A3(n1100), .ZN(n1219) );
AND2_X1 U896 ( .A1(G953), .A2(n1221), .ZN(n1100) );
XOR2_X1 U897 ( .A(KEYINPUT37), .B(G900), .Z(n1221) );
XNOR2_X1 U898 ( .A(G122), .B(n1222), .ZN(G24) );
NAND3_X1 U899 ( .A1(KEYINPUT14), .A2(n1223), .A3(n1224), .ZN(n1222) );
NOR3_X1 U900 ( .A1(n1153), .A2(n1205), .A3(n1206), .ZN(n1224) );
INV_X1 U901 ( .A(n1039), .ZN(n1153) );
NAND2_X1 U902 ( .A1(n1225), .A2(n1226), .ZN(n1039) );
OR2_X1 U903 ( .A1(n1227), .A2(KEYINPUT48), .ZN(n1226) );
NAND3_X1 U904 ( .A1(n1082), .A2(n1228), .A3(KEYINPUT48), .ZN(n1225) );
XNOR2_X1 U905 ( .A(G119), .B(n1193), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1223), .A2(n1037), .A3(n1191), .ZN(n1193) );
NOR2_X1 U907 ( .A1(n1228), .A2(n1082), .ZN(n1191) );
INV_X1 U908 ( .A(n1229), .ZN(n1228) );
XNOR2_X1 U909 ( .A(G116), .B(n1198), .ZN(G18) );
NAND3_X1 U910 ( .A1(n1050), .A2(n1057), .A3(n1223), .ZN(n1198) );
NOR2_X1 U911 ( .A1(n1202), .A2(n1205), .ZN(n1057) );
INV_X1 U912 ( .A(n1203), .ZN(n1205) );
XNOR2_X1 U913 ( .A(G113), .B(n1197), .ZN(G15) );
NAND3_X1 U914 ( .A1(n1056), .A2(n1050), .A3(n1223), .ZN(n1197) );
AND2_X1 U915 ( .A1(n1151), .A2(n1038), .ZN(n1223) );
NOR2_X1 U916 ( .A1(n1229), .A2(n1082), .ZN(n1050) );
NOR2_X1 U917 ( .A1(n1203), .A2(n1206), .ZN(n1056) );
XOR2_X1 U918 ( .A(n1196), .B(n1230), .Z(G12) );
NOR2_X1 U919 ( .A1(G110), .A2(KEYINPUT20), .ZN(n1230) );
NAND2_X1 U920 ( .A1(n1218), .A2(n1049), .ZN(n1196) );
INV_X1 U921 ( .A(n1227), .ZN(n1049) );
NAND2_X1 U922 ( .A1(n1082), .A2(n1229), .ZN(n1227) );
XNOR2_X1 U923 ( .A(n1231), .B(n1075), .ZN(n1229) );
AND2_X1 U924 ( .A1(G217), .A2(n1232), .ZN(n1075) );
NAND2_X1 U925 ( .A1(KEYINPUT61), .A2(n1073), .ZN(n1231) );
NOR2_X1 U926 ( .A1(G902), .A2(n1138), .ZN(n1073) );
AND2_X1 U927 ( .A1(n1233), .A2(n1234), .ZN(n1138) );
NAND2_X1 U928 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U929 ( .A(n1237), .B(n1238), .ZN(n1235) );
XOR2_X1 U930 ( .A(n1239), .B(KEYINPUT50), .Z(n1233) );
NAND2_X1 U931 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XNOR2_X1 U932 ( .A(n1238), .B(n1242), .ZN(n1241) );
INV_X1 U933 ( .A(n1237), .ZN(n1242) );
XOR2_X1 U934 ( .A(G110), .B(n1243), .Z(n1237) );
XNOR2_X1 U935 ( .A(n1217), .B(G119), .ZN(n1243) );
INV_X1 U936 ( .A(G128), .ZN(n1217) );
NOR2_X1 U937 ( .A1(KEYINPUT32), .A2(n1244), .ZN(n1238) );
XNOR2_X1 U938 ( .A(G146), .B(n1102), .ZN(n1244) );
XNOR2_X1 U939 ( .A(G140), .B(n1245), .ZN(n1102) );
INV_X1 U940 ( .A(n1236), .ZN(n1240) );
XNOR2_X1 U941 ( .A(n1246), .B(G137), .ZN(n1236) );
NAND2_X1 U942 ( .A1(G221), .A2(n1247), .ZN(n1246) );
XOR2_X1 U943 ( .A(n1248), .B(G472), .Z(n1082) );
NAND2_X1 U944 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XNOR2_X1 U945 ( .A(n1251), .B(n1159), .ZN(n1249) );
XNOR2_X1 U946 ( .A(n1252), .B(G101), .ZN(n1159) );
NAND2_X1 U947 ( .A1(n1253), .A2(G210), .ZN(n1252) );
NAND2_X1 U948 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
OR2_X1 U949 ( .A1(n1158), .A2(n1161), .ZN(n1255) );
NAND2_X1 U950 ( .A1(n1256), .A2(n1158), .ZN(n1254) );
INV_X1 U951 ( .A(n1177), .ZN(n1158) );
XNOR2_X1 U952 ( .A(n1161), .B(KEYINPUT24), .ZN(n1256) );
XNOR2_X1 U953 ( .A(n1257), .B(n1258), .ZN(n1161) );
AND3_X1 U954 ( .A1(n1151), .A2(n1063), .A3(n1037), .ZN(n1218) );
NOR2_X1 U955 ( .A1(n1203), .A2(n1202), .ZN(n1037) );
INV_X1 U956 ( .A(n1206), .ZN(n1202) );
XOR2_X1 U957 ( .A(n1078), .B(G475), .Z(n1206) );
NAND2_X1 U958 ( .A1(n1146), .A2(n1250), .ZN(n1078) );
XOR2_X1 U959 ( .A(n1259), .B(n1260), .Z(n1146) );
XOR2_X1 U960 ( .A(G104), .B(n1261), .Z(n1260) );
NOR2_X1 U961 ( .A1(KEYINPUT3), .A2(n1262), .ZN(n1261) );
XOR2_X1 U962 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U963 ( .A(n1265), .B(n1266), .Z(n1264) );
NAND2_X1 U964 ( .A1(n1253), .A2(G214), .ZN(n1265) );
NOR2_X1 U965 ( .A1(G953), .A2(G237), .ZN(n1253) );
XOR2_X1 U966 ( .A(n1267), .B(G131), .Z(n1263) );
NAND4_X1 U967 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
OR2_X1 U968 ( .A1(n1245), .A2(KEYINPUT36), .ZN(n1271) );
NAND3_X1 U969 ( .A1(n1272), .A2(n1245), .A3(KEYINPUT36), .ZN(n1270) );
XNOR2_X1 U970 ( .A(KEYINPUT45), .B(n1207), .ZN(n1272) );
NAND3_X1 U971 ( .A1(KEYINPUT7), .A2(n1273), .A3(n1207), .ZN(n1269) );
OR2_X1 U972 ( .A1(n1274), .A2(KEYINPUT45), .ZN(n1273) );
NAND3_X1 U973 ( .A1(n1275), .A2(n1276), .A3(G140), .ZN(n1268) );
INV_X1 U974 ( .A(KEYINPUT7), .ZN(n1276) );
NAND2_X1 U975 ( .A1(KEYINPUT45), .A2(n1245), .ZN(n1275) );
XNOR2_X1 U976 ( .A(G113), .B(G122), .ZN(n1259) );
NAND2_X1 U977 ( .A1(n1277), .A2(n1278), .ZN(n1203) );
NAND2_X1 U978 ( .A1(n1279), .A2(n1076), .ZN(n1278) );
XNOR2_X1 U979 ( .A(KEYINPUT60), .B(n1144), .ZN(n1279) );
INV_X1 U980 ( .A(G478), .ZN(n1144) );
XOR2_X1 U981 ( .A(KEYINPUT25), .B(n1091), .Z(n1277) );
NOR2_X1 U982 ( .A1(n1076), .A2(G478), .ZN(n1091) );
NAND2_X1 U983 ( .A1(n1141), .A2(n1250), .ZN(n1076) );
XNOR2_X1 U984 ( .A(n1280), .B(n1281), .ZN(n1141) );
AND2_X1 U985 ( .A1(n1247), .A2(G217), .ZN(n1281) );
AND2_X1 U986 ( .A1(G234), .A2(n1028), .ZN(n1247) );
NAND2_X1 U987 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND2_X1 U988 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U989 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
OR2_X1 U990 ( .A1(n1288), .A2(KEYINPUT55), .ZN(n1287) );
INV_X1 U991 ( .A(KEYINPUT15), .ZN(n1286) );
NAND2_X1 U992 ( .A1(n1288), .A2(n1289), .ZN(n1282) );
NAND2_X1 U993 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
OR2_X1 U994 ( .A1(n1284), .A2(KEYINPUT15), .ZN(n1291) );
XOR2_X1 U995 ( .A(G128), .B(n1292), .Z(n1284) );
XNOR2_X1 U996 ( .A(G143), .B(n1210), .ZN(n1292) );
INV_X1 U997 ( .A(G134), .ZN(n1210) );
INV_X1 U998 ( .A(KEYINPUT55), .ZN(n1290) );
XOR2_X1 U999 ( .A(n1293), .B(n1294), .Z(n1288) );
XNOR2_X1 U1000 ( .A(KEYINPUT62), .B(n1295), .ZN(n1294) );
INV_X1 U1001 ( .A(G122), .ZN(n1295) );
XNOR2_X1 U1002 ( .A(G116), .B(n1296), .ZN(n1293) );
NAND2_X1 U1003 ( .A1(n1297), .A2(n1298), .ZN(n1063) );
OR3_X1 U1004 ( .A1(n1061), .A2(n1062), .A3(KEYINPUT29), .ZN(n1298) );
INV_X1 U1005 ( .A(n1299), .ZN(n1062) );
NAND2_X1 U1006 ( .A1(KEYINPUT29), .A2(n1038), .ZN(n1297) );
NOR2_X1 U1007 ( .A1(n1299), .A2(n1061), .ZN(n1038) );
INV_X1 U1008 ( .A(n1066), .ZN(n1061) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1232), .ZN(n1066) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1250), .ZN(n1232) );
NAND3_X1 U1011 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1299) );
INV_X1 U1012 ( .A(n1092), .ZN(n1302) );
NOR2_X1 U1013 ( .A1(n1093), .A2(G469), .ZN(n1092) );
NAND2_X1 U1014 ( .A1(KEYINPUT18), .A2(n1175), .ZN(n1301) );
INV_X1 U1015 ( .A(G469), .ZN(n1175) );
NAND3_X1 U1016 ( .A1(n1093), .A2(n1303), .A3(G469), .ZN(n1300) );
INV_X1 U1017 ( .A(KEYINPUT18), .ZN(n1303) );
NAND2_X1 U1018 ( .A1(n1304), .A2(n1250), .ZN(n1093) );
XOR2_X1 U1019 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1020 ( .A(n1307), .B(n1177), .ZN(n1306) );
XNOR2_X1 U1021 ( .A(n1308), .B(n1309), .ZN(n1177) );
XOR2_X1 U1022 ( .A(G131), .B(n1310), .Z(n1309) );
NOR2_X1 U1023 ( .A1(KEYINPUT43), .A2(n1111), .ZN(n1310) );
XNOR2_X1 U1024 ( .A(G134), .B(n1311), .ZN(n1111) );
XOR2_X1 U1025 ( .A(KEYINPUT23), .B(G137), .Z(n1311) );
XNOR2_X1 U1026 ( .A(KEYINPUT9), .B(KEYINPUT26), .ZN(n1308) );
NAND2_X1 U1027 ( .A1(n1312), .A2(n1313), .ZN(n1307) );
NAND2_X1 U1028 ( .A1(n1106), .A2(n1176), .ZN(n1313) );
XOR2_X1 U1029 ( .A(KEYINPUT0), .B(n1314), .Z(n1312) );
NOR2_X1 U1030 ( .A1(n1106), .A2(n1176), .ZN(n1314) );
XNOR2_X1 U1031 ( .A(n1315), .B(G101), .ZN(n1176) );
NAND2_X1 U1032 ( .A1(KEYINPUT4), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1033 ( .A(G128), .B(n1317), .Z(n1106) );
XOR2_X1 U1034 ( .A(KEYINPUT49), .B(n1318), .Z(n1305) );
NOR3_X1 U1035 ( .A1(n1319), .A2(KEYINPUT40), .A3(n1171), .ZN(n1318) );
AND2_X1 U1036 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U1037 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1038 ( .A(KEYINPUT42), .B(n1173), .ZN(n1321) );
XNOR2_X1 U1039 ( .A(n1322), .B(n1207), .ZN(n1173) );
INV_X1 U1040 ( .A(G140), .ZN(n1207) );
XOR2_X1 U1041 ( .A(KEYINPUT31), .B(n1172), .Z(n1320) );
AND2_X1 U1042 ( .A1(G227), .A2(n1028), .ZN(n1172) );
AND2_X1 U1043 ( .A1(n1215), .A2(n1323), .ZN(n1151) );
NAND2_X1 U1044 ( .A1(n1064), .A2(n1324), .ZN(n1323) );
NAND4_X1 U1045 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1325), .ZN(n1324) );
INV_X1 U1046 ( .A(G898), .ZN(n1325) );
NAND3_X1 U1047 ( .A1(n1220), .A2(n1028), .A3(G952), .ZN(n1064) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1220) );
NOR2_X1 U1049 ( .A1(n1043), .A2(n1051), .ZN(n1215) );
INV_X1 U1050 ( .A(n1046), .ZN(n1051) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1326), .ZN(n1046) );
XOR2_X1 U1052 ( .A(n1087), .B(n1327), .Z(n1043) );
NOR2_X1 U1053 ( .A1(n1090), .A2(KEYINPUT33), .ZN(n1327) );
INV_X1 U1054 ( .A(n1084), .ZN(n1090) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1326), .ZN(n1084) );
NAND2_X1 U1056 ( .A1(n1328), .A2(n1250), .ZN(n1326) );
INV_X1 U1057 ( .A(G902), .ZN(n1250) );
INV_X1 U1058 ( .A(G237), .ZN(n1328) );
NOR2_X1 U1059 ( .A1(n1180), .A2(G902), .ZN(n1087) );
XNOR2_X1 U1060 ( .A(n1329), .B(n1330), .ZN(n1180) );
XOR2_X1 U1061 ( .A(n1331), .B(n1332), .Z(n1330) );
NAND2_X1 U1062 ( .A1(G224), .A2(n1028), .ZN(n1332) );
INV_X1 U1063 ( .A(G953), .ZN(n1028) );
NAND3_X1 U1064 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1331) );
NAND2_X1 U1065 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
NAND2_X1 U1066 ( .A1(KEYINPUT41), .A2(n1338), .ZN(n1334) );
NAND3_X1 U1067 ( .A1(n1339), .A2(n1340), .A3(n1131), .ZN(n1338) );
INV_X1 U1068 ( .A(n1336), .ZN(n1131) );
NOR2_X1 U1069 ( .A1(n1341), .A2(n1342), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(n1337), .A2(n1343), .ZN(n1340) );
NAND3_X1 U1071 ( .A1(n1341), .A2(n1130), .A3(n1342), .ZN(n1339) );
INV_X1 U1072 ( .A(n1337), .ZN(n1130) );
NAND2_X1 U1073 ( .A1(n1127), .A2(n1344), .ZN(n1333) );
INV_X1 U1074 ( .A(KEYINPUT41), .ZN(n1344) );
NAND2_X1 U1075 ( .A1(n1345), .A2(n1346), .ZN(n1127) );
NAND2_X1 U1076 ( .A1(n1347), .A2(n1341), .ZN(n1346) );
XNOR2_X1 U1077 ( .A(n1337), .B(n1342), .ZN(n1347) );
INV_X1 U1078 ( .A(n1343), .ZN(n1342) );
OR3_X1 U1079 ( .A1(n1343), .A2(n1337), .A3(n1341), .ZN(n1345) );
XOR2_X1 U1080 ( .A(n1348), .B(n1349), .Z(n1341) );
XOR2_X1 U1081 ( .A(KEYINPUT58), .B(G101), .Z(n1349) );
NAND2_X1 U1082 ( .A1(KEYINPUT47), .A2(n1316), .ZN(n1348) );
XNOR2_X1 U1083 ( .A(G104), .B(n1296), .ZN(n1316) );
XOR2_X1 U1084 ( .A(G107), .B(KEYINPUT12), .Z(n1296) );
XOR2_X1 U1085 ( .A(n1258), .B(KEYINPUT34), .Z(n1337) );
XOR2_X1 U1086 ( .A(G113), .B(n1350), .Z(n1258) );
XOR2_X1 U1087 ( .A(G119), .B(G116), .Z(n1350) );
NAND2_X1 U1088 ( .A1(n1351), .A2(n1352), .ZN(n1343) );
NAND2_X1 U1089 ( .A1(G122), .A2(n1322), .ZN(n1352) );
XOR2_X1 U1090 ( .A(KEYINPUT57), .B(n1353), .Z(n1351) );
NOR2_X1 U1091 ( .A1(G122), .A2(n1322), .ZN(n1353) );
INV_X1 U1092 ( .A(G110), .ZN(n1322) );
XNOR2_X1 U1093 ( .A(n1257), .B(n1245), .ZN(n1329) );
INV_X1 U1094 ( .A(n1274), .ZN(n1245) );
XOR2_X1 U1095 ( .A(G125), .B(KEYINPUT10), .Z(n1274) );
XOR2_X1 U1096 ( .A(n1354), .B(n1317), .Z(n1257) );
XOR2_X1 U1097 ( .A(n1266), .B(KEYINPUT63), .Z(n1317) );
XOR2_X1 U1098 ( .A(G143), .B(G146), .Z(n1266) );
NAND2_X1 U1099 ( .A1(KEYINPUT35), .A2(G128), .ZN(n1354) );
endmodule


