//Key = 1000110001010111000001001011110000110110111100011011110110110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425, n1426, n1427, n1428;

XNOR2_X1 U785 ( .A(n1084), .B(n1085), .ZN(G9) );
NOR2_X1 U786 ( .A1(n1086), .A2(n1087), .ZN(G75) );
NOR4_X1 U787 ( .A1(n1088), .A2(n1089), .A3(G953), .A4(n1090), .ZN(n1087) );
NOR3_X1 U788 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
NAND3_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1088) );
NAND2_X1 U796 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
XOR2_X1 U797 ( .A(KEYINPUT60), .B(n1111), .Z(n1106) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
AND2_X1 U799 ( .A1(n1114), .A2(n1109), .ZN(n1113) );
NOR3_X1 U800 ( .A1(n1099), .A2(n1093), .A3(n1097), .ZN(n1109) );
INV_X1 U801 ( .A(n1115), .ZN(n1097) );
NOR3_X1 U802 ( .A1(n1091), .A2(n1116), .A3(n1093), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U804 ( .A1(n1119), .A2(n1099), .ZN(n1118) );
NOR3_X1 U805 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
AND2_X1 U806 ( .A1(n1115), .A2(KEYINPUT20), .ZN(n1122) );
NOR4_X1 U807 ( .A1(KEYINPUT20), .A2(n1123), .A3(n1103), .A4(n1124), .ZN(n1121) );
AND2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
AND3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1115), .ZN(n1117) );
NOR2_X1 U810 ( .A1(n1105), .A2(n1103), .ZN(n1115) );
NOR3_X1 U811 ( .A1(n1090), .A2(G953), .A3(G952), .ZN(n1086) );
AND4_X1 U812 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1090) );
NOR4_X1 U813 ( .A1(n1127), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1132) );
XOR2_X1 U814 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U815 ( .A(KEYINPUT25), .B(n1138), .ZN(n1136) );
NOR2_X1 U816 ( .A1(KEYINPUT12), .A2(n1139), .ZN(n1138) );
XNOR2_X1 U817 ( .A(G475), .B(n1140), .ZN(n1134) );
NOR2_X1 U818 ( .A1(n1141), .A2(KEYINPUT32), .ZN(n1140) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1144), .B(n1145), .Z(n1130) );
XNOR2_X1 U821 ( .A(KEYINPUT54), .B(n1146), .ZN(n1145) );
XOR2_X1 U822 ( .A(n1147), .B(KEYINPUT27), .Z(n1129) );
NAND2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XNOR2_X1 U824 ( .A(KEYINPUT59), .B(n1150), .ZN(n1148) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(G72) );
NOR2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n1157), .A2(n1158), .ZN(n1151) );
NAND2_X1 U829 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U830 ( .A(n1161), .B(n1162), .Z(n1159) );
NAND3_X1 U831 ( .A1(G900), .A2(n1162), .A3(G953), .ZN(n1157) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U833 ( .A(n1165), .B(n1166), .ZN(n1164) );
XOR2_X1 U834 ( .A(n1167), .B(KEYINPUT53), .Z(n1163) );
NAND2_X1 U835 ( .A1(KEYINPUT56), .A2(n1168), .ZN(n1167) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(G69) );
XOR2_X1 U837 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U838 ( .A1(n1173), .A2(n1154), .ZN(n1172) );
XNOR2_X1 U839 ( .A(G953), .B(KEYINPUT22), .ZN(n1154) );
AND2_X1 U840 ( .A1(G224), .A2(G898), .ZN(n1173) );
NAND2_X1 U841 ( .A1(n1160), .A2(n1174), .ZN(n1171) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
INV_X1 U843 ( .A(n1177), .ZN(n1176) );
XNOR2_X1 U844 ( .A(n1178), .B(KEYINPUT39), .ZN(n1175) );
NAND2_X1 U845 ( .A1(n1179), .A2(n1180), .ZN(n1169) );
INV_X1 U846 ( .A(n1181), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1183), .ZN(G66) );
XOR2_X1 U848 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U849 ( .A1(n1186), .A2(G217), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1182), .A2(n1187), .ZN(G63) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND3_X1 U852 ( .A1(n1186), .A2(G478), .A3(KEYINPUT52), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1182), .A2(n1190), .ZN(G60) );
NOR3_X1 U854 ( .A1(n1141), .A2(n1191), .A3(n1192), .ZN(n1190) );
AND3_X1 U855 ( .A1(n1193), .A2(G475), .A3(n1186), .ZN(n1192) );
NOR2_X1 U856 ( .A1(n1194), .A2(n1193), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1108), .A2(n1195), .ZN(n1194) );
INV_X1 U858 ( .A(G475), .ZN(n1195) );
XNOR2_X1 U859 ( .A(G104), .B(n1196), .ZN(G6) );
NOR2_X1 U860 ( .A1(n1182), .A2(n1197), .ZN(G57) );
XOR2_X1 U861 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U862 ( .A(n1200), .B(n1201), .ZN(n1199) );
XOR2_X1 U863 ( .A(n1202), .B(n1203), .Z(n1198) );
XOR2_X1 U864 ( .A(n1204), .B(n1205), .Z(n1203) );
NAND2_X1 U865 ( .A1(KEYINPUT34), .A2(n1206), .ZN(n1205) );
INV_X1 U866 ( .A(n1207), .ZN(n1206) );
NAND2_X1 U867 ( .A1(n1186), .A2(G472), .ZN(n1204) );
NOR2_X1 U868 ( .A1(n1182), .A2(n1208), .ZN(G54) );
XOR2_X1 U869 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U870 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U871 ( .A1(n1186), .A2(G469), .ZN(n1211) );
XOR2_X1 U872 ( .A(n1213), .B(n1214), .Z(n1209) );
XNOR2_X1 U873 ( .A(n1215), .B(KEYINPUT35), .ZN(n1214) );
NAND2_X1 U874 ( .A1(KEYINPUT58), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U875 ( .A(n1168), .B(n1217), .ZN(n1216) );
XNOR2_X1 U876 ( .A(n1218), .B(n1219), .ZN(n1217) );
NAND2_X1 U877 ( .A1(KEYINPUT11), .A2(n1220), .ZN(n1218) );
XOR2_X1 U878 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U879 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U880 ( .A(G101), .B(G128), .ZN(n1221) );
NOR3_X1 U881 ( .A1(n1155), .A2(KEYINPUT23), .A3(G953), .ZN(n1213) );
INV_X1 U882 ( .A(G227), .ZN(n1155) );
NOR2_X1 U883 ( .A1(n1182), .A2(n1225), .ZN(G51) );
XOR2_X1 U884 ( .A(n1226), .B(n1227), .Z(n1225) );
NAND2_X1 U885 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U886 ( .A1(n1179), .A2(n1230), .ZN(n1229) );
XOR2_X1 U887 ( .A(KEYINPUT0), .B(n1231), .Z(n1228) );
NOR2_X1 U888 ( .A1(n1179), .A2(n1230), .ZN(n1231) );
XOR2_X1 U889 ( .A(n1232), .B(n1233), .Z(n1230) );
NAND2_X1 U890 ( .A1(n1234), .A2(KEYINPUT62), .ZN(n1233) );
XNOR2_X1 U891 ( .A(n1235), .B(G125), .ZN(n1234) );
NAND3_X1 U892 ( .A1(n1236), .A2(n1237), .A3(n1137), .ZN(n1226) );
OR2_X1 U893 ( .A1(n1186), .A2(KEYINPUT7), .ZN(n1237) );
NOR2_X1 U894 ( .A1(n1238), .A2(n1108), .ZN(n1186) );
NAND2_X1 U895 ( .A1(KEYINPUT7), .A2(n1239), .ZN(n1236) );
NAND2_X1 U896 ( .A1(n1108), .A2(G902), .ZN(n1239) );
NOR3_X1 U897 ( .A1(n1177), .A2(n1178), .A3(n1161), .ZN(n1108) );
NAND4_X1 U898 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1161) );
NOR3_X1 U899 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
INV_X1 U900 ( .A(n1247), .ZN(n1245) );
NAND3_X1 U901 ( .A1(n1114), .A2(n1248), .A3(n1249), .ZN(n1242) );
NAND2_X1 U902 ( .A1(n1126), .A2(n1250), .ZN(n1241) );
NAND4_X1 U903 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
NAND2_X1 U904 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U905 ( .A(KEYINPUT47), .ZN(n1256) );
NAND2_X1 U906 ( .A1(n1257), .A2(n1110), .ZN(n1255) );
NAND2_X1 U907 ( .A1(n1257), .A2(n1258), .ZN(n1253) );
NAND2_X1 U908 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND2_X1 U909 ( .A1(KEYINPUT47), .A2(n1110), .ZN(n1260) );
XNOR2_X1 U910 ( .A(n1114), .B(KEYINPUT49), .ZN(n1259) );
OR2_X1 U911 ( .A1(n1261), .A2(KEYINPUT45), .ZN(n1252) );
NAND2_X1 U912 ( .A1(n1262), .A2(n1249), .ZN(n1251) );
NAND3_X1 U913 ( .A1(KEYINPUT45), .A2(n1263), .A3(n1105), .ZN(n1240) );
INV_X1 U914 ( .A(n1261), .ZN(n1263) );
NAND4_X1 U915 ( .A1(n1196), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1177) );
NOR4_X1 U916 ( .A1(n1267), .A2(n1085), .A3(n1268), .A4(n1269), .ZN(n1266) );
INV_X1 U917 ( .A(n1270), .ZN(n1269) );
NOR3_X1 U918 ( .A1(n1103), .A2(n1271), .A3(n1272), .ZN(n1085) );
INV_X1 U919 ( .A(n1273), .ZN(n1103) );
NAND4_X1 U920 ( .A1(n1262), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1265) );
XNOR2_X1 U921 ( .A(KEYINPUT1), .B(n1096), .ZN(n1276) );
NAND3_X1 U922 ( .A1(n1273), .A2(n1277), .A3(n1110), .ZN(n1196) );
NOR2_X1 U923 ( .A1(n1160), .A2(G952), .ZN(n1182) );
XNOR2_X1 U924 ( .A(n1278), .B(n1244), .ZN(G48) );
AND3_X1 U925 ( .A1(n1110), .A2(n1248), .A3(n1249), .ZN(n1244) );
XOR2_X1 U926 ( .A(G143), .B(n1246), .Z(G45) );
AND4_X1 U927 ( .A1(n1279), .A2(n1257), .A3(n1248), .A4(n1143), .ZN(n1246) );
XNOR2_X1 U928 ( .A(n1280), .B(n1281), .ZN(G42) );
NOR2_X1 U929 ( .A1(n1261), .A2(n1105), .ZN(n1281) );
INV_X1 U930 ( .A(n1126), .ZN(n1105) );
NAND4_X1 U931 ( .A1(n1125), .A2(n1110), .A3(n1282), .A4(n1283), .ZN(n1261) );
XNOR2_X1 U932 ( .A(G137), .B(n1284), .ZN(G39) );
NAND4_X1 U933 ( .A1(KEYINPUT40), .A2(n1126), .A3(n1262), .A4(n1249), .ZN(n1284) );
XOR2_X1 U934 ( .A(G134), .B(n1285), .Z(G36) );
NOR3_X1 U935 ( .A1(n1286), .A2(KEYINPUT6), .A3(n1272), .ZN(n1285) );
INV_X1 U936 ( .A(n1114), .ZN(n1272) );
XNOR2_X1 U937 ( .A(G131), .B(n1287), .ZN(G33) );
NAND2_X1 U938 ( .A1(n1288), .A2(n1110), .ZN(n1287) );
INV_X1 U939 ( .A(n1286), .ZN(n1288) );
NAND2_X1 U940 ( .A1(n1126), .A2(n1257), .ZN(n1286) );
NOR3_X1 U941 ( .A1(n1096), .A2(n1289), .A3(n1104), .ZN(n1257) );
INV_X1 U942 ( .A(n1282), .ZN(n1096) );
NOR2_X1 U943 ( .A1(n1124), .A2(n1133), .ZN(n1126) );
XNOR2_X1 U944 ( .A(G128), .B(n1290), .ZN(G30) );
NAND4_X1 U945 ( .A1(n1291), .A2(KEYINPUT55), .A3(n1249), .A4(n1114), .ZN(n1290) );
AND4_X1 U946 ( .A1(n1282), .A2(n1142), .A3(n1283), .A4(n1292), .ZN(n1249) );
XNOR2_X1 U947 ( .A(n1248), .B(KEYINPUT9), .ZN(n1291) );
XNOR2_X1 U948 ( .A(n1293), .B(n1294), .ZN(G3) );
NOR3_X1 U949 ( .A1(n1091), .A2(n1271), .A3(n1104), .ZN(n1294) );
INV_X1 U950 ( .A(n1262), .ZN(n1091) );
XNOR2_X1 U951 ( .A(n1295), .B(n1296), .ZN(G27) );
NOR2_X1 U952 ( .A1(KEYINPUT57), .A2(n1247), .ZN(n1296) );
NAND3_X1 U953 ( .A1(n1125), .A2(n1110), .A3(n1297), .ZN(n1247) );
NOR3_X1 U954 ( .A1(n1099), .A2(n1289), .A3(n1102), .ZN(n1297) );
INV_X1 U955 ( .A(n1248), .ZN(n1102) );
INV_X1 U956 ( .A(n1283), .ZN(n1289) );
NAND2_X1 U957 ( .A1(n1093), .A2(n1298), .ZN(n1283) );
NAND4_X1 U958 ( .A1(G902), .A2(G953), .A3(n1299), .A4(n1156), .ZN(n1298) );
INV_X1 U959 ( .A(G900), .ZN(n1156) );
XNOR2_X1 U960 ( .A(G122), .B(n1264), .ZN(G24) );
NAND4_X1 U961 ( .A1(n1279), .A2(n1300), .A3(n1273), .A4(n1143), .ZN(n1264) );
NOR2_X1 U962 ( .A1(n1292), .A2(n1142), .ZN(n1273) );
XNOR2_X1 U963 ( .A(G119), .B(n1270), .ZN(G21) );
NAND4_X1 U964 ( .A1(n1262), .A2(n1300), .A3(n1142), .A4(n1292), .ZN(n1270) );
NAND2_X1 U965 ( .A1(n1301), .A2(n1302), .ZN(G18) );
NAND2_X1 U966 ( .A1(n1178), .A2(n1303), .ZN(n1302) );
XOR2_X1 U967 ( .A(KEYINPUT15), .B(n1304), .Z(n1301) );
NOR2_X1 U968 ( .A1(n1178), .A2(n1303), .ZN(n1304) );
AND3_X1 U969 ( .A1(n1300), .A2(n1114), .A3(n1274), .ZN(n1178) );
NOR2_X1 U970 ( .A1(n1305), .A2(n1279), .ZN(n1114) );
INV_X1 U971 ( .A(n1143), .ZN(n1305) );
XOR2_X1 U972 ( .A(G113), .B(n1268), .Z(G15) );
AND3_X1 U973 ( .A1(n1274), .A2(n1300), .A3(n1110), .ZN(n1268) );
AND2_X1 U974 ( .A1(n1306), .A2(n1279), .ZN(n1110) );
XNOR2_X1 U975 ( .A(n1143), .B(KEYINPUT46), .ZN(n1306) );
NOR2_X1 U976 ( .A1(n1099), .A2(n1307), .ZN(n1300) );
NAND2_X1 U977 ( .A1(n1128), .A2(n1308), .ZN(n1099) );
INV_X1 U978 ( .A(n1104), .ZN(n1274) );
NAND2_X1 U979 ( .A1(n1309), .A2(n1142), .ZN(n1104) );
XOR2_X1 U980 ( .A(n1267), .B(n1310), .Z(G12) );
NOR2_X1 U981 ( .A1(KEYINPUT44), .A2(n1311), .ZN(n1310) );
AND3_X1 U982 ( .A1(n1125), .A2(n1277), .A3(n1262), .ZN(n1267) );
NOR2_X1 U983 ( .A1(n1143), .A2(n1279), .ZN(n1262) );
XOR2_X1 U984 ( .A(G475), .B(n1312), .Z(n1279) );
NOR2_X1 U985 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NOR2_X1 U986 ( .A1(KEYINPUT30), .A2(n1141), .ZN(n1314) );
NOR2_X1 U987 ( .A1(KEYINPUT26), .A2(n1315), .ZN(n1313) );
INV_X1 U988 ( .A(n1141), .ZN(n1315) );
NOR2_X1 U989 ( .A1(n1193), .A2(G902), .ZN(n1141) );
XNOR2_X1 U990 ( .A(n1316), .B(n1317), .ZN(n1193) );
XNOR2_X1 U991 ( .A(n1318), .B(n1319), .ZN(n1317) );
NOR3_X1 U992 ( .A1(n1320), .A2(KEYINPUT31), .A3(n1321), .ZN(n1319) );
NOR2_X1 U993 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U994 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U995 ( .A(KEYINPUT50), .B(KEYINPUT28), .Z(n1325) );
NOR2_X1 U996 ( .A1(n1326), .A2(n1324), .ZN(n1322) );
AND2_X1 U997 ( .A1(n1327), .A2(KEYINPUT24), .ZN(n1326) );
NOR2_X1 U998 ( .A1(n1328), .A2(n1327), .ZN(n1320) );
XOR2_X1 U999 ( .A(n1329), .B(n1166), .Z(n1327) );
XOR2_X1 U1000 ( .A(G125), .B(G140), .Z(n1166) );
XNOR2_X1 U1001 ( .A(G146), .B(KEYINPUT3), .ZN(n1329) );
NOR2_X1 U1002 ( .A1(n1324), .A2(n1330), .ZN(n1328) );
INV_X1 U1003 ( .A(KEYINPUT24), .ZN(n1330) );
XNOR2_X1 U1004 ( .A(n1331), .B(n1332), .ZN(n1324) );
XNOR2_X1 U1005 ( .A(n1333), .B(n1219), .ZN(n1331) );
INV_X1 U1006 ( .A(G131), .ZN(n1219) );
NAND2_X1 U1007 ( .A1(G214), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1008 ( .A(G113), .B(G122), .ZN(n1316) );
XNOR2_X1 U1009 ( .A(n1335), .B(G478), .ZN(n1143) );
NAND2_X1 U1010 ( .A1(n1189), .A2(n1238), .ZN(n1335) );
XOR2_X1 U1011 ( .A(n1336), .B(n1337), .Z(n1189) );
XOR2_X1 U1012 ( .A(n1338), .B(n1339), .Z(n1337) );
XNOR2_X1 U1013 ( .A(n1303), .B(G107), .ZN(n1339) );
INV_X1 U1014 ( .A(G116), .ZN(n1303) );
XOR2_X1 U1015 ( .A(G128), .B(G122), .Z(n1338) );
XOR2_X1 U1016 ( .A(n1340), .B(n1341), .Z(n1336) );
XNOR2_X1 U1017 ( .A(n1342), .B(n1332), .ZN(n1340) );
NAND3_X1 U1018 ( .A1(n1343), .A2(n1160), .A3(G217), .ZN(n1342) );
XNOR2_X1 U1019 ( .A(KEYINPUT18), .B(n1344), .ZN(n1343) );
INV_X1 U1020 ( .A(n1271), .ZN(n1277) );
NAND2_X1 U1021 ( .A1(n1282), .A2(n1275), .ZN(n1271) );
INV_X1 U1022 ( .A(n1307), .ZN(n1275) );
NAND2_X1 U1023 ( .A1(n1248), .A2(n1345), .ZN(n1307) );
NAND2_X1 U1024 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND3_X1 U1025 ( .A1(n1181), .A2(n1299), .A3(G902), .ZN(n1347) );
NOR2_X1 U1026 ( .A1(n1160), .A2(G898), .ZN(n1181) );
XNOR2_X1 U1027 ( .A(KEYINPUT41), .B(n1093), .ZN(n1346) );
NAND3_X1 U1028 ( .A1(n1299), .A2(n1160), .A3(G952), .ZN(n1093) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1299) );
NOR2_X1 U1030 ( .A1(n1348), .A2(n1133), .ZN(n1248) );
INV_X1 U1031 ( .A(n1123), .ZN(n1133) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1349), .ZN(n1123) );
INV_X1 U1033 ( .A(n1124), .ZN(n1348) );
XOR2_X1 U1034 ( .A(n1139), .B(n1137), .Z(n1124) );
AND2_X1 U1035 ( .A1(G210), .A2(n1349), .ZN(n1137) );
NAND2_X1 U1036 ( .A1(n1350), .A2(n1238), .ZN(n1349) );
INV_X1 U1037 ( .A(G237), .ZN(n1350) );
AND2_X1 U1038 ( .A1(n1351), .A2(n1238), .ZN(n1139) );
XOR2_X1 U1039 ( .A(n1179), .B(n1352), .Z(n1351) );
XOR2_X1 U1040 ( .A(n1232), .B(n1353), .Z(n1352) );
NAND2_X1 U1041 ( .A1(KEYINPUT38), .A2(n1354), .ZN(n1353) );
XNOR2_X1 U1042 ( .A(G125), .B(n1355), .ZN(n1354) );
INV_X1 U1043 ( .A(n1235), .ZN(n1355) );
NAND2_X1 U1044 ( .A1(G224), .A2(n1160), .ZN(n1232) );
XOR2_X1 U1045 ( .A(n1356), .B(n1357), .Z(n1179) );
XNOR2_X1 U1046 ( .A(G122), .B(n1311), .ZN(n1357) );
XOR2_X1 U1047 ( .A(n1358), .B(n1359), .Z(n1356) );
NOR2_X1 U1048 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NOR2_X1 U1049 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
XNOR2_X1 U1050 ( .A(n1364), .B(n1293), .ZN(n1363) );
INV_X1 U1051 ( .A(G101), .ZN(n1293) );
XNOR2_X1 U1052 ( .A(KEYINPUT21), .B(KEYINPUT14), .ZN(n1364) );
NOR3_X1 U1053 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1362) );
NOR2_X1 U1054 ( .A1(n1084), .A2(n1368), .ZN(n1367) );
NOR2_X1 U1055 ( .A1(KEYINPUT37), .A2(G107), .ZN(n1366) );
NOR2_X1 U1056 ( .A1(G101), .A2(n1369), .ZN(n1360) );
XNOR2_X1 U1057 ( .A(n1368), .B(n1084), .ZN(n1369) );
NAND2_X1 U1058 ( .A1(KEYINPUT37), .A2(n1318), .ZN(n1368) );
NAND2_X1 U1059 ( .A1(n1370), .A2(n1371), .ZN(n1358) );
OR2_X1 U1060 ( .A1(n1372), .A2(G113), .ZN(n1371) );
XOR2_X1 U1061 ( .A(n1373), .B(KEYINPUT33), .Z(n1370) );
NAND2_X1 U1062 ( .A1(G113), .A2(n1372), .ZN(n1373) );
XNOR2_X1 U1063 ( .A(G116), .B(n1374), .ZN(n1372) );
NOR2_X1 U1064 ( .A1(n1128), .A2(n1127), .ZN(n1282) );
INV_X1 U1065 ( .A(n1308), .ZN(n1127) );
NAND2_X1 U1066 ( .A1(G221), .A2(n1375), .ZN(n1308) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1238), .ZN(n1375) );
XOR2_X1 U1068 ( .A(n1376), .B(n1144), .Z(n1128) );
NAND4_X1 U1069 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1238), .ZN(n1144) );
NAND3_X1 U1070 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1379) );
NAND2_X1 U1071 ( .A1(G227), .A2(n1160), .ZN(n1382) );
NAND2_X1 U1072 ( .A1(n1383), .A2(n1384), .ZN(n1380) );
NAND2_X1 U1073 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
INV_X1 U1074 ( .A(KEYINPUT63), .ZN(n1386) );
NAND3_X1 U1075 ( .A1(n1387), .A2(n1160), .A3(G227), .ZN(n1378) );
NAND2_X1 U1076 ( .A1(n1381), .A2(n1388), .ZN(n1387) );
OR3_X1 U1077 ( .A1(n1385), .A2(KEYINPUT63), .A3(n1389), .ZN(n1388) );
NAND2_X1 U1078 ( .A1(n1385), .A2(n1389), .ZN(n1381) );
NOR2_X1 U1079 ( .A1(KEYINPUT36), .A2(n1212), .ZN(n1385) );
XNOR2_X1 U1080 ( .A(G110), .B(G140), .ZN(n1212) );
NAND2_X1 U1081 ( .A1(KEYINPUT63), .A2(n1389), .ZN(n1377) );
INV_X1 U1082 ( .A(n1383), .ZN(n1389) );
XNOR2_X1 U1083 ( .A(n1390), .B(n1391), .ZN(n1383) );
XNOR2_X1 U1084 ( .A(n1224), .B(n1165), .ZN(n1391) );
XOR2_X1 U1085 ( .A(n1223), .B(n1200), .Z(n1165) );
XOR2_X1 U1086 ( .A(G131), .B(G128), .Z(n1200) );
NAND2_X1 U1087 ( .A1(KEYINPUT61), .A2(n1392), .ZN(n1223) );
XNOR2_X1 U1088 ( .A(G146), .B(n1332), .ZN(n1392) );
NOR2_X1 U1089 ( .A1(n1393), .A2(n1365), .ZN(n1224) );
NOR2_X1 U1090 ( .A1(n1318), .A2(G107), .ZN(n1365) );
INV_X1 U1091 ( .A(G104), .ZN(n1318) );
XNOR2_X1 U1092 ( .A(KEYINPUT48), .B(n1394), .ZN(n1393) );
NOR2_X1 U1093 ( .A1(G104), .A2(n1084), .ZN(n1394) );
INV_X1 U1094 ( .A(G107), .ZN(n1084) );
NAND2_X1 U1095 ( .A1(KEYINPUT29), .A2(n1146), .ZN(n1376) );
INV_X1 U1096 ( .A(G469), .ZN(n1146) );
NOR2_X1 U1097 ( .A1(n1142), .A2(n1309), .ZN(n1125) );
INV_X1 U1098 ( .A(n1292), .ZN(n1309) );
NAND2_X1 U1099 ( .A1(n1150), .A2(n1149), .ZN(n1292) );
NAND2_X1 U1100 ( .A1(G217), .A2(n1395), .ZN(n1149) );
NAND2_X1 U1101 ( .A1(n1238), .A2(n1396), .ZN(n1395) );
OR2_X1 U1102 ( .A1(n1184), .A2(G234), .ZN(n1396) );
NAND3_X1 U1103 ( .A1(n1184), .A2(n1238), .A3(n1397), .ZN(n1150) );
NAND2_X1 U1104 ( .A1(G217), .A2(n1344), .ZN(n1397) );
INV_X1 U1105 ( .A(G234), .ZN(n1344) );
NAND2_X1 U1106 ( .A1(n1398), .A2(n1399), .ZN(n1184) );
OR2_X1 U1107 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
XOR2_X1 U1108 ( .A(n1402), .B(KEYINPUT2), .Z(n1398) );
NAND2_X1 U1109 ( .A1(n1401), .A2(n1400), .ZN(n1402) );
NAND2_X1 U1110 ( .A1(n1403), .A2(n1404), .ZN(n1400) );
NAND2_X1 U1111 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
XOR2_X1 U1112 ( .A(n1407), .B(KEYINPUT16), .Z(n1403) );
OR2_X1 U1113 ( .A1(n1406), .A2(n1405), .ZN(n1407) );
NAND3_X1 U1114 ( .A1(G234), .A2(n1160), .A3(G221), .ZN(n1405) );
INV_X1 U1115 ( .A(G953), .ZN(n1160) );
INV_X1 U1116 ( .A(G137), .ZN(n1406) );
XNOR2_X1 U1117 ( .A(n1408), .B(n1409), .ZN(n1401) );
XNOR2_X1 U1118 ( .A(n1311), .B(n1410), .ZN(n1409) );
NOR2_X1 U1119 ( .A1(KEYINPUT8), .A2(n1411), .ZN(n1410) );
NOR3_X1 U1120 ( .A1(n1412), .A2(n1413), .A3(n1414), .ZN(n1411) );
NOR2_X1 U1121 ( .A1(n1415), .A2(n1278), .ZN(n1414) );
AND3_X1 U1122 ( .A1(n1278), .A2(n1415), .A3(KEYINPUT43), .ZN(n1413) );
NOR2_X1 U1123 ( .A1(KEYINPUT19), .A2(n1416), .ZN(n1415) );
NOR2_X1 U1124 ( .A1(KEYINPUT43), .A2(n1417), .ZN(n1412) );
INV_X1 U1125 ( .A(n1416), .ZN(n1417) );
XOR2_X1 U1126 ( .A(n1418), .B(n1295), .Z(n1416) );
INV_X1 U1127 ( .A(G125), .ZN(n1295) );
NAND2_X1 U1128 ( .A1(KEYINPUT51), .A2(n1280), .ZN(n1418) );
INV_X1 U1129 ( .A(G140), .ZN(n1280) );
INV_X1 U1130 ( .A(G110), .ZN(n1311) );
XNOR2_X1 U1131 ( .A(G119), .B(G128), .ZN(n1408) );
XNOR2_X1 U1132 ( .A(n1419), .B(G472), .ZN(n1142) );
NAND2_X1 U1133 ( .A1(n1420), .A2(n1238), .ZN(n1419) );
INV_X1 U1134 ( .A(G902), .ZN(n1238) );
XOR2_X1 U1135 ( .A(n1421), .B(n1422), .Z(n1420) );
XOR2_X1 U1136 ( .A(n1423), .B(n1201), .Z(n1422) );
XOR2_X1 U1137 ( .A(n1424), .B(n1425), .Z(n1201) );
XOR2_X1 U1138 ( .A(G113), .B(n1426), .Z(n1425) );
XNOR2_X1 U1139 ( .A(KEYINPUT42), .B(n1374), .ZN(n1426) );
INV_X1 U1140 ( .A(G119), .ZN(n1374) );
XOR2_X1 U1141 ( .A(n1390), .B(n1427), .Z(n1424) );
NOR2_X1 U1142 ( .A1(G116), .A2(KEYINPUT10), .ZN(n1427) );
XNOR2_X1 U1143 ( .A(n1168), .B(G101), .ZN(n1390) );
XOR2_X1 U1144 ( .A(G137), .B(n1341), .Z(n1168) );
XOR2_X1 U1145 ( .A(G134), .B(KEYINPUT13), .Z(n1341) );
NAND2_X1 U1146 ( .A1(KEYINPUT4), .A2(n1235), .ZN(n1423) );
XNOR2_X1 U1147 ( .A(n1202), .B(G128), .ZN(n1235) );
XNOR2_X1 U1148 ( .A(n1428), .B(n1278), .ZN(n1202) );
INV_X1 U1149 ( .A(G146), .ZN(n1278) );
NAND2_X1 U1150 ( .A1(KEYINPUT5), .A2(n1332), .ZN(n1428) );
XNOR2_X1 U1151 ( .A(G143), .B(KEYINPUT17), .ZN(n1332) );
XNOR2_X1 U1152 ( .A(G131), .B(n1207), .ZN(n1421) );
NAND2_X1 U1153 ( .A1(G210), .A2(n1334), .ZN(n1207) );
NOR2_X1 U1154 ( .A1(G953), .A2(G237), .ZN(n1334) );
endmodule


