//Key = 0001100110010101111000100011111001010110100111010000101100110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;

XOR2_X1 U776 ( .A(G107), .B(n1061), .Z(G9) );
NOR2_X1 U777 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR3_X1 U778 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NAND3_X1 U779 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1064) );
NAND2_X1 U780 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U781 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U782 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U783 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND3_X1 U784 ( .A1(n1079), .A2(n1080), .A3(KEYINPUT19), .ZN(n1077) );
NAND3_X1 U785 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1074) );
NAND2_X1 U786 ( .A1(n1079), .A2(n1084), .ZN(n1082) );
NAND2_X1 U787 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
OR2_X1 U788 ( .A1(n1087), .A2(KEYINPUT19), .ZN(n1086) );
INV_X1 U789 ( .A(n1088), .ZN(n1085) );
NAND2_X1 U790 ( .A1(n1089), .A2(n1090), .ZN(n1081) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U792 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U793 ( .A1(n1089), .A2(n1095), .A3(n1079), .ZN(n1072) );
NAND2_X1 U794 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U795 ( .A1(n1083), .A2(n1098), .ZN(n1097) );
NAND2_X1 U796 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U797 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U798 ( .A1(n1076), .A2(n1103), .ZN(n1096) );
NAND2_X1 U799 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
INV_X1 U801 ( .A(n1108), .ZN(n1070) );
NOR3_X1 U802 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1062) );
INV_X1 U803 ( .A(n1067), .ZN(n1109) );
NAND4_X1 U804 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1067) );
NOR4_X1 U805 ( .A1(n1114), .A2(n1093), .A3(n1115), .A4(n1078), .ZN(n1113) );
XNOR2_X1 U806 ( .A(n1116), .B(KEYINPUT27), .ZN(n1115) );
NOR3_X1 U807 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1112) );
NOR3_X1 U808 ( .A1(n1120), .A2(G902), .A3(n1121), .ZN(n1119) );
AND2_X1 U809 ( .A1(n1122), .A2(n1120), .ZN(n1118) );
XOR2_X1 U810 ( .A(G472), .B(KEYINPUT9), .Z(n1120) );
XNOR2_X1 U811 ( .A(G478), .B(n1123), .ZN(n1117) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1111) );
NOR2_X1 U813 ( .A1(KEYINPUT56), .A2(n1126), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1127), .B(KEYINPUT31), .Z(n1110) );
NAND2_X1 U815 ( .A1(G475), .A2(n1128), .ZN(n1127) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(G72) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U818 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XNOR2_X1 U819 ( .A(G953), .B(KEYINPUT26), .ZN(n1134) );
INV_X1 U820 ( .A(n1066), .ZN(n1133) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1068), .ZN(n1131) );
NOR2_X1 U822 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U823 ( .A(G900), .B(KEYINPUT2), .ZN(n1136) );
NOR2_X1 U824 ( .A1(n1138), .A2(n1139), .ZN(n1129) );
XOR2_X1 U825 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U826 ( .A(n1142), .B(n1143), .Z(n1140) );
NOR2_X1 U827 ( .A1(KEYINPUT57), .A2(n1144), .ZN(n1143) );
XNOR2_X1 U828 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U829 ( .A1(G134), .A2(KEYINPUT53), .ZN(n1146) );
NAND4_X1 U830 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1142) );
NAND3_X1 U831 ( .A1(KEYINPUT7), .A2(n1151), .A3(n1152), .ZN(n1150) );
NAND2_X1 U832 ( .A1(n1153), .A2(G125), .ZN(n1149) );
INV_X1 U833 ( .A(n1152), .ZN(n1153) );
XNOR2_X1 U834 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n1152) );
NAND2_X1 U835 ( .A1(G140), .A2(n1154), .ZN(n1147) );
INV_X1 U836 ( .A(KEYINPUT7), .ZN(n1154) );
NAND2_X1 U837 ( .A1(n1155), .A2(n1156), .ZN(G69) );
NAND2_X1 U838 ( .A1(n1157), .A2(n1068), .ZN(n1156) );
XNOR2_X1 U839 ( .A(n1065), .B(n1158), .ZN(n1157) );
NAND2_X1 U840 ( .A1(n1159), .A2(G953), .ZN(n1155) );
NAND2_X1 U841 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U842 ( .A1(n1158), .A2(n1162), .ZN(n1161) );
NAND2_X1 U843 ( .A1(G224), .A2(n1163), .ZN(n1160) );
NAND2_X1 U844 ( .A1(G898), .A2(n1158), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NAND2_X1 U846 ( .A1(G953), .A2(n1166), .ZN(n1165) );
XOR2_X1 U847 ( .A(n1167), .B(n1168), .Z(n1164) );
NAND2_X1 U848 ( .A1(KEYINPUT58), .A2(n1169), .ZN(n1167) );
NOR2_X1 U849 ( .A1(n1170), .A2(n1171), .ZN(G66) );
XNOR2_X1 U850 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U851 ( .A1(n1124), .A2(n1174), .ZN(n1173) );
NOR2_X1 U852 ( .A1(n1170), .A2(n1175), .ZN(G63) );
NOR2_X1 U853 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U854 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U855 ( .A1(KEYINPUT5), .A2(n1180), .ZN(n1179) );
NOR2_X1 U856 ( .A1(n1181), .A2(n1174), .ZN(n1178) );
AND2_X1 U857 ( .A1(n1180), .A2(KEYINPUT5), .ZN(n1176) );
NOR2_X1 U858 ( .A1(n1170), .A2(n1182), .ZN(G60) );
NOR2_X1 U859 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NOR2_X1 U860 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U861 ( .A(n1187), .ZN(n1186) );
NOR2_X1 U862 ( .A1(n1188), .A2(n1189), .ZN(n1183) );
XNOR2_X1 U863 ( .A(n1187), .B(KEYINPUT15), .ZN(n1189) );
XNOR2_X1 U864 ( .A(n1185), .B(KEYINPUT39), .ZN(n1188) );
NOR2_X1 U865 ( .A1(n1174), .A2(n1190), .ZN(n1185) );
INV_X1 U866 ( .A(G475), .ZN(n1190) );
XNOR2_X1 U867 ( .A(n1191), .B(n1192), .ZN(G6) );
NOR2_X1 U868 ( .A1(n1193), .A2(n1194), .ZN(G57) );
XOR2_X1 U869 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U870 ( .A(n1197), .B(n1198), .Z(n1196) );
NAND2_X1 U871 ( .A1(KEYINPUT47), .A2(n1199), .ZN(n1197) );
XOR2_X1 U872 ( .A(n1200), .B(n1201), .Z(n1195) );
XOR2_X1 U873 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U874 ( .A1(KEYINPUT51), .A2(n1204), .ZN(n1203) );
INV_X1 U875 ( .A(n1205), .ZN(n1204) );
NOR2_X1 U876 ( .A1(n1206), .A2(n1174), .ZN(n1200) );
NOR2_X1 U877 ( .A1(G952), .A2(n1207), .ZN(n1193) );
XNOR2_X1 U878 ( .A(G953), .B(KEYINPUT61), .ZN(n1207) );
NOR2_X1 U879 ( .A1(n1170), .A2(n1208), .ZN(G54) );
XOR2_X1 U880 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U881 ( .A1(n1211), .A2(n1174), .ZN(n1210) );
NAND2_X1 U882 ( .A1(n1212), .A2(KEYINPUT35), .ZN(n1209) );
XOR2_X1 U883 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND2_X1 U884 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
NAND2_X1 U885 ( .A1(KEYINPUT11), .A2(n1217), .ZN(n1216) );
NAND3_X1 U886 ( .A1(G140), .A2(n1218), .A3(n1219), .ZN(n1215) );
INV_X1 U887 ( .A(KEYINPUT11), .ZN(n1219) );
NOR2_X1 U888 ( .A1(n1170), .A2(n1220), .ZN(G51) );
XOR2_X1 U889 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U890 ( .A(n1223), .B(n1224), .ZN(n1222) );
NOR3_X1 U891 ( .A1(n1174), .A2(KEYINPUT23), .A3(n1225), .ZN(n1224) );
NAND2_X1 U892 ( .A1(n1226), .A2(n1227), .ZN(n1174) );
OR2_X1 U893 ( .A1(n1066), .A2(n1065), .ZN(n1227) );
NAND4_X1 U894 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1065) );
NOR4_X1 U895 ( .A1(n1061), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1231) );
INV_X1 U896 ( .A(n1235), .ZN(n1234) );
AND2_X1 U897 ( .A1(n1088), .A2(n1236), .ZN(n1061) );
NOR2_X1 U898 ( .A1(n1237), .A2(n1192), .ZN(n1230) );
AND2_X1 U899 ( .A1(n1080), .A2(n1236), .ZN(n1192) );
AND3_X1 U900 ( .A1(n1238), .A2(n1076), .A3(n1239), .ZN(n1236) );
NAND2_X1 U901 ( .A1(n1240), .A2(n1241), .ZN(n1229) );
NAND2_X1 U902 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND3_X1 U903 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
INV_X1 U904 ( .A(KEYINPUT33), .ZN(n1245) );
XOR2_X1 U905 ( .A(n1247), .B(KEYINPUT63), .Z(n1242) );
NAND2_X1 U906 ( .A1(KEYINPUT33), .A2(n1248), .ZN(n1228) );
NAND4_X1 U907 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1066) );
NOR4_X1 U908 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1252) );
NOR3_X1 U909 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1251) );
NOR4_X1 U910 ( .A1(n1260), .A2(n1261), .A3(n1099), .A4(n1087), .ZN(n1259) );
INV_X1 U911 ( .A(n1080), .ZN(n1087) );
INV_X1 U912 ( .A(n1262), .ZN(n1099) );
NAND3_X1 U913 ( .A1(n1263), .A2(n1091), .A3(n1083), .ZN(n1261) );
INV_X1 U914 ( .A(n1239), .ZN(n1091) );
INV_X1 U915 ( .A(KEYINPUT32), .ZN(n1260) );
NOR2_X1 U916 ( .A1(KEYINPUT32), .A2(n1264), .ZN(n1258) );
XNOR2_X1 U917 ( .A(G902), .B(KEYINPUT44), .ZN(n1226) );
NAND2_X1 U918 ( .A1(KEYINPUT29), .A2(n1265), .ZN(n1223) );
XOR2_X1 U919 ( .A(G125), .B(n1266), .Z(n1265) );
NOR2_X1 U920 ( .A1(KEYINPUT50), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U921 ( .A(n1268), .B(KEYINPUT62), .ZN(n1267) );
NOR2_X1 U922 ( .A1(n1068), .A2(G952), .ZN(n1170) );
XNOR2_X1 U923 ( .A(n1269), .B(n1257), .ZN(G48) );
AND3_X1 U924 ( .A1(n1270), .A2(n1240), .A3(n1080), .ZN(n1257) );
XOR2_X1 U925 ( .A(G143), .B(n1256), .Z(G45) );
AND4_X1 U926 ( .A1(n1271), .A2(n1240), .A3(n1272), .A4(n1273), .ZN(n1256) );
XNOR2_X1 U927 ( .A(G140), .B(n1249), .ZN(G42) );
NAND3_X1 U928 ( .A1(n1101), .A2(n1102), .A3(n1274), .ZN(n1249) );
XOR2_X1 U929 ( .A(n1255), .B(n1275), .Z(G39) );
NOR2_X1 U930 ( .A1(KEYINPUT10), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U931 ( .A(G137), .B(KEYINPUT49), .ZN(n1276) );
AND3_X1 U932 ( .A1(n1270), .A2(n1083), .A3(n1089), .ZN(n1255) );
XOR2_X1 U933 ( .A(G134), .B(n1254), .Z(G36) );
AND3_X1 U934 ( .A1(n1083), .A2(n1088), .A3(n1271), .ZN(n1254) );
AND3_X1 U935 ( .A1(n1239), .A2(n1263), .A3(n1262), .ZN(n1271) );
XNOR2_X1 U936 ( .A(G131), .B(n1264), .ZN(G33) );
NAND2_X1 U937 ( .A1(n1274), .A2(n1262), .ZN(n1264) );
AND4_X1 U938 ( .A1(n1080), .A2(n1083), .A3(n1239), .A4(n1263), .ZN(n1274) );
INV_X1 U939 ( .A(n1078), .ZN(n1083) );
NAND2_X1 U940 ( .A1(n1107), .A2(n1277), .ZN(n1078) );
XNOR2_X1 U941 ( .A(G128), .B(n1278), .ZN(G30) );
NAND2_X1 U942 ( .A1(KEYINPUT37), .A2(n1253), .ZN(n1278) );
AND3_X1 U943 ( .A1(n1088), .A2(n1240), .A3(n1270), .ZN(n1253) );
AND4_X1 U944 ( .A1(n1239), .A2(n1102), .A3(n1263), .A4(n1279), .ZN(n1270) );
XOR2_X1 U945 ( .A(G101), .B(n1280), .Z(G3) );
NOR2_X1 U946 ( .A1(n1104), .A2(n1247), .ZN(n1280) );
NAND4_X1 U947 ( .A1(n1089), .A2(n1262), .A3(n1239), .A4(n1281), .ZN(n1247) );
NAND2_X1 U948 ( .A1(n1282), .A2(n1283), .ZN(G27) );
OR2_X1 U949 ( .A1(n1250), .A2(G125), .ZN(n1283) );
XOR2_X1 U950 ( .A(n1284), .B(KEYINPUT1), .Z(n1282) );
NAND2_X1 U951 ( .A1(G125), .A2(n1250), .ZN(n1284) );
NAND4_X1 U952 ( .A1(n1102), .A2(n1263), .A3(n1240), .A4(n1285), .ZN(n1250) );
AND3_X1 U953 ( .A1(n1079), .A2(n1101), .A3(n1080), .ZN(n1285) );
NAND2_X1 U954 ( .A1(n1108), .A2(n1286), .ZN(n1263) );
NAND3_X1 U955 ( .A1(G902), .A2(n1287), .A3(n1138), .ZN(n1286) );
NOR2_X1 U956 ( .A1(n1068), .A2(G900), .ZN(n1138) );
XNOR2_X1 U957 ( .A(n1288), .B(n1248), .ZN(G24) );
AND2_X1 U958 ( .A1(n1246), .A2(n1238), .ZN(n1248) );
AND4_X1 U959 ( .A1(n1079), .A2(n1076), .A3(n1272), .A4(n1273), .ZN(n1246) );
NOR2_X1 U960 ( .A1(n1279), .A2(n1102), .ZN(n1076) );
XNOR2_X1 U961 ( .A(n1237), .B(n1289), .ZN(G21) );
NAND2_X1 U962 ( .A1(KEYINPUT13), .A2(G119), .ZN(n1289) );
AND3_X1 U963 ( .A1(n1079), .A2(n1279), .A3(n1290), .ZN(n1237) );
XNOR2_X1 U964 ( .A(n1291), .B(n1292), .ZN(G18) );
NOR2_X1 U965 ( .A1(KEYINPUT12), .A2(n1235), .ZN(n1292) );
NAND2_X1 U966 ( .A1(n1293), .A2(n1088), .ZN(n1235) );
NOR2_X1 U967 ( .A1(n1273), .A2(n1294), .ZN(n1088) );
INV_X1 U968 ( .A(n1272), .ZN(n1294) );
NAND2_X1 U969 ( .A1(n1295), .A2(n1296), .ZN(G15) );
NAND2_X1 U970 ( .A1(n1233), .A2(n1297), .ZN(n1296) );
XOR2_X1 U971 ( .A(KEYINPUT52), .B(n1298), .Z(n1295) );
NOR2_X1 U972 ( .A1(n1233), .A2(n1297), .ZN(n1298) );
AND2_X1 U973 ( .A1(n1293), .A2(n1080), .ZN(n1233) );
NOR2_X1 U974 ( .A1(n1272), .A2(n1299), .ZN(n1080) );
AND3_X1 U975 ( .A1(n1262), .A2(n1238), .A3(n1079), .ZN(n1293) );
NOR2_X1 U976 ( .A1(n1116), .A2(n1093), .ZN(n1079) );
NOR2_X1 U977 ( .A1(n1102), .A2(n1101), .ZN(n1262) );
XNOR2_X1 U978 ( .A(n1218), .B(n1232), .ZN(G12) );
AND3_X1 U979 ( .A1(n1239), .A2(n1101), .A3(n1290), .ZN(n1232) );
AND3_X1 U980 ( .A1(n1238), .A2(n1102), .A3(n1089), .ZN(n1290) );
NOR2_X1 U981 ( .A1(n1272), .A2(n1273), .ZN(n1089) );
INV_X1 U982 ( .A(n1299), .ZN(n1273) );
NOR2_X1 U983 ( .A1(n1300), .A2(n1114), .ZN(n1299) );
NOR2_X1 U984 ( .A1(n1128), .A2(G475), .ZN(n1114) );
AND2_X1 U985 ( .A1(n1301), .A2(n1128), .ZN(n1300) );
NAND2_X1 U986 ( .A1(n1187), .A2(n1302), .ZN(n1128) );
XNOR2_X1 U987 ( .A(n1303), .B(n1304), .ZN(n1187) );
XNOR2_X1 U988 ( .A(n1288), .B(n1305), .ZN(n1304) );
XNOR2_X1 U989 ( .A(n1269), .B(G131), .ZN(n1305) );
XOR2_X1 U990 ( .A(n1306), .B(n1307), .Z(n1303) );
NOR2_X1 U991 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NOR2_X1 U992 ( .A1(G104), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U993 ( .A(G125), .B(G140), .ZN(n1310) );
NOR2_X1 U994 ( .A1(n1311), .A2(n1191), .ZN(n1308) );
INV_X1 U995 ( .A(G104), .ZN(n1191) );
NOR2_X1 U996 ( .A1(n1151), .A2(n1312), .ZN(n1311) );
INV_X1 U997 ( .A(n1148), .ZN(n1312) );
XNOR2_X1 U998 ( .A(n1313), .B(n1297), .ZN(n1306) );
NAND2_X1 U999 ( .A1(KEYINPUT40), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1000 ( .A(n1315), .B(n1316), .Z(n1314) );
NOR2_X1 U1001 ( .A1(G143), .A2(KEYINPUT60), .ZN(n1316) );
AND3_X1 U1002 ( .A1(G214), .A2(n1068), .A3(n1317), .ZN(n1315) );
XNOR2_X1 U1003 ( .A(G475), .B(KEYINPUT43), .ZN(n1301) );
XNOR2_X1 U1004 ( .A(n1123), .B(n1318), .ZN(n1272) );
NOR2_X1 U1005 ( .A1(KEYINPUT48), .A2(n1181), .ZN(n1318) );
INV_X1 U1006 ( .A(G478), .ZN(n1181) );
OR2_X1 U1007 ( .A1(n1180), .A2(G902), .ZN(n1123) );
XOR2_X1 U1008 ( .A(n1319), .B(n1320), .Z(n1180) );
XOR2_X1 U1009 ( .A(n1321), .B(n1322), .Z(n1320) );
NAND2_X1 U1010 ( .A1(G217), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1011 ( .A1(KEYINPUT30), .A2(n1288), .ZN(n1321) );
XOR2_X1 U1012 ( .A(n1324), .B(n1325), .Z(n1319) );
NOR2_X1 U1013 ( .A1(KEYINPUT24), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1014 ( .A(G134), .B(n1327), .Z(n1326) );
NOR2_X1 U1015 ( .A1(KEYINPUT21), .A2(n1328), .ZN(n1327) );
XNOR2_X1 U1016 ( .A(G128), .B(G143), .ZN(n1328) );
XNOR2_X1 U1017 ( .A(G107), .B(G116), .ZN(n1324) );
XOR2_X1 U1018 ( .A(n1126), .B(n1124), .Z(n1102) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1329), .ZN(n1124) );
NAND2_X1 U1020 ( .A1(n1330), .A2(n1302), .ZN(n1126) );
XOR2_X1 U1021 ( .A(n1172), .B(KEYINPUT0), .Z(n1330) );
NAND2_X1 U1022 ( .A1(n1331), .A2(n1332), .ZN(n1172) );
NAND2_X1 U1023 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XOR2_X1 U1024 ( .A(n1335), .B(KEYINPUT6), .Z(n1331) );
OR2_X1 U1025 ( .A1(n1334), .A2(n1333), .ZN(n1335) );
XNOR2_X1 U1026 ( .A(n1336), .B(n1337), .ZN(n1333) );
XOR2_X1 U1027 ( .A(n1338), .B(n1339), .Z(n1337) );
NAND2_X1 U1028 ( .A1(KEYINPUT18), .A2(n1269), .ZN(n1339) );
NAND3_X1 U1029 ( .A1(n1340), .A2(n1341), .A3(n1148), .ZN(n1338) );
NAND2_X1 U1030 ( .A1(G125), .A2(G140), .ZN(n1148) );
NAND2_X1 U1031 ( .A1(n1342), .A2(n1151), .ZN(n1341) );
NOR2_X1 U1032 ( .A1(G125), .A2(G140), .ZN(n1151) );
INV_X1 U1033 ( .A(n1343), .ZN(n1342) );
NAND2_X1 U1034 ( .A1(n1343), .A2(G140), .ZN(n1340) );
XOR2_X1 U1035 ( .A(KEYINPUT42), .B(KEYINPUT34), .Z(n1343) );
XNOR2_X1 U1036 ( .A(G110), .B(n1344), .ZN(n1336) );
XNOR2_X1 U1037 ( .A(n1345), .B(G119), .ZN(n1344) );
INV_X1 U1038 ( .A(G128), .ZN(n1345) );
XNOR2_X1 U1039 ( .A(n1346), .B(G137), .ZN(n1334) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1323), .ZN(n1346) );
AND2_X1 U1041 ( .A1(G234), .A2(n1068), .ZN(n1323) );
NOR2_X1 U1042 ( .A1(n1104), .A2(n1244), .ZN(n1238) );
INV_X1 U1043 ( .A(n1281), .ZN(n1244) );
NAND2_X1 U1044 ( .A1(n1108), .A2(n1347), .ZN(n1281) );
NAND4_X1 U1045 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1166), .ZN(n1347) );
INV_X1 U1046 ( .A(G898), .ZN(n1166) );
NAND3_X1 U1047 ( .A1(n1287), .A2(n1068), .A3(G952), .ZN(n1108) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1287) );
INV_X1 U1049 ( .A(n1240), .ZN(n1104) );
NOR2_X1 U1050 ( .A1(n1107), .A2(n1106), .ZN(n1240) );
INV_X1 U1051 ( .A(n1277), .ZN(n1106) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1348), .ZN(n1277) );
XNOR2_X1 U1053 ( .A(n1349), .B(n1225), .ZN(n1107) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1348), .ZN(n1225) );
NAND2_X1 U1055 ( .A1(n1317), .A2(n1302), .ZN(n1348) );
NAND2_X1 U1056 ( .A1(n1350), .A2(n1302), .ZN(n1349) );
XOR2_X1 U1057 ( .A(n1351), .B(n1352), .Z(n1350) );
XOR2_X1 U1058 ( .A(KEYINPUT14), .B(n1353), .Z(n1352) );
NOR2_X1 U1059 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1353) );
XNOR2_X1 U1060 ( .A(n1221), .B(n1199), .ZN(n1351) );
INV_X1 U1061 ( .A(n1268), .ZN(n1199) );
XNOR2_X1 U1062 ( .A(n1168), .B(n1354), .ZN(n1221) );
XOR2_X1 U1063 ( .A(n1355), .B(n1169), .Z(n1354) );
XNOR2_X1 U1064 ( .A(n1218), .B(n1356), .ZN(n1169) );
XNOR2_X1 U1065 ( .A(KEYINPUT16), .B(n1288), .ZN(n1356) );
INV_X1 U1066 ( .A(G122), .ZN(n1288) );
NOR2_X1 U1067 ( .A1(G953), .A2(n1162), .ZN(n1355) );
INV_X1 U1068 ( .A(G224), .ZN(n1162) );
XNOR2_X1 U1069 ( .A(n1357), .B(n1358), .ZN(n1168) );
XNOR2_X1 U1070 ( .A(n1297), .B(n1359), .ZN(n1358) );
XNOR2_X1 U1071 ( .A(G119), .B(n1291), .ZN(n1359) );
INV_X1 U1072 ( .A(G116), .ZN(n1291) );
XNOR2_X1 U1073 ( .A(n1360), .B(n1361), .ZN(n1357) );
NAND2_X1 U1074 ( .A1(KEYINPUT45), .A2(n1362), .ZN(n1360) );
INV_X1 U1075 ( .A(n1279), .ZN(n1101) );
NAND3_X1 U1076 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1279) );
NAND2_X1 U1077 ( .A1(n1366), .A2(n1206), .ZN(n1365) );
OR3_X1 U1078 ( .A1(n1206), .A2(n1366), .A3(n1367), .ZN(n1364) );
NOR2_X1 U1079 ( .A1(KEYINPUT25), .A2(n1122), .ZN(n1366) );
INV_X1 U1080 ( .A(G472), .ZN(n1206) );
NAND2_X1 U1081 ( .A1(n1368), .A2(n1367), .ZN(n1363) );
INV_X1 U1082 ( .A(KEYINPUT59), .ZN(n1367) );
NAND2_X1 U1083 ( .A1(G472), .A2(n1122), .ZN(n1368) );
OR2_X1 U1084 ( .A1(n1121), .A2(G902), .ZN(n1122) );
XOR2_X1 U1085 ( .A(n1369), .B(n1361), .Z(n1121) );
INV_X1 U1086 ( .A(n1370), .ZN(n1361) );
XNOR2_X1 U1087 ( .A(n1371), .B(n1372), .ZN(n1369) );
NAND2_X1 U1088 ( .A1(KEYINPUT22), .A2(n1202), .ZN(n1372) );
AND3_X1 U1089 ( .A1(n1317), .A2(n1068), .A3(G210), .ZN(n1202) );
INV_X1 U1090 ( .A(G953), .ZN(n1068) );
INV_X1 U1091 ( .A(G237), .ZN(n1317) );
NAND3_X1 U1092 ( .A1(KEYINPUT28), .A2(n1373), .A3(n1374), .ZN(n1371) );
XOR2_X1 U1093 ( .A(n1375), .B(KEYINPUT46), .Z(n1374) );
NAND2_X1 U1094 ( .A1(n1376), .A2(n1205), .ZN(n1375) );
OR2_X1 U1095 ( .A1(n1205), .A2(n1376), .ZN(n1373) );
XNOR2_X1 U1096 ( .A(n1377), .B(n1378), .ZN(n1376) );
XNOR2_X1 U1097 ( .A(n1268), .B(KEYINPUT55), .ZN(n1377) );
XOR2_X1 U1098 ( .A(G128), .B(n1379), .Z(n1268) );
XNOR2_X1 U1099 ( .A(n1380), .B(n1381), .ZN(n1205) );
XNOR2_X1 U1100 ( .A(n1297), .B(n1382), .ZN(n1381) );
NOR2_X1 U1101 ( .A1(G119), .A2(KEYINPUT41), .ZN(n1382) );
INV_X1 U1102 ( .A(G113), .ZN(n1297) );
XNOR2_X1 U1103 ( .A(G116), .B(KEYINPUT54), .ZN(n1380) );
NOR2_X1 U1104 ( .A1(n1094), .A2(n1093), .ZN(n1239) );
AND2_X1 U1105 ( .A1(G221), .A2(n1329), .ZN(n1093) );
NAND2_X1 U1106 ( .A1(G234), .A2(n1302), .ZN(n1329) );
INV_X1 U1107 ( .A(n1116), .ZN(n1094) );
XOR2_X1 U1108 ( .A(n1383), .B(n1211), .Z(n1116) );
INV_X1 U1109 ( .A(G469), .ZN(n1211) );
NAND2_X1 U1110 ( .A1(n1384), .A2(n1302), .ZN(n1383) );
INV_X1 U1111 ( .A(G902), .ZN(n1302) );
XOR2_X1 U1112 ( .A(n1217), .B(n1214), .Z(n1384) );
XOR2_X1 U1113 ( .A(n1385), .B(n1386), .Z(n1214) );
XOR2_X1 U1114 ( .A(n1387), .B(n1362), .Z(n1386) );
XOR2_X1 U1115 ( .A(G107), .B(G104), .Z(n1362) );
NOR2_X1 U1116 ( .A1(G953), .A2(n1137), .ZN(n1387) );
INV_X1 U1117 ( .A(G227), .ZN(n1137) );
XOR2_X1 U1118 ( .A(n1198), .B(n1141), .Z(n1385) );
XNOR2_X1 U1119 ( .A(n1388), .B(n1389), .ZN(n1141) );
NOR2_X1 U1120 ( .A1(KEYINPUT36), .A2(n1379), .ZN(n1389) );
XNOR2_X1 U1121 ( .A(G143), .B(n1269), .ZN(n1379) );
INV_X1 U1122 ( .A(G146), .ZN(n1269) );
XNOR2_X1 U1123 ( .A(G128), .B(KEYINPUT38), .ZN(n1388) );
XNOR2_X1 U1124 ( .A(n1370), .B(n1378), .ZN(n1198) );
XNOR2_X1 U1125 ( .A(n1390), .B(n1145), .ZN(n1378) );
XOR2_X1 U1126 ( .A(G131), .B(G137), .Z(n1145) );
XNOR2_X1 U1127 ( .A(G134), .B(KEYINPUT8), .ZN(n1390) );
XOR2_X1 U1128 ( .A(G101), .B(KEYINPUT3), .Z(n1370) );
XNOR2_X1 U1129 ( .A(G110), .B(G140), .ZN(n1217) );
INV_X1 U1130 ( .A(G110), .ZN(n1218) );
endmodule


