//Key = 0000001111010111110111111101100001111110101111010110100000111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346;

XOR2_X1 U743 ( .A(G107), .B(n1012), .Z(G9) );
NOR2_X1 U744 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U745 ( .A1(G953), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1014) );
NOR2_X1 U746 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U747 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR4_X1 U748 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
NOR4_X1 U749 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1023) );
NOR2_X1 U750 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XOR2_X1 U751 ( .A(n1032), .B(KEYINPUT5), .Z(n1030) );
NOR2_X1 U752 ( .A1(n1033), .A2(n1034), .ZN(n1028) );
NOR2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U754 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U755 ( .A1(n1039), .A2(n1032), .ZN(n1027) );
NOR2_X1 U756 ( .A1(n1040), .A2(n1041), .ZN(n1022) );
NOR2_X1 U757 ( .A1(n1034), .A2(n1032), .ZN(n1040) );
NOR4_X1 U758 ( .A1(n1026), .A2(n1042), .A3(n1034), .A4(n1032), .ZN(n1020) );
NOR2_X1 U759 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U760 ( .A1(n1045), .A2(n1024), .ZN(n1044) );
NOR2_X1 U761 ( .A1(n1046), .A2(n1025), .ZN(n1043) );
INV_X1 U762 ( .A(n1047), .ZN(n1025) );
NOR2_X1 U763 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U764 ( .A1(n1015), .A2(G953), .A3(G952), .ZN(n1013) );
AND4_X1 U765 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1015) );
NOR4_X1 U766 ( .A1(n1054), .A2(n1026), .A3(n1055), .A4(n1024), .ZN(n1053) );
INV_X1 U767 ( .A(n1056), .ZN(n1024) );
NOR2_X1 U768 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
INV_X1 U769 ( .A(n1041), .ZN(n1026) );
NOR3_X1 U770 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1052) );
NOR2_X1 U771 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U772 ( .A(KEYINPUT9), .ZN(n1063) );
NOR2_X1 U773 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
AND3_X1 U774 ( .A1(KEYINPUT60), .A2(n1058), .A3(n1057), .ZN(n1065) );
NOR2_X1 U775 ( .A1(KEYINPUT60), .A2(n1057), .ZN(n1064) );
NOR2_X1 U776 ( .A1(KEYINPUT9), .A2(n1066), .ZN(n1060) );
NOR2_X1 U777 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U778 ( .A(KEYINPUT60), .B(n1057), .Z(n1068) );
INV_X1 U779 ( .A(n1058), .ZN(n1067) );
XOR2_X1 U780 ( .A(G469), .B(n1069), .Z(n1059) );
NAND2_X1 U781 ( .A1(KEYINPUT62), .A2(n1034), .ZN(n1051) );
INV_X1 U782 ( .A(n1070), .ZN(n1034) );
NAND2_X1 U783 ( .A1(n1071), .A2(n1072), .ZN(n1050) );
INV_X1 U784 ( .A(KEYINPUT62), .ZN(n1072) );
OR2_X1 U785 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
XOR2_X1 U786 ( .A(n1075), .B(n1076), .Z(G72) );
XOR2_X1 U787 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U788 ( .A1(G953), .A2(n1079), .ZN(n1078) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1079) );
NAND3_X1 U790 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
NAND2_X1 U791 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U792 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U793 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U794 ( .A1(n1088), .A2(KEYINPUT12), .ZN(n1087) );
NAND3_X1 U795 ( .A1(n1089), .A2(n1090), .A3(n1088), .ZN(n1080) );
INV_X1 U796 ( .A(KEYINPUT55), .ZN(n1088) );
NAND2_X1 U797 ( .A1(n1086), .A2(n1091), .ZN(n1090) );
OR2_X1 U798 ( .A1(n1084), .A2(KEYINPUT12), .ZN(n1091) );
XNOR2_X1 U799 ( .A(n1092), .B(n1093), .ZN(n1084) );
NOR2_X1 U800 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND3_X1 U801 ( .A1(KEYINPUT57), .A2(n1096), .A3(G131), .ZN(n1095) );
NOR2_X1 U802 ( .A1(KEYINPUT57), .A2(n1097), .ZN(n1094) );
XOR2_X1 U803 ( .A(n1098), .B(KEYINPUT58), .Z(n1092) );
OR2_X1 U804 ( .A1(n1086), .A2(KEYINPUT12), .ZN(n1089) );
XOR2_X1 U805 ( .A(n1099), .B(n1100), .Z(n1086) );
NOR2_X1 U806 ( .A1(n1101), .A2(G953), .ZN(n1075) );
XOR2_X1 U807 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U808 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND3_X1 U809 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
XOR2_X1 U810 ( .A(n1109), .B(KEYINPUT51), .Z(n1108) );
OR2_X1 U811 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U812 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NAND2_X1 U813 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND2_X1 U814 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U815 ( .A(KEYINPUT6), .B(n1116), .Z(n1114) );
NAND2_X1 U816 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
XOR2_X1 U817 ( .A(n1119), .B(KEYINPUT37), .Z(n1118) );
INV_X1 U818 ( .A(n1115), .ZN(n1117) );
NAND2_X1 U819 ( .A1(G953), .A2(n1120), .ZN(n1106) );
NAND2_X1 U820 ( .A1(n1121), .A2(n1122), .ZN(n1104) );
XOR2_X1 U821 ( .A(KEYINPUT49), .B(G953), .Z(n1121) );
NOR2_X1 U822 ( .A1(n1123), .A2(n1124), .ZN(n1102) );
NOR2_X1 U823 ( .A1(n1125), .A2(n1120), .ZN(n1123) );
NOR2_X1 U824 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U825 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND4_X1 U826 ( .A1(KEYINPUT47), .A2(n1130), .A3(G217), .A4(n1131), .ZN(n1128) );
NOR2_X1 U827 ( .A1(n1126), .A2(n1132), .ZN(G63) );
XNOR2_X1 U828 ( .A(n1133), .B(n1134), .ZN(n1132) );
AND2_X1 U829 ( .A1(G478), .A2(n1130), .ZN(n1134) );
NOR2_X1 U830 ( .A1(n1126), .A2(n1135), .ZN(G60) );
XOR2_X1 U831 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U832 ( .A1(KEYINPUT24), .A2(n1138), .ZN(n1136) );
NAND2_X1 U833 ( .A1(n1130), .A2(G475), .ZN(n1138) );
XOR2_X1 U834 ( .A(G104), .B(n1139), .Z(G6) );
NOR2_X1 U835 ( .A1(n1126), .A2(n1140), .ZN(G57) );
XOR2_X1 U836 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U837 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U838 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U839 ( .A1(G472), .A2(n1130), .ZN(n1146) );
NAND2_X1 U840 ( .A1(n1147), .A2(KEYINPUT25), .ZN(n1145) );
XOR2_X1 U841 ( .A(n1148), .B(KEYINPUT10), .Z(n1147) );
XNOR2_X1 U842 ( .A(n1149), .B(n1150), .ZN(n1141) );
XOR2_X1 U843 ( .A(KEYINPUT54), .B(G101), .Z(n1150) );
NOR2_X1 U844 ( .A1(n1126), .A2(n1151), .ZN(G54) );
XOR2_X1 U845 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U846 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U847 ( .A(n1156), .B(n1157), .Z(n1152) );
XOR2_X1 U848 ( .A(KEYINPUT61), .B(n1158), .Z(n1157) );
AND2_X1 U849 ( .A1(G469), .A2(n1130), .ZN(n1158) );
NOR2_X1 U850 ( .A1(n1126), .A2(n1159), .ZN(G51) );
XOR2_X1 U851 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR3_X1 U852 ( .A1(n1162), .A2(KEYINPUT46), .A3(n1163), .ZN(n1161) );
NOR2_X1 U853 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U854 ( .A(KEYINPUT41), .B(n1166), .Z(n1165) );
NOR2_X1 U855 ( .A1(n1167), .A2(n1166), .ZN(n1164) );
NOR2_X1 U856 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U857 ( .A1(n1170), .A2(n1171), .ZN(n1162) );
NOR2_X1 U858 ( .A1(n1166), .A2(n1169), .ZN(n1170) );
INV_X1 U859 ( .A(KEYINPUT11), .ZN(n1169) );
AND3_X1 U860 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1166) );
NAND2_X1 U861 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
INV_X1 U862 ( .A(KEYINPUT29), .ZN(n1176) );
NAND2_X1 U863 ( .A1(KEYINPUT29), .A2(n1177), .ZN(n1172) );
NAND2_X1 U864 ( .A1(n1130), .A2(n1057), .ZN(n1160) );
INV_X1 U865 ( .A(n1178), .ZN(n1057) );
AND2_X1 U866 ( .A1(n1179), .A2(n1017), .ZN(n1130) );
NAND2_X1 U867 ( .A1(n1101), .A2(n1180), .ZN(n1017) );
INV_X1 U868 ( .A(n1122), .ZN(n1180) );
NAND4_X1 U869 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1122) );
NOR4_X1 U870 ( .A1(n1012), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
INV_X1 U871 ( .A(n1188), .ZN(n1186) );
AND2_X1 U872 ( .A1(n1048), .A2(n1189), .ZN(n1012) );
NOR3_X1 U873 ( .A1(n1139), .A2(n1190), .A3(n1191), .ZN(n1183) );
NOR2_X1 U874 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
INV_X1 U875 ( .A(KEYINPUT20), .ZN(n1192) );
NOR3_X1 U876 ( .A1(KEYINPUT20), .A2(n1194), .A3(n1195), .ZN(n1190) );
AND2_X1 U877 ( .A1(n1049), .A2(n1189), .ZN(n1139) );
AND3_X1 U878 ( .A1(n1036), .A2(n1070), .A3(n1196), .ZN(n1189) );
AND4_X1 U879 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1101) );
NOR4_X1 U880 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR3_X1 U881 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1204) );
XOR2_X1 U882 ( .A(KEYINPUT35), .B(n1208), .Z(n1205) );
INV_X1 U883 ( .A(n1209), .ZN(n1202) );
INV_X1 U884 ( .A(n1210), .ZN(n1201) );
NOR2_X1 U885 ( .A1(n1211), .A2(n1212), .ZN(n1199) );
XOR2_X1 U886 ( .A(n1213), .B(KEYINPUT34), .Z(n1179) );
NOR2_X1 U887 ( .A1(n1124), .A2(G952), .ZN(n1126) );
XOR2_X1 U888 ( .A(n1214), .B(n1210), .Z(G48) );
NAND3_X1 U889 ( .A1(n1215), .A2(n1216), .A3(n1049), .ZN(n1210) );
XNOR2_X1 U890 ( .A(G143), .B(n1197), .ZN(G45) );
NAND4_X1 U891 ( .A1(n1215), .A2(n1208), .A3(n1217), .A4(n1218), .ZN(n1197) );
XOR2_X1 U892 ( .A(n1203), .B(n1219), .Z(G42) );
NOR2_X1 U893 ( .A1(KEYINPUT4), .A2(n1100), .ZN(n1219) );
NOR3_X1 U894 ( .A1(n1220), .A2(n1207), .A3(n1031), .ZN(n1203) );
XNOR2_X1 U895 ( .A(G137), .B(n1198), .ZN(G39) );
NAND3_X1 U896 ( .A1(n1056), .A2(n1216), .A3(n1221), .ZN(n1198) );
XOR2_X1 U897 ( .A(G134), .B(n1222), .Z(G36) );
AND2_X1 U898 ( .A1(n1221), .A2(n1223), .ZN(n1222) );
XOR2_X1 U899 ( .A(G131), .B(n1212), .Z(G33) );
NOR3_X1 U900 ( .A1(n1207), .A2(n1039), .A3(n1220), .ZN(n1212) );
INV_X1 U901 ( .A(n1221), .ZN(n1207) );
NOR3_X1 U902 ( .A1(n1045), .A2(n1224), .A3(n1032), .ZN(n1221) );
OR2_X1 U903 ( .A1(n1038), .A2(n1225), .ZN(n1032) );
XOR2_X1 U904 ( .A(KEYINPUT36), .B(n1037), .Z(n1225) );
XOR2_X1 U905 ( .A(G128), .B(n1211), .Z(G30) );
AND3_X1 U906 ( .A1(n1048), .A2(n1216), .A3(n1215), .ZN(n1211) );
NOR3_X1 U907 ( .A1(n1045), .A2(n1195), .A3(n1224), .ZN(n1215) );
INV_X1 U908 ( .A(n1226), .ZN(n1045) );
XOR2_X1 U909 ( .A(n1227), .B(n1228), .Z(G3) );
NAND2_X1 U910 ( .A1(KEYINPUT23), .A2(n1229), .ZN(n1228) );
INV_X1 U911 ( .A(n1181), .ZN(n1229) );
NAND4_X1 U912 ( .A1(n1208), .A2(n1056), .A3(n1196), .A4(n1036), .ZN(n1181) );
XOR2_X1 U913 ( .A(n1099), .B(n1209), .Z(G27) );
NAND3_X1 U914 ( .A1(n1047), .A2(n1230), .A3(n1231), .ZN(n1209) );
NOR3_X1 U915 ( .A1(n1220), .A2(n1195), .A3(n1224), .ZN(n1231) );
NAND2_X1 U916 ( .A1(n1041), .A2(n1232), .ZN(n1224) );
NAND2_X1 U917 ( .A1(n1019), .A2(n1233), .ZN(n1232) );
NAND3_X1 U918 ( .A1(G953), .A2(n1083), .A3(n1234), .ZN(n1233) );
INV_X1 U919 ( .A(G900), .ZN(n1083) );
NAND2_X1 U920 ( .A1(n1235), .A2(n1236), .ZN(G24) );
NAND2_X1 U921 ( .A1(G122), .A2(n1182), .ZN(n1236) );
XOR2_X1 U922 ( .A(KEYINPUT16), .B(n1237), .Z(n1235) );
NOR2_X1 U923 ( .A1(G122), .A2(n1182), .ZN(n1237) );
NAND4_X1 U924 ( .A1(n1238), .A2(n1070), .A3(n1217), .A4(n1218), .ZN(n1182) );
NOR2_X1 U925 ( .A1(n1239), .A2(n1073), .ZN(n1070) );
XOR2_X1 U926 ( .A(G119), .B(n1187), .Z(G21) );
AND3_X1 U927 ( .A1(n1056), .A2(n1216), .A3(n1238), .ZN(n1187) );
NAND2_X1 U928 ( .A1(n1240), .A2(n1241), .ZN(n1216) );
NAND3_X1 U929 ( .A1(n1073), .A2(n1239), .A3(n1242), .ZN(n1241) );
INV_X1 U930 ( .A(KEYINPUT53), .ZN(n1242) );
NAND2_X1 U931 ( .A1(KEYINPUT53), .A2(n1208), .ZN(n1240) );
NAND2_X1 U932 ( .A1(n1243), .A2(n1244), .ZN(G18) );
NAND2_X1 U933 ( .A1(G116), .A2(n1188), .ZN(n1244) );
XOR2_X1 U934 ( .A(KEYINPUT13), .B(n1245), .Z(n1243) );
NOR2_X1 U935 ( .A1(G116), .A2(n1188), .ZN(n1245) );
NAND2_X1 U936 ( .A1(n1223), .A2(n1238), .ZN(n1188) );
NOR2_X1 U937 ( .A1(n1039), .A2(n1206), .ZN(n1223) );
INV_X1 U938 ( .A(n1048), .ZN(n1206) );
NOR2_X1 U939 ( .A1(n1218), .A2(n1246), .ZN(n1048) );
XOR2_X1 U940 ( .A(G113), .B(n1185), .Z(G15) );
AND3_X1 U941 ( .A1(n1049), .A2(n1208), .A3(n1238), .ZN(n1185) );
AND4_X1 U942 ( .A1(n1047), .A2(n1036), .A3(n1247), .A4(n1041), .ZN(n1238) );
XOR2_X1 U943 ( .A(n1226), .B(KEYINPUT59), .Z(n1047) );
INV_X1 U944 ( .A(n1039), .ZN(n1208) );
NAND2_X1 U945 ( .A1(n1074), .A2(n1073), .ZN(n1039) );
INV_X1 U946 ( .A(n1239), .ZN(n1074) );
INV_X1 U947 ( .A(n1220), .ZN(n1049) );
NAND2_X1 U948 ( .A1(n1246), .A2(n1218), .ZN(n1220) );
XOR2_X1 U949 ( .A(n1193), .B(n1248), .Z(G12) );
NOR2_X1 U950 ( .A1(G110), .A2(KEYINPUT1), .ZN(n1248) );
NAND2_X1 U951 ( .A1(n1194), .A2(n1036), .ZN(n1193) );
INV_X1 U952 ( .A(n1195), .ZN(n1036) );
NAND2_X1 U953 ( .A1(n1249), .A2(n1038), .ZN(n1195) );
XOR2_X1 U954 ( .A(n1058), .B(n1178), .Z(n1038) );
NAND2_X1 U955 ( .A1(G210), .A2(n1250), .ZN(n1178) );
NAND2_X1 U956 ( .A1(n1251), .A2(n1213), .ZN(n1058) );
XOR2_X1 U957 ( .A(n1252), .B(n1168), .Z(n1251) );
INV_X1 U958 ( .A(n1171), .ZN(n1168) );
XOR2_X1 U959 ( .A(n1253), .B(n1111), .Z(n1171) );
XOR2_X1 U960 ( .A(G110), .B(G122), .Z(n1111) );
NAND2_X1 U961 ( .A1(n1254), .A2(KEYINPUT40), .ZN(n1253) );
XOR2_X1 U962 ( .A(n1115), .B(n1255), .Z(n1254) );
XOR2_X1 U963 ( .A(KEYINPUT18), .B(n1116), .Z(n1255) );
INV_X1 U964 ( .A(n1119), .ZN(n1116) );
XNOR2_X1 U965 ( .A(G113), .B(n1256), .ZN(n1119) );
NOR2_X1 U966 ( .A1(KEYINPUT32), .A2(n1257), .ZN(n1256) );
XOR2_X1 U967 ( .A(G116), .B(n1258), .Z(n1257) );
XOR2_X1 U968 ( .A(KEYINPUT17), .B(G119), .Z(n1258) );
XOR2_X1 U969 ( .A(n1227), .B(n1259), .Z(n1115) );
INV_X1 U970 ( .A(G101), .ZN(n1227) );
NOR2_X1 U971 ( .A1(n1175), .A2(n1260), .ZN(n1252) );
INV_X1 U972 ( .A(n1174), .ZN(n1260) );
NAND2_X1 U973 ( .A1(n1177), .A2(n1261), .ZN(n1174) );
NAND2_X1 U974 ( .A1(G224), .A2(n1124), .ZN(n1261) );
NOR3_X1 U975 ( .A1(n1177), .A2(G953), .A3(n1125), .ZN(n1175) );
INV_X1 U976 ( .A(G224), .ZN(n1125) );
XNOR2_X1 U977 ( .A(n1148), .B(n1099), .ZN(n1177) );
XOR2_X1 U978 ( .A(KEYINPUT36), .B(n1054), .Z(n1249) );
INV_X1 U979 ( .A(n1037), .ZN(n1054) );
NAND2_X1 U980 ( .A1(G214), .A2(n1250), .ZN(n1037) );
NAND2_X1 U981 ( .A1(n1262), .A2(n1213), .ZN(n1250) );
AND3_X1 U982 ( .A1(n1056), .A2(n1196), .A3(n1230), .ZN(n1194) );
INV_X1 U983 ( .A(n1031), .ZN(n1230) );
NAND2_X1 U984 ( .A1(n1263), .A2(n1264), .ZN(n1031) );
XOR2_X1 U985 ( .A(KEYINPUT33), .B(n1073), .Z(n1264) );
XNOR2_X1 U986 ( .A(n1265), .B(G472), .ZN(n1073) );
NAND2_X1 U987 ( .A1(n1266), .A2(n1213), .ZN(n1265) );
XOR2_X1 U988 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U989 ( .A(n1269), .B(G101), .Z(n1268) );
NAND2_X1 U990 ( .A1(KEYINPUT7), .A2(n1270), .ZN(n1269) );
XOR2_X1 U991 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U992 ( .A(n1273), .B(KEYINPUT63), .ZN(n1272) );
NAND2_X1 U993 ( .A1(KEYINPUT52), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U994 ( .A(KEYINPUT10), .B(n1148), .ZN(n1274) );
XOR2_X1 U995 ( .A(n1275), .B(n1276), .Z(n1148) );
NAND2_X1 U996 ( .A1(KEYINPUT21), .A2(n1277), .ZN(n1275) );
XOR2_X1 U997 ( .A(G146), .B(G143), .Z(n1277) );
INV_X1 U998 ( .A(n1143), .ZN(n1271) );
XOR2_X1 U999 ( .A(n1097), .B(n1278), .Z(n1143) );
XNOR2_X1 U1000 ( .A(G113), .B(n1279), .ZN(n1278) );
NAND2_X1 U1001 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U1002 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U1003 ( .A(KEYINPUT44), .B(G116), .Z(n1283) );
XOR2_X1 U1004 ( .A(n1284), .B(KEYINPUT56), .Z(n1282) );
NAND2_X1 U1005 ( .A1(n1285), .A2(n1286), .ZN(n1280) );
XOR2_X1 U1006 ( .A(KEYINPUT26), .B(G119), .Z(n1286) );
XOR2_X1 U1007 ( .A(KEYINPUT44), .B(n1287), .Z(n1285) );
INV_X1 U1008 ( .A(n1156), .ZN(n1097) );
NAND2_X1 U1009 ( .A1(KEYINPUT15), .A2(n1149), .ZN(n1267) );
AND3_X1 U1010 ( .A1(n1262), .A2(n1124), .A3(G210), .ZN(n1149) );
XOR2_X1 U1011 ( .A(n1239), .B(KEYINPUT53), .Z(n1263) );
NAND3_X1 U1012 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1239) );
OR2_X1 U1013 ( .A1(n1291), .A2(n1129), .ZN(n1290) );
NAND3_X1 U1014 ( .A1(n1129), .A2(n1291), .A3(n1213), .ZN(n1289) );
NAND2_X1 U1015 ( .A1(G217), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1016 ( .A(n1293), .B(n1294), .Z(n1129) );
XOR2_X1 U1017 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1018 ( .A(G125), .B(G110), .Z(n1296) );
XOR2_X1 U1019 ( .A(KEYINPUT50), .B(G137), .Z(n1295) );
XNOR2_X1 U1020 ( .A(n1297), .B(n1298), .ZN(n1293) );
XOR2_X1 U1021 ( .A(n1299), .B(n1300), .Z(n1298) );
NAND2_X1 U1022 ( .A1(G221), .A2(n1301), .ZN(n1300) );
NAND2_X1 U1023 ( .A1(n1302), .A2(n1303), .ZN(n1299) );
NAND2_X1 U1024 ( .A1(G119), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1025 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1026 ( .A1(G128), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1027 ( .A1(n1308), .A2(n1309), .ZN(n1302) );
INV_X1 U1028 ( .A(G128), .ZN(n1309) );
NAND2_X1 U1029 ( .A1(n1307), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1030 ( .A1(n1284), .A2(n1305), .ZN(n1310) );
INV_X1 U1031 ( .A(KEYINPUT39), .ZN(n1305) );
INV_X1 U1032 ( .A(G119), .ZN(n1284) );
INV_X1 U1033 ( .A(KEYINPUT2), .ZN(n1307) );
NAND2_X1 U1034 ( .A1(G902), .A2(G217), .ZN(n1288) );
AND3_X1 U1035 ( .A1(n1247), .A2(n1041), .A3(n1226), .ZN(n1196) );
XOR2_X1 U1036 ( .A(n1311), .B(G469), .Z(n1226) );
NAND2_X1 U1037 ( .A1(n1312), .A2(KEYINPUT27), .ZN(n1311) );
XNOR2_X1 U1038 ( .A(n1069), .B(KEYINPUT30), .ZN(n1312) );
AND2_X1 U1039 ( .A1(n1313), .A2(n1213), .ZN(n1069) );
XNOR2_X1 U1040 ( .A(n1154), .B(n1314), .ZN(n1313) );
NOR2_X1 U1041 ( .A1(KEYINPUT31), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1042 ( .A(n1156), .B(n1316), .Z(n1315) );
XNOR2_X1 U1043 ( .A(n1317), .B(KEYINPUT8), .ZN(n1316) );
NAND2_X1 U1044 ( .A1(KEYINPUT43), .A2(n1155), .ZN(n1317) );
XNOR2_X1 U1045 ( .A(n1098), .B(n1318), .ZN(n1155) );
XOR2_X1 U1046 ( .A(n1319), .B(n1259), .Z(n1318) );
XOR2_X1 U1047 ( .A(G104), .B(G107), .Z(n1259) );
NOR2_X1 U1048 ( .A1(G101), .A2(KEYINPUT0), .ZN(n1319) );
XOR2_X1 U1049 ( .A(n1320), .B(n1276), .Z(n1098) );
XOR2_X1 U1050 ( .A(G128), .B(KEYINPUT45), .Z(n1276) );
XOR2_X1 U1051 ( .A(n1321), .B(G143), .Z(n1320) );
NAND2_X1 U1052 ( .A1(KEYINPUT38), .A2(n1214), .ZN(n1321) );
INV_X1 U1053 ( .A(G146), .ZN(n1214) );
XOR2_X1 U1054 ( .A(G131), .B(n1096), .Z(n1156) );
XOR2_X1 U1055 ( .A(G134), .B(G137), .Z(n1096) );
XNOR2_X1 U1056 ( .A(n1322), .B(n1323), .ZN(n1154) );
XOR2_X1 U1057 ( .A(G140), .B(G110), .Z(n1323) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1124), .ZN(n1322) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1131), .ZN(n1041) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1213), .ZN(n1131) );
NAND2_X1 U1061 ( .A1(n1019), .A2(n1324), .ZN(n1247) );
NAND3_X1 U1062 ( .A1(n1234), .A2(n1120), .A3(n1325), .ZN(n1324) );
XOR2_X1 U1063 ( .A(n1124), .B(KEYINPUT28), .Z(n1325) );
INV_X1 U1064 ( .A(G898), .ZN(n1120) );
AND2_X1 U1065 ( .A1(n1326), .A2(n1327), .ZN(n1234) );
XOR2_X1 U1066 ( .A(KEYINPUT3), .B(G902), .Z(n1326) );
NAND3_X1 U1067 ( .A1(n1327), .A2(n1124), .A3(G952), .ZN(n1019) );
NAND2_X1 U1068 ( .A1(G237), .A2(G234), .ZN(n1327) );
NOR2_X1 U1069 ( .A1(n1217), .A2(n1218), .ZN(n1056) );
XNOR2_X1 U1070 ( .A(n1328), .B(G475), .ZN(n1218) );
OR2_X1 U1071 ( .A1(n1137), .A2(G902), .ZN(n1328) );
XNOR2_X1 U1072 ( .A(n1329), .B(n1330), .ZN(n1137) );
XOR2_X1 U1073 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1074 ( .A(n1333), .B(G104), .Z(n1332) );
NAND2_X1 U1075 ( .A1(KEYINPUT19), .A2(n1099), .ZN(n1333) );
INV_X1 U1076 ( .A(G125), .ZN(n1099) );
XNOR2_X1 U1077 ( .A(G113), .B(G131), .ZN(n1331) );
XNOR2_X1 U1078 ( .A(n1334), .B(n1335), .ZN(n1329) );
XOR2_X1 U1079 ( .A(n1336), .B(n1297), .Z(n1335) );
XNOR2_X1 U1080 ( .A(n1100), .B(G146), .ZN(n1297) );
INV_X1 U1081 ( .A(G140), .ZN(n1100) );
AND3_X1 U1082 ( .A1(G214), .A2(n1124), .A3(n1262), .ZN(n1336) );
INV_X1 U1083 ( .A(G237), .ZN(n1262) );
INV_X1 U1084 ( .A(G953), .ZN(n1124) );
INV_X1 U1085 ( .A(n1246), .ZN(n1217) );
XOR2_X1 U1086 ( .A(n1337), .B(G478), .Z(n1246) );
NAND2_X1 U1087 ( .A1(n1133), .A2(n1213), .ZN(n1337) );
INV_X1 U1088 ( .A(G902), .ZN(n1213) );
XNOR2_X1 U1089 ( .A(n1338), .B(n1339), .ZN(n1133) );
XOR2_X1 U1090 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1091 ( .A(G134), .B(G128), .Z(n1341) );
XOR2_X1 U1092 ( .A(KEYINPUT48), .B(KEYINPUT42), .Z(n1340) );
XOR2_X1 U1093 ( .A(n1342), .B(n1343), .Z(n1338) );
XNOR2_X1 U1094 ( .A(G107), .B(n1344), .ZN(n1343) );
NAND2_X1 U1095 ( .A1(n1345), .A2(n1287), .ZN(n1344) );
INV_X1 U1096 ( .A(G116), .ZN(n1287) );
XNOR2_X1 U1097 ( .A(KEYINPUT22), .B(KEYINPUT14), .ZN(n1345) );
XOR2_X1 U1098 ( .A(n1346), .B(n1334), .Z(n1342) );
XOR2_X1 U1099 ( .A(G122), .B(G143), .Z(n1334) );
NAND2_X1 U1100 ( .A1(G217), .A2(n1301), .ZN(n1346) );
NOR2_X1 U1101 ( .A1(n1292), .A2(G953), .ZN(n1301) );
INV_X1 U1102 ( .A(G234), .ZN(n1292) );
endmodule


