//Key = 1010111111011010000000011000010111000100101001101110100010111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366;

XNOR2_X1 U740 ( .A(G107), .B(n1026), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(G75) );
AND3_X1 U742 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR3_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR4_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1041), .A2(KEYINPUT60), .ZN(n1040) );
NOR3_X1 U747 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR3_X1 U748 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1039) );
NOR3_X1 U749 ( .A1(n1043), .A2(n1047), .A3(n1048), .ZN(n1046) );
AND2_X1 U750 ( .A1(n1049), .A2(KEYINPUT49), .ZN(n1048) );
NOR3_X1 U751 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
XOR2_X1 U752 ( .A(KEYINPUT20), .B(n1053), .Z(n1050) );
NOR2_X1 U753 ( .A1(n1054), .A2(n1055), .ZN(n1045) );
NOR2_X1 U754 ( .A1(KEYINPUT49), .A2(n1056), .ZN(n1055) );
INV_X1 U755 ( .A(n1049), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1038) );
INV_X1 U757 ( .A(n1059), .ZN(n1058) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
NOR3_X1 U759 ( .A1(n1044), .A2(n1062), .A3(n1043), .ZN(n1037) );
INV_X1 U760 ( .A(n1054), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U762 ( .A1(n1065), .A2(n1051), .ZN(n1064) );
AND2_X1 U763 ( .A1(n1066), .A2(KEYINPUT60), .ZN(n1063) );
NAND3_X1 U764 ( .A1(n1067), .A2(n1030), .A3(n1029), .ZN(n1032) );
NAND4_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1029) );
NOR4_X1 U766 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
AND2_X1 U767 ( .A1(n1076), .A2(G475), .ZN(n1073) );
NOR3_X1 U768 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1070) );
NOR2_X1 U769 ( .A1(KEYINPUT10), .A2(n1080), .ZN(n1079) );
NOR2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
AND2_X1 U771 ( .A1(G475), .A2(KEYINPUT63), .ZN(n1082) );
NOR3_X1 U772 ( .A1(KEYINPUT63), .A2(G475), .A3(n1076), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
INV_X1 U774 ( .A(KEYINPUT10), .ZN(n1084) );
NOR2_X1 U775 ( .A1(n1076), .A2(n1085), .ZN(n1083) );
XOR2_X1 U776 ( .A(KEYINPUT63), .B(G475), .Z(n1085) );
XNOR2_X1 U777 ( .A(n1086), .B(KEYINPUT29), .ZN(n1076) );
XNOR2_X1 U778 ( .A(n1087), .B(n1088), .ZN(n1077) );
XNOR2_X1 U779 ( .A(G478), .B(n1089), .ZN(n1069) );
XNOR2_X1 U780 ( .A(n1090), .B(KEYINPUT7), .ZN(n1068) );
NAND3_X1 U781 ( .A1(n1054), .A2(n1091), .A3(n1059), .ZN(n1067) );
NOR3_X1 U782 ( .A1(n1074), .A2(n1044), .A3(n1051), .ZN(n1059) );
INV_X1 U783 ( .A(n1092), .ZN(n1051) );
NAND2_X1 U784 ( .A1(KEYINPUT4), .A2(n1093), .ZN(n1044) );
NAND2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1072), .A2(n1096), .ZN(n1095) );
XOR2_X1 U787 ( .A(n1097), .B(n1098), .Z(G72) );
NOR3_X1 U788 ( .A1(KEYINPUT19), .A2(n1099), .A3(n1100), .ZN(n1098) );
AND3_X1 U789 ( .A1(n1101), .A2(n1030), .A3(n1102), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1103), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1030), .A2(n1106), .ZN(n1105) );
NOR2_X1 U793 ( .A1(G953), .A2(n1102), .ZN(n1104) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(n1101) );
XOR2_X1 U795 ( .A(n1109), .B(n1110), .Z(n1107) );
NAND2_X1 U796 ( .A1(KEYINPUT31), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U797 ( .A(n1112), .B(G125), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1097) );
NAND2_X1 U799 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U802 ( .A(n1119), .B(KEYINPUT17), .Z(n1115) );
OR2_X1 U803 ( .A1(n1118), .A2(n1117), .ZN(n1119) );
NAND2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
NAND2_X1 U805 ( .A1(n1122), .A2(n1030), .ZN(n1121) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1122) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND3_X1 U808 ( .A1(G898), .A2(n1123), .A3(G953), .ZN(n1120) );
NAND2_X1 U809 ( .A1(n1113), .A2(n1127), .ZN(n1118) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1127) );
XNOR2_X1 U811 ( .A(n1030), .B(KEYINPUT18), .ZN(n1113) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U813 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND3_X1 U814 ( .A1(G217), .A2(n1132), .A3(G902), .ZN(n1130) );
XNOR2_X1 U815 ( .A(KEYINPUT52), .B(n1034), .ZN(n1132) );
INV_X1 U816 ( .A(n1133), .ZN(n1034) );
NOR2_X1 U817 ( .A1(n1128), .A2(n1134), .ZN(G63) );
NOR3_X1 U818 ( .A1(n1089), .A2(n1135), .A3(n1136), .ZN(n1134) );
AND3_X1 U819 ( .A1(n1137), .A2(G478), .A3(n1138), .ZN(n1136) );
NOR2_X1 U820 ( .A1(n1139), .A2(n1137), .ZN(n1135) );
NOR2_X1 U821 ( .A1(n1133), .A2(n1140), .ZN(n1139) );
NOR2_X1 U822 ( .A1(n1128), .A2(n1141), .ZN(G60) );
XNOR2_X1 U823 ( .A(n1142), .B(n1143), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1144), .B(KEYINPUT12), .Z(n1143) );
NAND2_X1 U825 ( .A1(n1138), .A2(G475), .ZN(n1144) );
XNOR2_X1 U826 ( .A(G104), .B(n1145), .ZN(G6) );
NOR2_X1 U827 ( .A1(n1128), .A2(n1146), .ZN(G57) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U829 ( .A(G101), .B(n1149), .ZN(n1148) );
NOR2_X1 U830 ( .A1(KEYINPUT16), .A2(n1150), .ZN(n1149) );
XOR2_X1 U831 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U832 ( .A1(n1138), .A2(G472), .ZN(n1151) );
NAND2_X1 U833 ( .A1(KEYINPUT59), .A2(n1153), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1128), .A2(n1154), .ZN(G54) );
XOR2_X1 U835 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U837 ( .A(n1112), .B(G110), .ZN(n1158) );
XOR2_X1 U838 ( .A(n1159), .B(n1110), .Z(n1155) );
XOR2_X1 U839 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U840 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U841 ( .A(n1164), .B(KEYINPUT6), .Z(n1163) );
NAND2_X1 U842 ( .A1(n1165), .A2(n1108), .ZN(n1164) );
NOR2_X1 U843 ( .A1(n1165), .A2(n1108), .ZN(n1162) );
NAND2_X1 U844 ( .A1(n1138), .A2(G469), .ZN(n1160) );
NOR2_X1 U845 ( .A1(n1128), .A2(n1166), .ZN(G51) );
XOR2_X1 U846 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U847 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1169) );
NAND2_X1 U849 ( .A1(n1138), .A2(n1087), .ZN(n1171) );
NOR2_X1 U850 ( .A1(n1173), .A2(n1133), .ZN(n1138) );
NOR3_X1 U851 ( .A1(n1126), .A2(n1174), .A3(n1102), .ZN(n1133) );
NAND2_X1 U852 ( .A1(n1175), .A2(n1176), .ZN(n1102) );
AND4_X1 U853 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR4_X1 U854 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1175) );
NOR2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U856 ( .A(KEYINPUT8), .ZN(n1186) );
NOR3_X1 U857 ( .A1(n1065), .A2(n1187), .A3(n1188), .ZN(n1182) );
NOR2_X1 U858 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR2_X1 U859 ( .A1(KEYINPUT8), .A2(n1191), .ZN(n1189) );
AND2_X1 U860 ( .A1(n1190), .A2(n1192), .ZN(n1187) );
XOR2_X1 U861 ( .A(KEYINPUT39), .B(n1125), .Z(n1174) );
NAND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1125) );
NOR2_X1 U863 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U864 ( .A1(n1199), .A2(n1200), .ZN(n1194) );
INV_X1 U865 ( .A(KEYINPUT15), .ZN(n1200) );
NAND4_X1 U866 ( .A1(n1049), .A2(n1201), .A3(n1202), .A4(KEYINPUT15), .ZN(n1193) );
AND2_X1 U867 ( .A1(n1203), .A2(n1061), .ZN(n1202) );
NAND4_X1 U868 ( .A1(n1204), .A2(n1145), .A3(n1205), .A4(n1026), .ZN(n1126) );
NAND3_X1 U869 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1026) );
NAND4_X1 U870 ( .A1(n1209), .A2(n1208), .A3(n1054), .A4(n1210), .ZN(n1145) );
OR3_X1 U871 ( .A1(n1075), .A2(n1065), .A3(n1211), .ZN(n1204) );
XOR2_X1 U872 ( .A(n1212), .B(n1213), .Z(n1167) );
NOR2_X1 U873 ( .A1(KEYINPUT43), .A2(n1214), .ZN(n1213) );
XNOR2_X1 U874 ( .A(n1215), .B(KEYINPUT21), .ZN(n1212) );
AND2_X1 U875 ( .A1(n1216), .A2(n1031), .ZN(n1128) );
INV_X1 U876 ( .A(G952), .ZN(n1031) );
XNOR2_X1 U877 ( .A(KEYINPUT62), .B(n1030), .ZN(n1216) );
XOR2_X1 U878 ( .A(G146), .B(n1181), .Z(G48) );
AND2_X1 U879 ( .A1(n1217), .A2(n1209), .ZN(n1181) );
XOR2_X1 U880 ( .A(n1185), .B(n1218), .Z(G45) );
NOR2_X1 U881 ( .A1(G143), .A2(KEYINPUT3), .ZN(n1218) );
NAND2_X1 U882 ( .A1(n1219), .A2(n1220), .ZN(n1185) );
INV_X1 U883 ( .A(n1191), .ZN(n1219) );
NAND4_X1 U884 ( .A1(n1221), .A2(n1061), .A3(n1203), .A4(n1222), .ZN(n1191) );
XNOR2_X1 U885 ( .A(G140), .B(n1179), .ZN(G42) );
NAND4_X1 U886 ( .A1(n1220), .A2(n1223), .A3(n1060), .A4(n1209), .ZN(n1179) );
XOR2_X1 U887 ( .A(G137), .B(n1224), .Z(G39) );
NOR3_X1 U888 ( .A1(n1192), .A2(n1225), .A3(n1065), .ZN(n1224) );
XOR2_X1 U889 ( .A(n1190), .B(KEYINPUT40), .Z(n1225) );
NAND4_X1 U890 ( .A1(n1223), .A2(n1092), .A3(n1075), .A4(n1226), .ZN(n1192) );
XNOR2_X1 U891 ( .A(G134), .B(n1178), .ZN(G36) );
NAND3_X1 U892 ( .A1(n1061), .A2(n1220), .A3(n1227), .ZN(n1178) );
NOR3_X1 U893 ( .A1(n1036), .A2(n1228), .A3(n1221), .ZN(n1227) );
XOR2_X1 U894 ( .A(n1229), .B(G131), .Z(G33) );
NAND2_X1 U895 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U896 ( .A1(n1183), .A2(n1232), .ZN(n1231) );
INV_X1 U897 ( .A(KEYINPUT34), .ZN(n1232) );
NOR2_X1 U898 ( .A1(n1233), .A2(n1036), .ZN(n1183) );
NAND3_X1 U899 ( .A1(n1223), .A2(n1233), .A3(KEYINPUT34), .ZN(n1230) );
NAND3_X1 U900 ( .A1(n1220), .A2(n1209), .A3(n1061), .ZN(n1233) );
INV_X1 U901 ( .A(n1036), .ZN(n1223) );
NAND2_X1 U902 ( .A1(n1096), .A2(n1234), .ZN(n1036) );
XNOR2_X1 U903 ( .A(G128), .B(n1180), .ZN(G30) );
NAND3_X1 U904 ( .A1(n1207), .A2(n1222), .A3(n1217), .ZN(n1180) );
AND4_X1 U905 ( .A1(n1220), .A2(n1203), .A3(n1075), .A4(n1226), .ZN(n1217) );
AND2_X1 U906 ( .A1(n1208), .A2(n1190), .ZN(n1220) );
XNOR2_X1 U907 ( .A(n1205), .B(n1235), .ZN(G3) );
NOR2_X1 U908 ( .A1(KEYINPUT27), .A2(n1236), .ZN(n1235) );
NAND3_X1 U909 ( .A1(n1092), .A2(n1208), .A3(n1237), .ZN(n1205) );
XNOR2_X1 U910 ( .A(G125), .B(n1177), .ZN(G27) );
NAND4_X1 U911 ( .A1(n1060), .A2(n1066), .A3(n1203), .A4(n1190), .ZN(n1177) );
NAND2_X1 U912 ( .A1(n1238), .A2(n1239), .ZN(n1190) );
NAND4_X1 U913 ( .A1(G953), .A2(G902), .A3(n1093), .A4(n1106), .ZN(n1239) );
INV_X1 U914 ( .A(G900), .ZN(n1106) );
NOR2_X1 U915 ( .A1(n1075), .A2(n1090), .ZN(n1060) );
INV_X1 U916 ( .A(n1226), .ZN(n1090) );
XNOR2_X1 U917 ( .A(G122), .B(n1195), .ZN(G24) );
NAND3_X1 U918 ( .A1(n1240), .A2(n1206), .A3(n1221), .ZN(n1195) );
AND3_X1 U919 ( .A1(n1210), .A2(n1222), .A3(n1054), .ZN(n1206) );
NOR2_X1 U920 ( .A1(n1226), .A2(n1075), .ZN(n1054) );
XNOR2_X1 U921 ( .A(n1198), .B(n1241), .ZN(G21) );
NAND2_X1 U922 ( .A1(KEYINPUT58), .A2(G119), .ZN(n1241) );
NOR3_X1 U923 ( .A1(n1074), .A2(n1242), .A3(n1211), .ZN(n1198) );
XOR2_X1 U924 ( .A(n1199), .B(n1243), .Z(G18) );
NOR2_X1 U925 ( .A1(KEYINPUT44), .A2(n1244), .ZN(n1243) );
AND2_X1 U926 ( .A1(n1049), .A2(n1237), .ZN(n1199) );
NOR3_X1 U927 ( .A1(n1221), .A2(n1228), .A3(n1074), .ZN(n1049) );
INV_X1 U928 ( .A(n1240), .ZN(n1074) );
INV_X1 U929 ( .A(n1222), .ZN(n1228) );
XOR2_X1 U930 ( .A(G113), .B(n1197), .Z(G15) );
AND2_X1 U931 ( .A1(n1237), .A2(n1066), .ZN(n1197) );
INV_X1 U932 ( .A(n1042), .ZN(n1066) );
NAND2_X1 U933 ( .A1(n1209), .A2(n1240), .ZN(n1042) );
NOR2_X1 U934 ( .A1(n1053), .A2(n1245), .ZN(n1240) );
INV_X1 U935 ( .A(n1052), .ZN(n1245) );
NOR2_X1 U936 ( .A1(n1207), .A2(n1222), .ZN(n1209) );
AND2_X1 U937 ( .A1(n1061), .A2(n1210), .ZN(n1237) );
NOR2_X1 U938 ( .A1(n1226), .A2(n1242), .ZN(n1061) );
INV_X1 U939 ( .A(n1075), .ZN(n1242) );
XNOR2_X1 U940 ( .A(n1246), .B(n1247), .ZN(G12) );
NOR3_X1 U941 ( .A1(n1211), .A2(n1248), .A3(n1075), .ZN(n1247) );
XNOR2_X1 U942 ( .A(n1249), .B(G472), .ZN(n1075) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1173), .ZN(n1249) );
XOR2_X1 U944 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U945 ( .A(n1152), .B(n1153), .Z(n1252) );
AND3_X1 U946 ( .A1(n1253), .A2(n1030), .A3(G210), .ZN(n1153) );
XOR2_X1 U947 ( .A(n1254), .B(n1255), .Z(n1152) );
XOR2_X1 U948 ( .A(G113), .B(n1256), .Z(n1255) );
NOR2_X1 U949 ( .A1(KEYINPUT51), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U950 ( .A(n1258), .B(G116), .ZN(n1257) );
XNOR2_X1 U951 ( .A(n1170), .B(n1110), .ZN(n1254) );
XNOR2_X1 U952 ( .A(n1259), .B(n1236), .ZN(n1251) );
XNOR2_X1 U953 ( .A(KEYINPUT33), .B(KEYINPUT2), .ZN(n1259) );
XNOR2_X1 U954 ( .A(n1208), .B(KEYINPUT1), .ZN(n1248) );
INV_X1 U955 ( .A(n1065), .ZN(n1208) );
NAND2_X1 U956 ( .A1(n1053), .A2(n1052), .ZN(n1065) );
NAND2_X1 U957 ( .A1(G221), .A2(n1260), .ZN(n1052) );
NAND2_X1 U958 ( .A1(G234), .A2(n1173), .ZN(n1260) );
XNOR2_X1 U959 ( .A(n1261), .B(G469), .ZN(n1053) );
NAND3_X1 U960 ( .A1(n1262), .A2(n1263), .A3(n1173), .ZN(n1261) );
NAND2_X1 U961 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
INV_X1 U962 ( .A(KEYINPUT32), .ZN(n1265) );
NAND2_X1 U963 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND3_X1 U964 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
INV_X1 U965 ( .A(KEYINPUT37), .ZN(n1269) );
NAND2_X1 U966 ( .A1(n1271), .A2(n1272), .ZN(n1266) );
NAND2_X1 U967 ( .A1(n1273), .A2(KEYINPUT32), .ZN(n1262) );
XNOR2_X1 U968 ( .A(n1271), .B(n1270), .ZN(n1273) );
INV_X1 U969 ( .A(n1272), .ZN(n1270) );
XNOR2_X1 U970 ( .A(n1274), .B(n1157), .ZN(n1272) );
AND2_X1 U971 ( .A1(G227), .A2(n1030), .ZN(n1157) );
NAND3_X1 U972 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1274) );
NAND2_X1 U973 ( .A1(KEYINPUT30), .A2(G110), .ZN(n1277) );
OR3_X1 U974 ( .A1(n1278), .A2(KEYINPUT30), .A3(G140), .ZN(n1276) );
NAND2_X1 U975 ( .A1(G140), .A2(n1278), .ZN(n1275) );
NAND2_X1 U976 ( .A1(KEYINPUT56), .A2(n1246), .ZN(n1278) );
AND2_X1 U977 ( .A1(KEYINPUT37), .A2(n1268), .ZN(n1271) );
XOR2_X1 U978 ( .A(n1279), .B(n1110), .Z(n1268) );
XOR2_X1 U979 ( .A(G131), .B(n1280), .Z(n1110) );
XOR2_X1 U980 ( .A(G137), .B(G134), .Z(n1280) );
NAND2_X1 U981 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NAND2_X1 U982 ( .A1(n1165), .A2(n1283), .ZN(n1282) );
XOR2_X1 U983 ( .A(KEYINPUT9), .B(n1284), .Z(n1281) );
NOR2_X1 U984 ( .A1(n1165), .A2(n1283), .ZN(n1284) );
XNOR2_X1 U985 ( .A(KEYINPUT45), .B(n1108), .ZN(n1283) );
XOR2_X1 U986 ( .A(n1285), .B(n1286), .Z(n1108) );
XNOR2_X1 U987 ( .A(G128), .B(KEYINPUT57), .ZN(n1285) );
XNOR2_X1 U988 ( .A(G101), .B(n1287), .ZN(n1165) );
NOR2_X1 U989 ( .A1(KEYINPUT25), .A2(n1288), .ZN(n1287) );
XNOR2_X1 U990 ( .A(n1289), .B(n1290), .ZN(n1288) );
NOR2_X1 U991 ( .A1(G104), .A2(KEYINPUT47), .ZN(n1290) );
INV_X1 U992 ( .A(G107), .ZN(n1289) );
NAND3_X1 U993 ( .A1(n1210), .A2(n1226), .A3(n1092), .ZN(n1211) );
NOR2_X1 U994 ( .A1(n1222), .A2(n1221), .ZN(n1092) );
INV_X1 U995 ( .A(n1207), .ZN(n1221) );
XNOR2_X1 U996 ( .A(n1086), .B(n1291), .ZN(n1207) );
NOR2_X1 U997 ( .A1(G475), .A2(KEYINPUT28), .ZN(n1291) );
NAND2_X1 U998 ( .A1(n1142), .A2(n1173), .ZN(n1086) );
XNOR2_X1 U999 ( .A(n1292), .B(n1293), .ZN(n1142) );
XOR2_X1 U1000 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1001 ( .A(G146), .B(n1112), .ZN(n1295) );
XOR2_X1 U1002 ( .A(KEYINPUT5), .B(KEYINPUT23), .Z(n1294) );
XOR2_X1 U1003 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U1004 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1005 ( .A1(KEYINPUT55), .A2(n1214), .ZN(n1298) );
XOR2_X1 U1006 ( .A(n1300), .B(G122), .Z(n1296) );
NAND2_X1 U1007 ( .A1(KEYINPUT61), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1008 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1009 ( .A(G143), .B(G131), .Z(n1303) );
NOR4_X1 U1010 ( .A1(KEYINPUT36), .A2(G953), .A3(G237), .A4(n1304), .ZN(n1302) );
INV_X1 U1011 ( .A(G214), .ZN(n1304) );
NAND3_X1 U1012 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1222) );
NAND2_X1 U1013 ( .A1(KEYINPUT22), .A2(n1089), .ZN(n1307) );
OR3_X1 U1014 ( .A1(n1089), .A2(KEYINPUT22), .A3(n1140), .ZN(n1306) );
NAND2_X1 U1015 ( .A1(n1308), .A2(n1140), .ZN(n1305) );
INV_X1 U1016 ( .A(G478), .ZN(n1140) );
NAND2_X1 U1017 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
INV_X1 U1018 ( .A(KEYINPUT22), .ZN(n1310) );
XNOR2_X1 U1019 ( .A(n1089), .B(KEYINPUT38), .ZN(n1309) );
NOR2_X1 U1020 ( .A1(n1137), .A2(G902), .ZN(n1089) );
XOR2_X1 U1021 ( .A(n1311), .B(n1312), .Z(n1137) );
NOR2_X1 U1022 ( .A1(KEYINPUT54), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1023 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1024 ( .A(n1316), .B(n1317), .ZN(n1315) );
XOR2_X1 U1025 ( .A(G143), .B(G134), .Z(n1317) );
XNOR2_X1 U1026 ( .A(G107), .B(n1318), .ZN(n1314) );
XNOR2_X1 U1027 ( .A(G122), .B(n1244), .ZN(n1318) );
NAND2_X1 U1028 ( .A1(n1319), .A2(G217), .ZN(n1311) );
NAND3_X1 U1029 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1226) );
NAND2_X1 U1030 ( .A1(G902), .A2(G217), .ZN(n1322) );
NAND3_X1 U1031 ( .A1(n1131), .A2(n1173), .A3(n1323), .ZN(n1321) );
OR2_X1 U1032 ( .A1(n1323), .A2(n1131), .ZN(n1320) );
XNOR2_X1 U1033 ( .A(n1324), .B(n1325), .ZN(n1131) );
XOR2_X1 U1034 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1035 ( .A(n1214), .B(G110), .ZN(n1327) );
XOR2_X1 U1036 ( .A(G146), .B(G137), .Z(n1326) );
XOR2_X1 U1037 ( .A(n1328), .B(n1329), .Z(n1324) );
XOR2_X1 U1038 ( .A(n1330), .B(n1331), .Z(n1329) );
NAND2_X1 U1039 ( .A1(KEYINPUT50), .A2(n1112), .ZN(n1331) );
INV_X1 U1040 ( .A(G140), .ZN(n1112) );
NAND3_X1 U1041 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1330) );
NAND2_X1 U1042 ( .A1(KEYINPUT26), .A2(n1258), .ZN(n1334) );
NAND3_X1 U1043 ( .A1(G119), .A2(n1335), .A3(n1316), .ZN(n1333) );
NAND2_X1 U1044 ( .A1(G128), .A2(n1336), .ZN(n1332) );
NAND2_X1 U1045 ( .A1(n1337), .A2(n1335), .ZN(n1336) );
INV_X1 U1046 ( .A(KEYINPUT26), .ZN(n1335) );
XNOR2_X1 U1047 ( .A(KEYINPUT53), .B(n1258), .ZN(n1337) );
NAND2_X1 U1048 ( .A1(n1319), .A2(G221), .ZN(n1328) );
NOR2_X1 U1049 ( .A1(n1338), .A2(G953), .ZN(n1319) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1338), .ZN(n1323) );
INV_X1 U1051 ( .A(G234), .ZN(n1338) );
NOR2_X1 U1052 ( .A1(n1094), .A2(n1201), .ZN(n1210) );
AND2_X1 U1053 ( .A1(n1238), .A2(n1339), .ZN(n1201) );
NAND4_X1 U1054 ( .A1(G953), .A2(G902), .A3(n1093), .A4(n1340), .ZN(n1339) );
INV_X1 U1055 ( .A(G898), .ZN(n1340) );
NAND3_X1 U1056 ( .A1(n1093), .A2(n1030), .A3(G952), .ZN(n1238) );
NAND2_X1 U1057 ( .A1(G237), .A2(G234), .ZN(n1093) );
INV_X1 U1058 ( .A(n1203), .ZN(n1094) );
NOR2_X1 U1059 ( .A1(n1096), .A2(n1072), .ZN(n1203) );
INV_X1 U1060 ( .A(n1234), .ZN(n1072) );
NAND2_X1 U1061 ( .A1(G214), .A2(n1341), .ZN(n1234) );
XNOR2_X1 U1062 ( .A(n1088), .B(n1342), .ZN(n1096) );
XOR2_X1 U1063 ( .A(KEYINPUT35), .B(n1343), .Z(n1342) );
NOR2_X1 U1064 ( .A1(KEYINPUT13), .A2(n1087), .ZN(n1343) );
AND2_X1 U1065 ( .A1(G210), .A2(n1341), .ZN(n1087) );
NAND2_X1 U1066 ( .A1(n1253), .A2(n1173), .ZN(n1341) );
INV_X1 U1067 ( .A(G237), .ZN(n1253) );
NAND2_X1 U1068 ( .A1(n1344), .A2(n1173), .ZN(n1088) );
INV_X1 U1069 ( .A(G902), .ZN(n1173) );
XOR2_X1 U1070 ( .A(n1345), .B(n1172), .Z(n1344) );
XNOR2_X1 U1071 ( .A(n1346), .B(KEYINPUT0), .ZN(n1172) );
INV_X1 U1072 ( .A(n1123), .ZN(n1346) );
XNOR2_X1 U1073 ( .A(n1347), .B(n1348), .ZN(n1123) );
XNOR2_X1 U1074 ( .A(n1236), .B(n1349), .ZN(n1348) );
XNOR2_X1 U1075 ( .A(n1246), .B(G107), .ZN(n1349) );
INV_X1 U1076 ( .A(G101), .ZN(n1236) );
XNOR2_X1 U1077 ( .A(n1299), .B(n1350), .ZN(n1347) );
XOR2_X1 U1078 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND2_X1 U1079 ( .A1(KEYINPUT48), .A2(G122), .ZN(n1352) );
NAND3_X1 U1080 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1351) );
NAND2_X1 U1081 ( .A1(G119), .A2(n1244), .ZN(n1355) );
INV_X1 U1082 ( .A(G116), .ZN(n1244) );
NAND2_X1 U1083 ( .A1(KEYINPUT41), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1084 ( .A1(n1357), .A2(n1258), .ZN(n1356) );
XNOR2_X1 U1085 ( .A(KEYINPUT42), .B(G116), .ZN(n1357) );
NAND2_X1 U1086 ( .A1(n1358), .A2(n1359), .ZN(n1353) );
INV_X1 U1087 ( .A(KEYINPUT41), .ZN(n1359) );
NAND2_X1 U1088 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
OR2_X1 U1089 ( .A1(G116), .A2(KEYINPUT42), .ZN(n1361) );
NAND3_X1 U1090 ( .A1(G116), .A2(n1258), .A3(KEYINPUT42), .ZN(n1360) );
INV_X1 U1091 ( .A(G119), .ZN(n1258) );
XOR2_X1 U1092 ( .A(G104), .B(G113), .Z(n1299) );
NAND2_X1 U1093 ( .A1(KEYINPUT46), .A2(n1362), .ZN(n1345) );
XNOR2_X1 U1094 ( .A(n1170), .B(n1363), .ZN(n1362) );
XNOR2_X1 U1095 ( .A(n1364), .B(n1214), .ZN(n1363) );
INV_X1 U1096 ( .A(G125), .ZN(n1214) );
NAND2_X1 U1097 ( .A1(KEYINPUT11), .A2(n1215), .ZN(n1364) );
AND2_X1 U1098 ( .A1(n1365), .A2(n1030), .ZN(n1215) );
INV_X1 U1099 ( .A(G953), .ZN(n1030) );
XNOR2_X1 U1100 ( .A(G224), .B(KEYINPUT14), .ZN(n1365) );
XNOR2_X1 U1101 ( .A(n1366), .B(n1286), .ZN(n1170) );
XOR2_X1 U1102 ( .A(G143), .B(G146), .Z(n1286) );
NAND2_X1 U1103 ( .A1(KEYINPUT24), .A2(n1316), .ZN(n1366) );
INV_X1 U1104 ( .A(G128), .ZN(n1316) );
INV_X1 U1105 ( .A(G110), .ZN(n1246) );
endmodule


