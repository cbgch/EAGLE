//Key = 1000001000000001000100011001011110100110011001100111110111001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346;

XNOR2_X1 U750 ( .A(G107), .B(n1020), .ZN(G9) );
NAND3_X1 U751 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
XOR2_X1 U752 ( .A(KEYINPUT11), .B(n1024), .Z(n1022) );
NOR2_X1 U753 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
INV_X1 U755 ( .A(G952), .ZN(n1029) );
XOR2_X1 U756 ( .A(KEYINPUT20), .B(n1031), .Z(n1028) );
NOR2_X1 U757 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U758 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U759 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U760 ( .A1(n1038), .A2(n1039), .ZN(n1034) );
INV_X1 U761 ( .A(n1040), .ZN(n1039) );
NOR2_X1 U762 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
NOR2_X1 U763 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U764 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
AND2_X1 U765 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U766 ( .A1(n1037), .A2(n1049), .ZN(n1041) );
XOR2_X1 U767 ( .A(KEYINPUT19), .B(n1024), .Z(n1049) );
NAND3_X1 U768 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1027) );
NAND2_X1 U769 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U770 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U771 ( .A1(n1057), .A2(n1023), .A3(n1058), .ZN(n1056) );
NAND2_X1 U772 ( .A1(n1040), .A2(n1059), .ZN(n1055) );
NAND2_X1 U773 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U774 ( .A1(n1062), .A2(n1058), .A3(n1063), .ZN(n1061) );
INV_X1 U775 ( .A(n1037), .ZN(n1058) );
NAND2_X1 U776 ( .A1(n1064), .A2(n1048), .ZN(n1037) );
NAND2_X1 U777 ( .A1(n1057), .A2(n1065), .ZN(n1060) );
NAND2_X1 U778 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U779 ( .A1(n1068), .A2(n1048), .A3(n1069), .ZN(n1067) );
NAND2_X1 U780 ( .A1(n1070), .A2(n1064), .ZN(n1066) );
INV_X1 U781 ( .A(n1033), .ZN(n1053) );
NOR3_X1 U782 ( .A1(n1071), .A2(G953), .A3(n1072), .ZN(n1025) );
INV_X1 U783 ( .A(n1050), .ZN(n1072) );
NAND4_X1 U784 ( .A1(n1073), .A2(n1040), .A3(n1074), .A4(n1075), .ZN(n1050) );
NOR4_X1 U785 ( .A1(n1069), .A2(n1063), .A3(n1076), .A4(n1077), .ZN(n1075) );
XOR2_X1 U786 ( .A(n1068), .B(KEYINPUT29), .Z(n1077) );
NOR2_X1 U787 ( .A1(G469), .A2(n1078), .ZN(n1076) );
NOR3_X1 U788 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1074) );
NOR2_X1 U789 ( .A1(KEYINPUT21), .A2(n1082), .ZN(n1081) );
NOR2_X1 U790 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
AND3_X1 U791 ( .A1(KEYINPUT51), .A2(n1078), .A3(G469), .ZN(n1084) );
NOR2_X1 U792 ( .A1(KEYINPUT51), .A2(G469), .ZN(n1083) );
NOR2_X1 U793 ( .A1(n1085), .A2(n1086), .ZN(n1080) );
INV_X1 U794 ( .A(KEYINPUT21), .ZN(n1086) );
NOR2_X1 U795 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XNOR2_X1 U796 ( .A(KEYINPUT51), .B(n1089), .ZN(n1088) );
INV_X1 U797 ( .A(n1078), .ZN(n1087) );
XOR2_X1 U798 ( .A(n1090), .B(n1091), .Z(n1079) );
XOR2_X1 U799 ( .A(n1092), .B(G472), .Z(n1091) );
XNOR2_X1 U800 ( .A(KEYINPUT53), .B(KEYINPUT27), .ZN(n1090) );
XNOR2_X1 U801 ( .A(G952), .B(KEYINPUT41), .ZN(n1071) );
XOR2_X1 U802 ( .A(n1093), .B(n1094), .Z(G72) );
XOR2_X1 U803 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U804 ( .A1(n1097), .A2(n1051), .ZN(n1096) );
AND2_X1 U805 ( .A1(G227), .A2(G900), .ZN(n1097) );
NAND2_X1 U806 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NAND2_X1 U807 ( .A1(G953), .A2(n1100), .ZN(n1099) );
XOR2_X1 U808 ( .A(n1101), .B(n1102), .Z(n1098) );
XOR2_X1 U809 ( .A(n1103), .B(n1104), .Z(n1102) );
XNOR2_X1 U810 ( .A(n1105), .B(n1106), .ZN(n1103) );
NAND2_X1 U811 ( .A1(KEYINPUT32), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U812 ( .A(G128), .B(n1108), .ZN(n1101) );
XOR2_X1 U813 ( .A(KEYINPUT36), .B(G143), .Z(n1108) );
NAND2_X1 U814 ( .A1(n1051), .A2(n1109), .ZN(n1093) );
NAND2_X1 U815 ( .A1(n1110), .A2(n1111), .ZN(G69) );
NAND2_X1 U816 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
OR2_X1 U817 ( .A1(n1051), .A2(G224), .ZN(n1113) );
NAND3_X1 U818 ( .A1(n1114), .A2(n1115), .A3(G953), .ZN(n1110) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1115) );
XOR2_X1 U820 ( .A(KEYINPUT30), .B(n1112), .Z(n1114) );
XNOR2_X1 U821 ( .A(n1116), .B(n1117), .ZN(n1112) );
NOR2_X1 U822 ( .A1(G953), .A2(n1118), .ZN(n1117) );
NOR2_X1 U823 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U824 ( .A(KEYINPUT24), .B(n1121), .Z(n1120) );
NOR2_X1 U825 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND3_X1 U826 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1116) );
XOR2_X1 U827 ( .A(KEYINPUT34), .B(n1127), .Z(n1126) );
NOR2_X1 U828 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U829 ( .A(n1130), .B(KEYINPUT37), .ZN(n1128) );
NAND2_X1 U830 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
XOR2_X1 U831 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U832 ( .A1(KEYINPUT59), .A2(n1133), .ZN(n1132) );
XOR2_X1 U833 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U834 ( .A(KEYINPUT60), .B(n1136), .ZN(n1135) );
XNOR2_X1 U835 ( .A(G101), .B(G104), .ZN(n1134) );
XNOR2_X1 U836 ( .A(G122), .B(n1137), .ZN(n1129) );
NAND2_X1 U837 ( .A1(G953), .A2(n1138), .ZN(n1124) );
NOR3_X1 U838 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(G66) );
NOR3_X1 U839 ( .A1(n1142), .A2(G953), .A3(G952), .ZN(n1141) );
AND2_X1 U840 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
INV_X1 U841 ( .A(KEYINPUT7), .ZN(n1142) );
XOR2_X1 U842 ( .A(n1144), .B(n1145), .Z(n1139) );
NOR2_X1 U843 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U844 ( .A1(KEYINPUT50), .A2(n1148), .ZN(n1144) );
NOR2_X1 U845 ( .A1(n1143), .A2(n1149), .ZN(G63) );
XOR2_X1 U846 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND3_X1 U847 ( .A1(n1152), .A2(G478), .A3(KEYINPUT49), .ZN(n1150) );
NOR2_X1 U848 ( .A1(n1153), .A2(n1154), .ZN(G60) );
XOR2_X1 U849 ( .A(KEYINPUT8), .B(n1143), .Z(n1154) );
XNOR2_X1 U850 ( .A(n1155), .B(n1156), .ZN(n1153) );
XOR2_X1 U851 ( .A(KEYINPUT43), .B(n1157), .Z(n1156) );
AND2_X1 U852 ( .A1(G475), .A2(n1152), .ZN(n1157) );
XNOR2_X1 U853 ( .A(G104), .B(n1158), .ZN(G6) );
NOR2_X1 U854 ( .A1(n1143), .A2(n1159), .ZN(G57) );
XOR2_X1 U855 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U856 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U857 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NAND2_X1 U858 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U859 ( .A(KEYINPUT26), .ZN(n1167) );
XNOR2_X1 U860 ( .A(n1168), .B(n1106), .ZN(n1166) );
NAND3_X1 U861 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT26), .ZN(n1164) );
XOR2_X1 U862 ( .A(n1170), .B(n1171), .Z(n1160) );
AND2_X1 U863 ( .A1(G472), .A2(n1152), .ZN(n1171) );
NOR2_X1 U864 ( .A1(n1143), .A2(n1172), .ZN(G54) );
XOR2_X1 U865 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U866 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U867 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U868 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
XNOR2_X1 U869 ( .A(KEYINPUT25), .B(n1181), .ZN(n1180) );
NOR2_X1 U870 ( .A1(n1089), .A2(n1147), .ZN(n1175) );
INV_X1 U871 ( .A(G469), .ZN(n1089) );
XOR2_X1 U872 ( .A(KEYINPUT48), .B(n1182), .Z(n1173) );
NOR2_X1 U873 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U874 ( .A(n1185), .B(KEYINPUT15), .ZN(n1184) );
NOR2_X1 U875 ( .A1(n1143), .A2(n1186), .ZN(G51) );
XOR2_X1 U876 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U877 ( .A(n1189), .B(n1190), .Z(n1188) );
NAND3_X1 U878 ( .A1(n1152), .A2(G210), .A3(KEYINPUT6), .ZN(n1189) );
INV_X1 U879 ( .A(n1147), .ZN(n1152) );
NAND2_X1 U880 ( .A1(G902), .A2(n1030), .ZN(n1147) );
OR4_X1 U881 ( .A1(n1109), .A2(n1119), .A3(n1123), .A4(n1191), .ZN(n1030) );
XNOR2_X1 U882 ( .A(KEYINPUT31), .B(n1122), .ZN(n1191) );
INV_X1 U883 ( .A(n1192), .ZN(n1122) );
NAND3_X1 U884 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1123) );
NAND4_X1 U885 ( .A1(n1196), .A2(n1158), .A3(n1197), .A4(n1198), .ZN(n1119) );
NAND3_X1 U886 ( .A1(n1021), .A2(n1024), .A3(n1199), .ZN(n1158) );
INV_X1 U887 ( .A(n1200), .ZN(n1199) );
NAND3_X1 U888 ( .A1(n1021), .A2(n1024), .A3(n1023), .ZN(n1196) );
NAND4_X1 U889 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1109) );
AND4_X1 U890 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NAND2_X1 U891 ( .A1(n1070), .A2(n1209), .ZN(n1203) );
NAND2_X1 U892 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U893 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U894 ( .A(KEYINPUT35), .B(n1214), .ZN(n1213) );
NAND2_X1 U895 ( .A1(n1215), .A2(n1216), .ZN(n1210) );
NAND3_X1 U896 ( .A1(n1046), .A2(n1217), .A3(n1218), .ZN(n1201) );
XNOR2_X1 U897 ( .A(n1023), .B(KEYINPUT42), .ZN(n1218) );
XOR2_X1 U898 ( .A(n1219), .B(KEYINPUT40), .Z(n1187) );
NAND2_X1 U899 ( .A1(KEYINPUT46), .A2(n1220), .ZN(n1219) );
NOR2_X1 U900 ( .A1(n1051), .A2(G952), .ZN(n1143) );
XNOR2_X1 U901 ( .A(G146), .B(n1202), .ZN(G48) );
NAND3_X1 U902 ( .A1(n1221), .A2(n1047), .A3(n1212), .ZN(n1202) );
XNOR2_X1 U903 ( .A(G143), .B(n1208), .ZN(G45) );
NAND4_X1 U904 ( .A1(n1222), .A2(n1223), .A3(n1047), .A4(n1224), .ZN(n1208) );
NOR2_X1 U905 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U906 ( .A(G140), .B(n1227), .ZN(G42) );
NAND3_X1 U907 ( .A1(n1070), .A2(n1212), .A3(n1228), .ZN(n1227) );
XNOR2_X1 U908 ( .A(n1064), .B(KEYINPUT23), .ZN(n1228) );
XOR2_X1 U909 ( .A(n1207), .B(n1229), .Z(G39) );
NOR2_X1 U910 ( .A1(G137), .A2(KEYINPUT62), .ZN(n1229) );
NAND4_X1 U911 ( .A1(n1064), .A2(n1217), .A3(n1221), .A4(n1040), .ZN(n1207) );
INV_X1 U912 ( .A(n1214), .ZN(n1064) );
XNOR2_X1 U913 ( .A(n1230), .B(n1231), .ZN(G36) );
AND3_X1 U914 ( .A1(n1046), .A2(n1023), .A3(n1217), .ZN(n1231) );
INV_X1 U915 ( .A(n1225), .ZN(n1217) );
XNOR2_X1 U916 ( .A(G131), .B(n1206), .ZN(G33) );
NAND2_X1 U917 ( .A1(n1212), .A2(n1046), .ZN(n1206) );
NOR2_X1 U918 ( .A1(n1214), .A2(n1226), .ZN(n1046) );
NAND2_X1 U919 ( .A1(n1068), .A2(n1232), .ZN(n1214) );
NOR2_X1 U920 ( .A1(n1200), .A2(n1225), .ZN(n1212) );
NAND2_X1 U921 ( .A1(n1233), .A2(n1234), .ZN(n1225) );
XNOR2_X1 U922 ( .A(n1024), .B(KEYINPUT19), .ZN(n1233) );
XNOR2_X1 U923 ( .A(G128), .B(n1205), .ZN(G30) );
NAND4_X1 U924 ( .A1(n1221), .A2(n1216), .A3(n1023), .A4(n1024), .ZN(n1205) );
XNOR2_X1 U925 ( .A(G101), .B(n1197), .ZN(G3) );
NAND2_X1 U926 ( .A1(n1235), .A2(n1236), .ZN(n1197) );
XNOR2_X1 U927 ( .A(G125), .B(n1237), .ZN(G27) );
NAND4_X1 U928 ( .A1(n1070), .A2(n1216), .A3(n1238), .A4(n1239), .ZN(n1237) );
NAND2_X1 U929 ( .A1(KEYINPUT0), .A2(n1036), .ZN(n1239) );
INV_X1 U930 ( .A(n1215), .ZN(n1036) );
NAND2_X1 U931 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
INV_X1 U932 ( .A(KEYINPUT0), .ZN(n1241) );
NAND2_X1 U933 ( .A1(n1057), .A2(n1200), .ZN(n1240) );
AND2_X1 U934 ( .A1(n1047), .A2(n1234), .ZN(n1216) );
NAND2_X1 U935 ( .A1(n1033), .A2(n1242), .ZN(n1234) );
NAND4_X1 U936 ( .A1(G953), .A2(G902), .A3(n1100), .A4(n1243), .ZN(n1242) );
XOR2_X1 U937 ( .A(KEYINPUT56), .B(G900), .Z(n1100) );
NAND2_X1 U938 ( .A1(n1244), .A2(n1245), .ZN(G24) );
NAND2_X1 U939 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U940 ( .A(KEYINPUT57), .B(n1248), .Z(n1244) );
NOR2_X1 U941 ( .A1(n1246), .A2(n1247), .ZN(n1248) );
INV_X1 U942 ( .A(n1195), .ZN(n1246) );
NAND4_X1 U943 ( .A1(n1057), .A2(n1021), .A3(n1222), .A4(n1223), .ZN(n1195) );
AND2_X1 U944 ( .A1(n1249), .A2(n1048), .ZN(n1021) );
AND2_X1 U945 ( .A1(n1073), .A2(n1250), .ZN(n1048) );
XNOR2_X1 U946 ( .A(G119), .B(n1193), .ZN(G21) );
NAND4_X1 U947 ( .A1(n1057), .A2(n1221), .A3(n1040), .A4(n1249), .ZN(n1193) );
AND2_X1 U948 ( .A1(n1251), .A2(n1252), .ZN(n1221) );
NAND2_X1 U949 ( .A1(n1253), .A2(n1254), .ZN(G18) );
NAND2_X1 U950 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U951 ( .A(KEYINPUT4), .B(n1194), .ZN(n1255) );
NAND2_X1 U952 ( .A1(G116), .A2(n1257), .ZN(n1253) );
XOR2_X1 U953 ( .A(n1194), .B(KEYINPUT33), .Z(n1257) );
NAND4_X1 U954 ( .A1(n1057), .A2(n1236), .A3(n1023), .A4(n1249), .ZN(n1194) );
NOR2_X1 U955 ( .A1(n1222), .A2(n1258), .ZN(n1023) );
INV_X1 U956 ( .A(n1044), .ZN(n1057) );
XNOR2_X1 U957 ( .A(G113), .B(n1192), .ZN(G15) );
NAND3_X1 U958 ( .A1(n1236), .A2(n1249), .A3(n1215), .ZN(n1192) );
NOR2_X1 U959 ( .A1(n1044), .A2(n1200), .ZN(n1215) );
NAND2_X1 U960 ( .A1(n1258), .A2(n1222), .ZN(n1200) );
INV_X1 U961 ( .A(n1223), .ZN(n1258) );
NAND2_X1 U962 ( .A1(n1259), .A2(n1260), .ZN(n1044) );
XOR2_X1 U963 ( .A(KEYINPUT17), .B(n1062), .Z(n1259) );
INV_X1 U964 ( .A(n1226), .ZN(n1236) );
NAND2_X1 U965 ( .A1(n1073), .A2(n1251), .ZN(n1226) );
XNOR2_X1 U966 ( .A(n1250), .B(KEYINPUT47), .ZN(n1251) );
INV_X1 U967 ( .A(n1252), .ZN(n1073) );
XNOR2_X1 U968 ( .A(n1198), .B(n1261), .ZN(G12) );
XNOR2_X1 U969 ( .A(KEYINPUT13), .B(n1262), .ZN(n1261) );
NAND2_X1 U970 ( .A1(n1235), .A2(n1070), .ZN(n1198) );
AND2_X1 U971 ( .A1(n1250), .A2(n1252), .ZN(n1070) );
XOR2_X1 U972 ( .A(n1263), .B(n1146), .Z(n1252) );
NAND2_X1 U973 ( .A1(G217), .A2(n1264), .ZN(n1146) );
NAND2_X1 U974 ( .A1(n1148), .A2(n1265), .ZN(n1263) );
XOR2_X1 U975 ( .A(n1266), .B(n1267), .Z(n1148) );
XOR2_X1 U976 ( .A(G137), .B(n1268), .Z(n1267) );
NOR2_X1 U977 ( .A1(KEYINPUT28), .A2(n1269), .ZN(n1268) );
XOR2_X1 U978 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U979 ( .A(n1272), .B(n1262), .ZN(n1271) );
INV_X1 U980 ( .A(G110), .ZN(n1262) );
NAND2_X1 U981 ( .A1(KEYINPUT52), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U982 ( .A(G119), .B(G128), .ZN(n1270) );
NAND2_X1 U983 ( .A1(G221), .A2(n1274), .ZN(n1266) );
XNOR2_X1 U984 ( .A(n1275), .B(n1092), .ZN(n1250) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1276), .ZN(n1092) );
XOR2_X1 U986 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U987 ( .A(n1279), .B(n1106), .ZN(n1278) );
NOR2_X1 U988 ( .A1(KEYINPUT39), .A2(n1170), .ZN(n1279) );
NAND2_X1 U989 ( .A1(G210), .A2(n1280), .ZN(n1170) );
NAND2_X1 U990 ( .A1(KEYINPUT38), .A2(G472), .ZN(n1275) );
AND3_X1 U991 ( .A1(n1024), .A2(n1249), .A3(n1040), .ZN(n1235) );
NOR2_X1 U992 ( .A1(n1223), .A2(n1222), .ZN(n1040) );
XNOR2_X1 U993 ( .A(n1281), .B(G475), .ZN(n1222) );
NAND2_X1 U994 ( .A1(n1265), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U995 ( .A(KEYINPUT12), .B(n1283), .ZN(n1282) );
INV_X1 U996 ( .A(n1155), .ZN(n1283) );
XNOR2_X1 U997 ( .A(n1284), .B(n1285), .ZN(n1155) );
XOR2_X1 U998 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U999 ( .A(G143), .B(n1288), .ZN(n1287) );
NOR2_X1 U1000 ( .A1(KEYINPUT16), .A2(G131), .ZN(n1286) );
XNOR2_X1 U1001 ( .A(n1273), .B(n1289), .ZN(n1284) );
XOR2_X1 U1002 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U1003 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U1004 ( .A1(G122), .A2(n1294), .ZN(n1293) );
INV_X1 U1005 ( .A(G113), .ZN(n1294) );
XOR2_X1 U1006 ( .A(n1295), .B(KEYINPUT5), .Z(n1292) );
NAND2_X1 U1007 ( .A1(G113), .A2(n1247), .ZN(n1295) );
INV_X1 U1008 ( .A(G122), .ZN(n1247) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1280), .ZN(n1290) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1280) );
XOR2_X1 U1011 ( .A(G140), .B(n1104), .Z(n1273) );
XOR2_X1 U1012 ( .A(G125), .B(G146), .Z(n1104) );
XNOR2_X1 U1013 ( .A(n1296), .B(G478), .ZN(n1223) );
NAND2_X1 U1014 ( .A1(n1265), .A2(n1151), .ZN(n1296) );
XOR2_X1 U1015 ( .A(n1297), .B(n1298), .Z(n1151) );
XOR2_X1 U1016 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1017 ( .A(G134), .B(G128), .ZN(n1300) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1274), .ZN(n1299) );
AND2_X1 U1019 ( .A1(G234), .A2(n1051), .ZN(n1274) );
XOR2_X1 U1020 ( .A(n1301), .B(n1302), .Z(n1297) );
XOR2_X1 U1021 ( .A(n1303), .B(n1304), .Z(n1302) );
NOR2_X1 U1022 ( .A1(G143), .A2(KEYINPUT54), .ZN(n1303) );
AND2_X1 U1023 ( .A1(n1047), .A2(n1305), .ZN(n1249) );
NAND2_X1 U1024 ( .A1(n1033), .A2(n1306), .ZN(n1305) );
NAND4_X1 U1025 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1138), .ZN(n1306) );
INV_X1 U1026 ( .A(G898), .ZN(n1138) );
NAND3_X1 U1027 ( .A1(n1243), .A2(n1051), .A3(G952), .ZN(n1033) );
NAND2_X1 U1028 ( .A1(G237), .A2(G234), .ZN(n1243) );
NOR2_X1 U1029 ( .A1(n1068), .A2(n1069), .ZN(n1047) );
INV_X1 U1030 ( .A(n1232), .ZN(n1069) );
NAND2_X1 U1031 ( .A1(n1307), .A2(n1308), .ZN(n1232) );
XOR2_X1 U1032 ( .A(KEYINPUT10), .B(G214), .Z(n1307) );
XOR2_X1 U1033 ( .A(n1309), .B(n1310), .Z(n1068) );
AND2_X1 U1034 ( .A1(n1308), .A2(G210), .ZN(n1310) );
OR2_X1 U1035 ( .A1(G902), .A2(G237), .ZN(n1308) );
NAND2_X1 U1036 ( .A1(n1265), .A2(n1311), .ZN(n1309) );
XNOR2_X1 U1037 ( .A(n1190), .B(n1220), .ZN(n1311) );
NAND2_X1 U1038 ( .A1(n1312), .A2(n1051), .ZN(n1220) );
XOR2_X1 U1039 ( .A(KEYINPUT44), .B(G224), .Z(n1312) );
XOR2_X1 U1040 ( .A(n1313), .B(n1314), .Z(n1190) );
XOR2_X1 U1041 ( .A(n1137), .B(n1301), .Z(n1314) );
XNOR2_X1 U1042 ( .A(G107), .B(G122), .ZN(n1301) );
XNOR2_X1 U1043 ( .A(KEYINPUT55), .B(n1315), .ZN(n1137) );
NOR2_X1 U1044 ( .A1(G110), .A2(KEYINPUT1), .ZN(n1315) );
XOR2_X1 U1045 ( .A(n1277), .B(n1316), .Z(n1313) );
XNOR2_X1 U1046 ( .A(G125), .B(n1288), .ZN(n1316) );
XOR2_X1 U1047 ( .A(n1163), .B(n1168), .Z(n1277) );
NAND2_X1 U1048 ( .A1(n1317), .A2(n1318), .ZN(n1168) );
OR2_X1 U1049 ( .A1(n1319), .A2(KEYINPUT9), .ZN(n1318) );
NAND3_X1 U1050 ( .A1(G128), .A2(n1320), .A3(KEYINPUT9), .ZN(n1317) );
XNOR2_X1 U1051 ( .A(G101), .B(n1321), .ZN(n1163) );
INV_X1 U1052 ( .A(n1131), .ZN(n1321) );
XNOR2_X1 U1053 ( .A(n1322), .B(n1304), .ZN(n1131) );
XNOR2_X1 U1054 ( .A(n1256), .B(KEYINPUT18), .ZN(n1304) );
INV_X1 U1055 ( .A(G116), .ZN(n1256) );
XNOR2_X1 U1056 ( .A(G119), .B(G113), .ZN(n1322) );
NOR2_X1 U1057 ( .A1(n1062), .A2(n1063), .ZN(n1024) );
INV_X1 U1058 ( .A(n1260), .ZN(n1063) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1264), .ZN(n1260) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1323), .ZN(n1264) );
INV_X1 U1061 ( .A(G902), .ZN(n1323) );
XOR2_X1 U1062 ( .A(G469), .B(n1324), .Z(n1062) );
NOR2_X1 U1063 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
AND2_X1 U1064 ( .A1(KEYINPUT3), .A2(n1078), .ZN(n1326) );
NOR2_X1 U1065 ( .A1(KEYINPUT58), .A2(n1078), .ZN(n1325) );
NAND4_X1 U1066 ( .A1(n1265), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1078) );
OR3_X1 U1067 ( .A1(n1179), .A2(n1330), .A3(n1181), .ZN(n1329) );
INV_X1 U1068 ( .A(n1331), .ZN(n1179) );
NAND2_X1 U1069 ( .A1(n1332), .A2(n1181), .ZN(n1328) );
XNOR2_X1 U1070 ( .A(n1331), .B(n1330), .ZN(n1332) );
NAND2_X1 U1071 ( .A1(n1178), .A2(n1330), .ZN(n1327) );
NOR3_X1 U1072 ( .A1(KEYINPUT22), .A2(n1183), .A3(n1185), .ZN(n1330) );
AND2_X1 U1073 ( .A1(n1333), .A2(n1169), .ZN(n1185) );
XNOR2_X1 U1074 ( .A(n1334), .B(n1335), .ZN(n1333) );
AND2_X1 U1075 ( .A1(n1336), .A2(n1106), .ZN(n1183) );
INV_X1 U1076 ( .A(n1169), .ZN(n1106) );
XOR2_X1 U1077 ( .A(G131), .B(n1337), .Z(n1169) );
XNOR2_X1 U1078 ( .A(G137), .B(n1230), .ZN(n1337) );
INV_X1 U1079 ( .A(G134), .ZN(n1230) );
XNOR2_X1 U1080 ( .A(n1335), .B(n1319), .ZN(n1336) );
INV_X1 U1081 ( .A(n1334), .ZN(n1319) );
XOR2_X1 U1082 ( .A(G128), .B(n1320), .Z(n1334) );
XOR2_X1 U1083 ( .A(G146), .B(G143), .Z(n1320) );
XOR2_X1 U1084 ( .A(n1338), .B(n1339), .Z(n1335) );
NOR2_X1 U1085 ( .A1(G101), .A2(KEYINPUT63), .ZN(n1339) );
NAND3_X1 U1086 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1338) );
NAND2_X1 U1087 ( .A1(KEYINPUT14), .A2(G104), .ZN(n1342) );
NAND3_X1 U1088 ( .A1(n1288), .A2(n1343), .A3(G107), .ZN(n1341) );
INV_X1 U1089 ( .A(G104), .ZN(n1288) );
NAND2_X1 U1090 ( .A1(n1344), .A2(n1136), .ZN(n1340) );
INV_X1 U1091 ( .A(G107), .ZN(n1136) );
NAND2_X1 U1092 ( .A1(n1345), .A2(n1343), .ZN(n1344) );
INV_X1 U1093 ( .A(KEYINPUT14), .ZN(n1343) );
XNOR2_X1 U1094 ( .A(G104), .B(KEYINPUT61), .ZN(n1345) );
NOR2_X1 U1095 ( .A1(n1181), .A2(n1331), .ZN(n1178) );
XNOR2_X1 U1096 ( .A(G110), .B(n1107), .ZN(n1331) );
INV_X1 U1097 ( .A(G140), .ZN(n1107) );
NAND2_X1 U1098 ( .A1(G227), .A2(n1346), .ZN(n1181) );
XNOR2_X1 U1099 ( .A(KEYINPUT45), .B(n1051), .ZN(n1346) );
INV_X1 U1100 ( .A(G953), .ZN(n1051) );
XNOR2_X1 U1101 ( .A(G902), .B(KEYINPUT2), .ZN(n1265) );
endmodule


