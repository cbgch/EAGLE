//Key = 0111011011011110000011010011011110111101000000111100101101101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294;

XOR2_X1 U715 ( .A(G107), .B(n988), .Z(G9) );
NOR2_X1 U716 ( .A1(n989), .A2(n990), .ZN(G75) );
NOR3_X1 U717 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NAND3_X1 U718 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n991) );
NAND2_X1 U719 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U720 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND3_X1 U721 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NAND3_X1 U722 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1002) );
NAND2_X1 U723 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1005) );
NAND2_X1 U725 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U726 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U727 ( .A1(n1015), .A2(n1016), .ZN(n1004) );
XOR2_X1 U728 ( .A(KEYINPUT42), .B(n1007), .Z(n1015) );
NAND3_X1 U729 ( .A1(n1009), .A2(n1017), .A3(n1007), .ZN(n999) );
NAND2_X1 U730 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U731 ( .A1(n1003), .A2(n1020), .ZN(n1019) );
OR2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U733 ( .A1(n1001), .A2(n1023), .ZN(n1018) );
NAND2_X1 U734 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XOR2_X1 U736 ( .A(KEYINPUT63), .B(n1028), .Z(n1027) );
INV_X1 U737 ( .A(n1029), .ZN(n997) );
NOR3_X1 U738 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n989) );
INV_X1 U739 ( .A(n994), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n994) );
NOR4_X1 U741 ( .A1(n1013), .A2(n1026), .A3(n1033), .A4(n1034), .ZN(n1032) );
NOR4_X1 U742 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1031) );
XNOR2_X1 U743 ( .A(G475), .B(n1039), .ZN(n1038) );
XNOR2_X1 U744 ( .A(n1040), .B(n1041), .ZN(n1037) );
XOR2_X1 U745 ( .A(n1042), .B(n1043), .Z(n1036) );
NAND2_X1 U746 ( .A1(KEYINPUT52), .A2(G472), .ZN(n1043) );
XOR2_X1 U747 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U748 ( .A1(n1046), .A2(n995), .ZN(n1045) );
AND2_X1 U749 ( .A1(G227), .A2(G900), .ZN(n1046) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NAND2_X1 U751 ( .A1(n1049), .A2(n995), .ZN(n1048) );
XOR2_X1 U752 ( .A(n992), .B(n1050), .Z(n1049) );
NAND3_X1 U753 ( .A1(n1050), .A2(n1051), .A3(G953), .ZN(n1047) );
INV_X1 U754 ( .A(n1052), .ZN(n1051) );
XNOR2_X1 U755 ( .A(n1053), .B(n1054), .ZN(n1050) );
XOR2_X1 U756 ( .A(n1055), .B(n1056), .Z(n1053) );
XOR2_X1 U757 ( .A(n1057), .B(n1058), .Z(G69) );
XOR2_X1 U758 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U759 ( .A1(n1061), .A2(n995), .ZN(n1060) );
AND2_X1 U760 ( .A1(G224), .A2(G898), .ZN(n1061) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NAND2_X1 U762 ( .A1(G953), .A2(n1064), .ZN(n1063) );
XOR2_X1 U763 ( .A(n1065), .B(n1066), .Z(n1062) );
NOR2_X1 U764 ( .A1(KEYINPUT40), .A2(n1067), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n995), .A2(n1068), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U767 ( .A(KEYINPUT26), .B(n1071), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XNOR2_X1 U769 ( .A(n1074), .B(KEYINPUT37), .ZN(n1073) );
XOR2_X1 U770 ( .A(n1075), .B(n1076), .Z(n1072) );
NOR2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U772 ( .A1(KEYINPUT29), .A2(n1079), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U775 ( .A1(KEYINPUT56), .A2(n1083), .ZN(n1082) );
AND2_X1 U776 ( .A1(G478), .A2(n1084), .ZN(n1081) );
NOR2_X1 U777 ( .A1(n1074), .A2(n1085), .ZN(G60) );
XOR2_X1 U778 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U779 ( .A1(n1084), .A2(G475), .ZN(n1086) );
XOR2_X1 U780 ( .A(n1088), .B(G104), .Z(G6) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
OR2_X1 U782 ( .A1(n1091), .A2(KEYINPUT24), .ZN(n1090) );
NAND3_X1 U783 ( .A1(n1092), .A2(n1024), .A3(KEYINPUT24), .ZN(n1089) );
INV_X1 U784 ( .A(n1093), .ZN(n1024) );
NOR2_X1 U785 ( .A1(n1074), .A2(n1094), .ZN(G57) );
XOR2_X1 U786 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U787 ( .A(KEYINPUT14), .B(n1097), .ZN(n1095) );
NOR2_X1 U788 ( .A1(KEYINPUT17), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U789 ( .A(n1099), .B(n1100), .ZN(n1098) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U791 ( .A1(KEYINPUT20), .A2(n1103), .ZN(n1102) );
AND2_X1 U792 ( .A1(KEYINPUT6), .A2(n1103), .ZN(n1101) );
AND2_X1 U793 ( .A1(n1084), .A2(G472), .ZN(n1103) );
NOR2_X1 U794 ( .A1(n1074), .A2(n1104), .ZN(G54) );
XOR2_X1 U795 ( .A(n1105), .B(n1106), .Z(n1104) );
AND2_X1 U796 ( .A1(G469), .A2(n1084), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1107), .A2(KEYINPUT27), .ZN(n1105) );
XOR2_X1 U798 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U799 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U801 ( .A1(G140), .A2(n1114), .ZN(n1113) );
NAND2_X1 U802 ( .A1(KEYINPUT32), .A2(n1115), .ZN(n1110) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1108) );
NOR2_X1 U804 ( .A1(n1074), .A2(n1118), .ZN(G51) );
XOR2_X1 U805 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U806 ( .A(n1121), .B(KEYINPUT13), .Z(n1119) );
NAND2_X1 U807 ( .A1(n1084), .A2(n1122), .ZN(n1121) );
INV_X1 U808 ( .A(n1078), .ZN(n1084) );
NAND2_X1 U809 ( .A1(G902), .A2(n1123), .ZN(n1078) );
NAND2_X1 U810 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U811 ( .A(KEYINPUT38), .B(n992), .ZN(n1125) );
NAND4_X1 U812 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n992) );
AND4_X1 U813 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U816 ( .A1(n1022), .A2(n1138), .ZN(n1137) );
XNOR2_X1 U817 ( .A(KEYINPUT50), .B(n1011), .ZN(n1138) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1001), .ZN(n1136) );
XNOR2_X1 U819 ( .A(n1007), .B(KEYINPUT30), .ZN(n1139) );
NAND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1126) );
XOR2_X1 U821 ( .A(n1142), .B(KEYINPUT31), .Z(n1140) );
INV_X1 U822 ( .A(n993), .ZN(n1124) );
NAND2_X1 U823 ( .A1(n1069), .A2(n1071), .ZN(n993) );
AND4_X1 U824 ( .A1(n1143), .A2(n1144), .A3(n1091), .A4(n1145), .ZN(n1069) );
NOR4_X1 U825 ( .A1(n1146), .A2(n1147), .A3(n988), .A4(n1148), .ZN(n1145) );
AND4_X1 U826 ( .A1(n1093), .A2(n1149), .A3(n1022), .A4(n1009), .ZN(n988) );
NAND2_X1 U827 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND3_X1 U828 ( .A1(n1149), .A2(n1009), .A3(n1021), .ZN(n1092) );
NOR2_X1 U829 ( .A1(n995), .A2(G952), .ZN(n1074) );
XOR2_X1 U830 ( .A(n1127), .B(n1150), .Z(G48) );
XNOR2_X1 U831 ( .A(KEYINPUT36), .B(n1151), .ZN(n1150) );
NAND2_X1 U832 ( .A1(n1152), .A2(n1021), .ZN(n1127) );
XOR2_X1 U833 ( .A(G143), .B(n1153), .Z(G45) );
NOR2_X1 U834 ( .A1(n1011), .A2(n1142), .ZN(n1153) );
NAND4_X1 U835 ( .A1(n1154), .A2(n1155), .A3(n1008), .A4(n1035), .ZN(n1142) );
XNOR2_X1 U836 ( .A(n1156), .B(n1157), .ZN(G42) );
NOR2_X1 U837 ( .A1(KEYINPUT0), .A2(n1133), .ZN(n1157) );
NAND3_X1 U838 ( .A1(n1021), .A2(n1016), .A3(n1158), .ZN(n1133) );
XOR2_X1 U839 ( .A(G137), .B(n1159), .Z(G39) );
AND3_X1 U840 ( .A1(n1134), .A2(n1001), .A3(n1007), .ZN(n1159) );
INV_X1 U841 ( .A(n1160), .ZN(n1134) );
NAND3_X1 U842 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(G36) );
OR2_X1 U843 ( .A1(G134), .A2(KEYINPUT55), .ZN(n1163) );
NAND3_X1 U844 ( .A1(KEYINPUT55), .A2(G134), .A3(n1132), .ZN(n1162) );
NAND2_X1 U845 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
NAND2_X1 U846 ( .A1(KEYINPUT55), .A2(n1166), .ZN(n1165) );
XOR2_X1 U847 ( .A(KEYINPUT51), .B(G134), .Z(n1166) );
INV_X1 U848 ( .A(n1132), .ZN(n1164) );
NAND3_X1 U849 ( .A1(n1008), .A2(n1022), .A3(n1158), .ZN(n1132) );
XNOR2_X1 U850 ( .A(G131), .B(n1131), .ZN(G33) );
NAND3_X1 U851 ( .A1(n1021), .A2(n1008), .A3(n1158), .ZN(n1131) );
AND2_X1 U852 ( .A1(n1007), .A2(n1155), .ZN(n1158) );
NOR2_X1 U853 ( .A1(n1167), .A2(n1013), .ZN(n1007) );
XNOR2_X1 U854 ( .A(G128), .B(n1168), .ZN(G30) );
NAND2_X1 U855 ( .A1(n1152), .A2(n1022), .ZN(n1168) );
NOR2_X1 U856 ( .A1(n1160), .A2(n1011), .ZN(n1152) );
INV_X1 U857 ( .A(n1141), .ZN(n1011) );
NAND3_X1 U858 ( .A1(n1169), .A2(n1033), .A3(n1155), .ZN(n1160) );
AND2_X1 U859 ( .A1(n1093), .A2(n1170), .ZN(n1155) );
XNOR2_X1 U860 ( .A(G101), .B(n1171), .ZN(G3) );
NAND2_X1 U861 ( .A1(KEYINPUT47), .A2(n1147), .ZN(n1171) );
AND4_X1 U862 ( .A1(n1008), .A2(n1001), .A3(n1093), .A4(n1149), .ZN(n1147) );
XNOR2_X1 U863 ( .A(G125), .B(n1130), .ZN(G27) );
NAND3_X1 U864 ( .A1(n1021), .A2(n1003), .A3(n1172), .ZN(n1130) );
AND3_X1 U865 ( .A1(n1141), .A2(n1170), .A3(n1016), .ZN(n1172) );
NAND2_X1 U866 ( .A1(n1173), .A2(n1029), .ZN(n1170) );
NAND2_X1 U867 ( .A1(n1174), .A2(n1052), .ZN(n1173) );
XOR2_X1 U868 ( .A(G900), .B(KEYINPUT34), .Z(n1052) );
XNOR2_X1 U869 ( .A(G122), .B(n1143), .ZN(G24) );
NAND4_X1 U870 ( .A1(n1154), .A2(n1175), .A3(n1009), .A4(n1035), .ZN(n1143) );
XNOR2_X1 U871 ( .A(G119), .B(n1144), .ZN(G21) );
NAND4_X1 U872 ( .A1(n1175), .A2(n1001), .A3(n1169), .A4(n1033), .ZN(n1144) );
NAND2_X1 U873 ( .A1(n1176), .A2(n1177), .ZN(G18) );
NAND2_X1 U874 ( .A1(n1146), .A2(n1178), .ZN(n1177) );
XOR2_X1 U875 ( .A(KEYINPUT23), .B(n1179), .Z(n1176) );
NOR2_X1 U876 ( .A1(n1146), .A2(n1178), .ZN(n1179) );
AND3_X1 U877 ( .A1(n1008), .A2(n1022), .A3(n1175), .ZN(n1146) );
NOR2_X1 U878 ( .A1(n1180), .A2(n1154), .ZN(n1022) );
XOR2_X1 U879 ( .A(G113), .B(n1148), .Z(G15) );
AND3_X1 U880 ( .A1(n1175), .A2(n1008), .A3(n1021), .ZN(n1148) );
AND2_X1 U881 ( .A1(n1154), .A2(n1180), .ZN(n1021) );
INV_X1 U882 ( .A(n1035), .ZN(n1180) );
AND2_X1 U883 ( .A1(n1181), .A2(n1169), .ZN(n1008) );
AND2_X1 U884 ( .A1(n1003), .A2(n1149), .ZN(n1175) );
AND2_X1 U885 ( .A1(n1028), .A2(n1182), .ZN(n1003) );
XNOR2_X1 U886 ( .A(n1183), .B(n1071), .ZN(G12) );
NAND4_X1 U887 ( .A1(n1001), .A2(n1093), .A3(n1149), .A4(n1016), .ZN(n1071) );
NAND2_X1 U888 ( .A1(n1184), .A2(n1185), .ZN(n1016) );
NAND2_X1 U889 ( .A1(n1009), .A2(n1186), .ZN(n1185) );
NOR2_X1 U890 ( .A1(n1033), .A2(n1169), .ZN(n1009) );
OR3_X1 U891 ( .A1(n1181), .A2(n1169), .A3(n1186), .ZN(n1184) );
INV_X1 U892 ( .A(KEYINPUT54), .ZN(n1186) );
XNOR2_X1 U893 ( .A(n1042), .B(G472), .ZN(n1169) );
NAND2_X1 U894 ( .A1(n1187), .A2(n1188), .ZN(n1042) );
XOR2_X1 U895 ( .A(n1189), .B(n1096), .Z(n1187) );
XNOR2_X1 U896 ( .A(n1190), .B(G101), .ZN(n1096) );
NAND2_X1 U897 ( .A1(n1191), .A2(G210), .ZN(n1190) );
NAND2_X1 U898 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U899 ( .A1(KEYINPUT58), .A2(n1100), .ZN(n1193) );
XOR2_X1 U900 ( .A(n1194), .B(n1195), .Z(n1100) );
OR3_X1 U901 ( .A1(n1194), .A2(n1195), .A3(KEYINPUT58), .ZN(n1192) );
XOR2_X1 U902 ( .A(n1196), .B(n1056), .Z(n1194) );
INV_X1 U903 ( .A(n1033), .ZN(n1181) );
XOR2_X1 U904 ( .A(n1197), .B(n1077), .Z(n1033) );
NAND2_X1 U905 ( .A1(G217), .A2(n1198), .ZN(n1077) );
NAND2_X1 U906 ( .A1(n1188), .A2(n1079), .ZN(n1197) );
NAND2_X1 U907 ( .A1(n1199), .A2(n1200), .ZN(n1079) );
NAND3_X1 U908 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
XOR2_X1 U909 ( .A(n1204), .B(n1205), .Z(n1203) );
NAND2_X1 U910 ( .A1(n1206), .A2(n1207), .ZN(n1199) );
NAND2_X1 U911 ( .A1(n1201), .A2(n1202), .ZN(n1207) );
NAND2_X1 U912 ( .A1(n1208), .A2(n1209), .ZN(n1202) );
XNOR2_X1 U913 ( .A(G146), .B(n1210), .ZN(n1209) );
XOR2_X1 U914 ( .A(n1211), .B(n1212), .Z(n1208) );
XNOR2_X1 U915 ( .A(KEYINPUT49), .B(n1213), .ZN(n1201) );
NAND2_X1 U916 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U917 ( .A(n1211), .B(n1212), .ZN(n1215) );
XNOR2_X1 U918 ( .A(G128), .B(n1114), .ZN(n1212) );
NAND2_X1 U919 ( .A1(KEYINPUT35), .A2(G119), .ZN(n1211) );
XNOR2_X1 U920 ( .A(n1210), .B(n1151), .ZN(n1214) );
INV_X1 U921 ( .A(G146), .ZN(n1151) );
NAND2_X1 U922 ( .A1(KEYINPUT5), .A2(n1216), .ZN(n1210) );
XOR2_X1 U923 ( .A(G125), .B(n1217), .Z(n1216) );
NOR2_X1 U924 ( .A1(KEYINPUT4), .A2(n1218), .ZN(n1217) );
XNOR2_X1 U925 ( .A(KEYINPUT16), .B(G140), .ZN(n1218) );
XNOR2_X1 U926 ( .A(n1204), .B(n1205), .ZN(n1206) );
NOR2_X1 U927 ( .A1(n1219), .A2(n1220), .ZN(n1205) );
INV_X1 U928 ( .A(KEYINPUT48), .ZN(n1219) );
NAND3_X1 U929 ( .A1(G234), .A2(n1221), .A3(G221), .ZN(n1204) );
XNOR2_X1 U930 ( .A(KEYINPUT57), .B(n995), .ZN(n1221) );
AND2_X1 U931 ( .A1(n1141), .A2(n1222), .ZN(n1149) );
NAND2_X1 U932 ( .A1(n1029), .A2(n1223), .ZN(n1222) );
NAND2_X1 U933 ( .A1(n1174), .A2(n1064), .ZN(n1223) );
INV_X1 U934 ( .A(G898), .ZN(n1064) );
AND3_X1 U935 ( .A1(G902), .A2(n1224), .A3(G953), .ZN(n1174) );
NAND3_X1 U936 ( .A1(n1224), .A2(n995), .A3(G952), .ZN(n1029) );
NAND2_X1 U937 ( .A1(G237), .A2(n1225), .ZN(n1224) );
XOR2_X1 U938 ( .A(KEYINPUT43), .B(G234), .Z(n1225) );
NOR2_X1 U939 ( .A1(n1014), .A2(n1013), .ZN(n1141) );
AND2_X1 U940 ( .A1(G214), .A2(n1226), .ZN(n1013) );
XNOR2_X1 U941 ( .A(KEYINPUT12), .B(n1227), .ZN(n1226) );
INV_X1 U942 ( .A(n1167), .ZN(n1014) );
NAND3_X1 U943 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1167) );
NAND2_X1 U944 ( .A1(n1122), .A2(n1231), .ZN(n1230) );
OR3_X1 U945 ( .A1(n1231), .A2(n1122), .A3(n1232), .ZN(n1229) );
INV_X1 U946 ( .A(n1041), .ZN(n1122) );
NOR2_X1 U947 ( .A1(n1040), .A2(KEYINPUT62), .ZN(n1231) );
NAND2_X1 U948 ( .A1(n1233), .A2(n1232), .ZN(n1228) );
INV_X1 U949 ( .A(KEYINPUT2), .ZN(n1232) );
NAND2_X1 U950 ( .A1(n1040), .A2(n1041), .ZN(n1233) );
NAND2_X1 U951 ( .A1(G210), .A2(n1227), .ZN(n1041) );
OR2_X1 U952 ( .A1(G902), .A2(G237), .ZN(n1227) );
NOR2_X1 U953 ( .A1(n1120), .A2(G902), .ZN(n1040) );
XNOR2_X1 U954 ( .A(n1234), .B(n1235), .ZN(n1120) );
XOR2_X1 U955 ( .A(n1196), .B(n1065), .Z(n1235) );
XNOR2_X1 U956 ( .A(n1236), .B(n1237), .ZN(n1065) );
NAND2_X1 U957 ( .A1(KEYINPUT21), .A2(n1114), .ZN(n1236) );
XOR2_X1 U958 ( .A(n1238), .B(n1239), .Z(n1196) );
XNOR2_X1 U959 ( .A(n1240), .B(KEYINPUT3), .ZN(n1238) );
XOR2_X1 U960 ( .A(n1241), .B(n1242), .Z(n1234) );
XOR2_X1 U961 ( .A(G125), .B(n1243), .Z(n1242) );
NOR3_X1 U962 ( .A1(KEYINPUT25), .A2(n1244), .A3(n1245), .ZN(n1243) );
NOR3_X1 U963 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1245) );
AND2_X1 U964 ( .A1(n1246), .A2(n1067), .ZN(n1244) );
XOR2_X1 U965 ( .A(n1248), .B(n1247), .Z(n1067) );
XNOR2_X1 U966 ( .A(n1195), .B(KEYINPUT41), .ZN(n1247) );
XOR2_X1 U967 ( .A(G113), .B(n1249), .Z(n1195) );
XNOR2_X1 U968 ( .A(G119), .B(n1178), .ZN(n1249) );
INV_X1 U969 ( .A(G116), .ZN(n1178) );
NAND2_X1 U970 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
OR2_X1 U971 ( .A1(n1252), .A2(G101), .ZN(n1251) );
XOR2_X1 U972 ( .A(n1253), .B(KEYINPUT33), .Z(n1250) );
NAND2_X1 U973 ( .A1(G101), .A2(n1252), .ZN(n1253) );
INV_X1 U974 ( .A(KEYINPUT18), .ZN(n1246) );
NAND2_X1 U975 ( .A1(G224), .A2(n995), .ZN(n1241) );
NOR2_X1 U976 ( .A1(n1028), .A2(n1026), .ZN(n1093) );
INV_X1 U977 ( .A(n1182), .ZN(n1026) );
NAND2_X1 U978 ( .A1(G221), .A2(n1198), .ZN(n1182) );
NAND2_X1 U979 ( .A1(G234), .A2(n1188), .ZN(n1198) );
XOR2_X1 U980 ( .A(n1034), .B(KEYINPUT9), .Z(n1028) );
XNOR2_X1 U981 ( .A(n1254), .B(n1255), .ZN(n1034) );
XOR2_X1 U982 ( .A(KEYINPUT53), .B(G469), .Z(n1255) );
NAND2_X1 U983 ( .A1(n1256), .A2(n1188), .ZN(n1254) );
XNOR2_X1 U984 ( .A(n1115), .B(n1257), .ZN(n1256) );
XOR2_X1 U985 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U986 ( .A1(n1260), .A2(KEYINPUT1), .ZN(n1259) );
XOR2_X1 U987 ( .A(n1261), .B(n1116), .Z(n1260) );
XNOR2_X1 U988 ( .A(n1262), .B(n1056), .ZN(n1116) );
XNOR2_X1 U989 ( .A(n1263), .B(n1220), .ZN(n1056) );
XOR2_X1 U990 ( .A(G137), .B(KEYINPUT45), .Z(n1220) );
XNOR2_X1 U991 ( .A(G131), .B(G134), .ZN(n1263) );
XOR2_X1 U992 ( .A(n1055), .B(KEYINPUT8), .Z(n1262) );
NAND3_X1 U993 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1055) );
NAND2_X1 U994 ( .A1(KEYINPUT10), .A2(n1239), .ZN(n1266) );
NAND3_X1 U995 ( .A1(n1267), .A2(n1268), .A3(n1240), .ZN(n1265) );
INV_X1 U996 ( .A(KEYINPUT10), .ZN(n1268) );
OR2_X1 U997 ( .A1(n1240), .A2(n1267), .ZN(n1264) );
NOR2_X1 U998 ( .A1(KEYINPUT44), .A2(n1239), .ZN(n1267) );
XOR2_X1 U999 ( .A(G128), .B(KEYINPUT15), .Z(n1239) );
XOR2_X1 U1000 ( .A(G146), .B(n1269), .Z(n1240) );
NAND2_X1 U1001 ( .A1(KEYINPUT60), .A2(n1117), .ZN(n1261) );
XOR2_X1 U1002 ( .A(n1270), .B(n1252), .Z(n1117) );
XOR2_X1 U1003 ( .A(G104), .B(G107), .Z(n1252) );
NAND2_X1 U1004 ( .A1(n1271), .A2(KEYINPUT46), .ZN(n1270) );
XNOR2_X1 U1005 ( .A(G101), .B(KEYINPUT39), .ZN(n1271) );
NAND2_X1 U1006 ( .A1(n1272), .A2(n1112), .ZN(n1258) );
NAND2_X1 U1007 ( .A1(G110), .A2(n1156), .ZN(n1112) );
NAND2_X1 U1008 ( .A1(n1273), .A2(n1114), .ZN(n1272) );
XNOR2_X1 U1009 ( .A(KEYINPUT19), .B(n1156), .ZN(n1273) );
AND2_X1 U1010 ( .A1(G227), .A2(n995), .ZN(n1115) );
NOR2_X1 U1011 ( .A1(n1035), .A2(n1154), .ZN(n1001) );
XOR2_X1 U1012 ( .A(n1039), .B(n1274), .Z(n1154) );
NOR2_X1 U1013 ( .A1(G475), .A2(KEYINPUT28), .ZN(n1274) );
NAND2_X1 U1014 ( .A1(n1275), .A2(n1188), .ZN(n1039) );
XOR2_X1 U1015 ( .A(n1087), .B(KEYINPUT7), .Z(n1275) );
XOR2_X1 U1016 ( .A(n1276), .B(G113), .Z(n1087) );
XOR2_X1 U1017 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1018 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U1019 ( .A(n1237), .B(G104), .ZN(n1280) );
XOR2_X1 U1020 ( .A(KEYINPUT16), .B(G131), .Z(n1279) );
XOR2_X1 U1021 ( .A(n1281), .B(n1282), .Z(n1277) );
XOR2_X1 U1022 ( .A(n1269), .B(n1054), .Z(n1282) );
XNOR2_X1 U1023 ( .A(G125), .B(n1156), .ZN(n1054) );
INV_X1 U1024 ( .A(G140), .ZN(n1156) );
XOR2_X1 U1025 ( .A(n1283), .B(n1284), .Z(n1281) );
NOR2_X1 U1026 ( .A1(G146), .A2(KEYINPUT59), .ZN(n1284) );
NAND2_X1 U1027 ( .A1(n1191), .A2(G214), .ZN(n1283) );
NOR2_X1 U1028 ( .A1(G953), .A2(G237), .ZN(n1191) );
XNOR2_X1 U1029 ( .A(n1285), .B(G478), .ZN(n1035) );
NAND2_X1 U1030 ( .A1(n1083), .A2(n1188), .ZN(n1285) );
INV_X1 U1031 ( .A(G902), .ZN(n1188) );
XNOR2_X1 U1032 ( .A(n1286), .B(n1287), .ZN(n1083) );
XOR2_X1 U1033 ( .A(n1288), .B(n1269), .Z(n1287) );
XOR2_X1 U1034 ( .A(G143), .B(KEYINPUT61), .Z(n1269) );
AND3_X1 U1035 ( .A1(G217), .A2(n995), .A3(G234), .ZN(n1288) );
INV_X1 U1036 ( .A(G953), .ZN(n995) );
XOR2_X1 U1037 ( .A(n1289), .B(n1290), .Z(n1286) );
XOR2_X1 U1038 ( .A(G134), .B(G128), .Z(n1290) );
NAND2_X1 U1039 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
OR2_X1 U1040 ( .A1(n1293), .A2(G107), .ZN(n1292) );
XOR2_X1 U1041 ( .A(n1294), .B(KEYINPUT22), .Z(n1291) );
NAND2_X1 U1042 ( .A1(G107), .A2(n1293), .ZN(n1294) );
XNOR2_X1 U1043 ( .A(G116), .B(n1237), .ZN(n1293) );
INV_X1 U1044 ( .A(G122), .ZN(n1237) );
NAND2_X1 U1045 ( .A1(KEYINPUT11), .A2(n1114), .ZN(n1183) );
INV_X1 U1046 ( .A(G110), .ZN(n1114) );
endmodule


