//Key = 0100100000001100101101000110111111010001001111100110000011111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;

XOR2_X1 U718 ( .A(n1000), .B(n1001), .Z(G9) );
NOR2_X1 U719 ( .A1(KEYINPUT41), .A2(n1002), .ZN(n1001) );
NOR2_X1 U720 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR3_X1 U721 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NOR4_X1 U722 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1006) );
NOR2_X1 U723 ( .A1(n1012), .A2(n1013), .ZN(n1008) );
NOR2_X1 U724 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
INV_X1 U725 ( .A(n1016), .ZN(n1015) );
NOR2_X1 U726 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
NOR2_X1 U727 ( .A1(n1019), .A2(n1020), .ZN(n1012) );
INV_X1 U728 ( .A(n1021), .ZN(n1020) );
NOR2_X1 U729 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NOR2_X1 U730 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NAND3_X1 U731 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1005) );
NAND4_X1 U732 ( .A1(n1016), .A2(n1021), .A3(n1029), .A4(n1030), .ZN(n1028) );
NAND2_X1 U733 ( .A1(n1031), .A2(n1011), .ZN(n1030) );
NAND2_X1 U734 ( .A1(KEYINPUT15), .A2(n1032), .ZN(n1031) );
NAND4_X1 U735 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1029) );
INV_X1 U736 ( .A(n1011), .ZN(n1036) );
NAND2_X1 U737 ( .A1(n1032), .A2(n1037), .ZN(n1035) );
INV_X1 U738 ( .A(KEYINPUT15), .ZN(n1037) );
NAND3_X1 U739 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1034) );
NAND2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1033) );
OR2_X1 U741 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U742 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1003) );
INV_X1 U743 ( .A(n1026), .ZN(n1045) );
NAND4_X1 U744 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1026) );
NOR3_X1 U745 ( .A1(n1050), .A2(n1009), .A3(n1051), .ZN(n1049) );
NAND3_X1 U746 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1050) );
XOR2_X1 U747 ( .A(n1055), .B(KEYINPUT20), .Z(n1054) );
NAND2_X1 U748 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
OR2_X1 U749 ( .A1(n1058), .A2(KEYINPUT44), .ZN(n1053) );
NAND3_X1 U750 ( .A1(n1058), .A2(n1059), .A3(KEYINPUT44), .ZN(n1052) );
NOR3_X1 U751 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1060) );
XOR2_X1 U753 ( .A(n1063), .B(KEYINPUT13), .Z(n1056) );
XOR2_X1 U754 ( .A(n1064), .B(n1065), .Z(n1047) );
NAND2_X1 U755 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XNOR2_X1 U756 ( .A(KEYINPUT62), .B(KEYINPUT32), .ZN(n1066) );
XOR2_X1 U757 ( .A(n1068), .B(n1069), .Z(G72) );
XOR2_X1 U758 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U759 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U760 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U761 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U762 ( .A1(KEYINPUT46), .A2(n1078), .ZN(n1077) );
NOR2_X1 U763 ( .A1(G900), .A2(n1027), .ZN(n1072) );
NAND2_X1 U764 ( .A1(n1079), .A2(n1027), .ZN(n1070) );
NAND2_X1 U765 ( .A1(G953), .A2(n1080), .ZN(n1068) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1080) );
XOR2_X1 U767 ( .A(n1081), .B(n1082), .Z(G69) );
XOR2_X1 U768 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR3_X1 U769 ( .A1(n1085), .A2(KEYINPUT9), .A3(G953), .ZN(n1084) );
NOR2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U771 ( .A(n1088), .B(KEYINPUT59), .Z(n1086) );
NAND2_X1 U772 ( .A1(n1089), .A2(n1090), .ZN(n1083) );
NAND2_X1 U773 ( .A1(G953), .A2(n1091), .ZN(n1090) );
XOR2_X1 U774 ( .A(n1092), .B(KEYINPUT39), .Z(n1089) );
NAND2_X1 U775 ( .A1(G953), .A2(n1093), .ZN(n1081) );
NAND2_X1 U776 ( .A1(G898), .A2(G224), .ZN(n1093) );
NOR2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(G66) );
XOR2_X1 U778 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1100), .ZN(G63) );
NOR3_X1 U781 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
AND3_X1 U782 ( .A1(n1104), .A2(G478), .A3(n1105), .ZN(n1103) );
NOR2_X1 U783 ( .A1(n1106), .A2(n1104), .ZN(n1102) );
NOR2_X1 U784 ( .A1(n1107), .A2(n1064), .ZN(n1106) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1108), .ZN(G60) );
XOR2_X1 U786 ( .A(n1109), .B(n1110), .Z(n1108) );
AND2_X1 U787 ( .A1(G475), .A2(n1105), .ZN(n1109) );
XOR2_X1 U788 ( .A(G104), .B(n1111), .Z(G6) );
NOR3_X1 U789 ( .A1(n1094), .A2(n1112), .A3(n1113), .ZN(G57) );
NOR2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
AND2_X1 U792 ( .A1(KEYINPUT34), .A2(n1118), .ZN(n1117) );
NOR3_X1 U793 ( .A1(KEYINPUT34), .A2(n1118), .A3(n1119), .ZN(n1116) );
INV_X1 U794 ( .A(n1120), .ZN(n1114) );
NOR2_X1 U795 ( .A1(n1121), .A2(n1120), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1122), .B(n1123), .Z(n1120) );
NOR2_X1 U797 ( .A1(KEYINPUT54), .A2(n1124), .ZN(n1123) );
NAND2_X1 U798 ( .A1(n1105), .A2(G472), .ZN(n1122) );
NOR2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1121) );
INV_X1 U800 ( .A(KEYINPUT29), .ZN(n1119) );
XNOR2_X1 U801 ( .A(n1125), .B(G101), .ZN(n1118) );
NOR2_X1 U802 ( .A1(n1094), .A2(n1126), .ZN(G54) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U804 ( .A1(n1105), .A2(G469), .ZN(n1128) );
INV_X1 U805 ( .A(n1099), .ZN(n1105) );
NAND2_X1 U806 ( .A1(KEYINPUT57), .A2(n1129), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U808 ( .A1(n1094), .A2(n1132), .ZN(G51) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U810 ( .A1(n1057), .A2(n1099), .ZN(n1133) );
NAND2_X1 U811 ( .A1(G902), .A2(n1007), .ZN(n1099) );
INV_X1 U812 ( .A(n1107), .ZN(n1007) );
NOR3_X1 U813 ( .A1(n1079), .A2(n1111), .A3(n1087), .ZN(n1107) );
NAND4_X1 U814 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1087) );
NOR4_X1 U815 ( .A1(n1000), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1138) );
INV_X1 U816 ( .A(n1142), .ZN(n1141) );
AND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1000) );
NAND3_X1 U818 ( .A1(n1145), .A2(n1146), .A3(n1039), .ZN(n1137) );
XNOR2_X1 U819 ( .A(KEYINPUT47), .B(n1147), .ZN(n1146) );
NAND4_X1 U820 ( .A1(n1018), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1135) );
XOR2_X1 U821 ( .A(KEYINPUT24), .B(n1039), .Z(n1150) );
INV_X1 U822 ( .A(n1088), .ZN(n1111) );
NAND3_X1 U823 ( .A1(n1144), .A2(n1149), .A3(n1043), .ZN(n1088) );
AND2_X1 U824 ( .A1(n1148), .A2(n1021), .ZN(n1144) );
NAND4_X1 U825 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1079) );
AND4_X1 U826 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
NAND3_X1 U827 ( .A1(n1159), .A2(n1044), .A3(n1016), .ZN(n1153) );
NAND3_X1 U828 ( .A1(n1023), .A2(n1160), .A3(n1161), .ZN(n1151) );
OR2_X1 U829 ( .A1(n1162), .A2(n1143), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1027), .A2(G952), .ZN(n1094) );
XOR2_X1 U831 ( .A(n1163), .B(n1164), .Z(G48) );
NAND3_X1 U832 ( .A1(n1162), .A2(n1161), .A3(n1165), .ZN(n1164) );
XNOR2_X1 U833 ( .A(n1023), .B(KEYINPUT31), .ZN(n1165) );
AND2_X1 U834 ( .A1(n1166), .A2(n1043), .ZN(n1162) );
XOR2_X1 U835 ( .A(n1152), .B(n1167), .Z(G45) );
XOR2_X1 U836 ( .A(KEYINPUT19), .B(G143), .Z(n1167) );
NAND4_X1 U837 ( .A1(n1159), .A2(n1023), .A3(n1168), .A4(n1169), .ZN(n1152) );
XNOR2_X1 U838 ( .A(G140), .B(n1158), .ZN(G42) );
NAND3_X1 U839 ( .A1(n1166), .A2(n1170), .A3(n1016), .ZN(n1158) );
XNOR2_X1 U840 ( .A(G137), .B(n1157), .ZN(G39) );
NAND3_X1 U841 ( .A1(n1032), .A2(n1016), .A3(n1161), .ZN(n1157) );
AND2_X1 U842 ( .A1(n1166), .A2(n1039), .ZN(n1032) );
XOR2_X1 U843 ( .A(G134), .B(n1171), .Z(G36) );
NOR3_X1 U844 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
XOR2_X1 U845 ( .A(KEYINPUT4), .B(n1016), .Z(n1172) );
XNOR2_X1 U846 ( .A(G131), .B(n1156), .ZN(G33) );
NAND3_X1 U847 ( .A1(n1159), .A2(n1043), .A3(n1016), .ZN(n1156) );
NOR2_X1 U848 ( .A1(n1024), .A2(n1062), .ZN(n1016) );
INV_X1 U849 ( .A(n1025), .ZN(n1062) );
INV_X1 U850 ( .A(n1174), .ZN(n1159) );
NAND3_X1 U851 ( .A1(n1017), .A2(n1175), .A3(n1166), .ZN(n1174) );
XNOR2_X1 U852 ( .A(n1149), .B(KEYINPUT42), .ZN(n1166) );
XOR2_X1 U853 ( .A(n1176), .B(n1177), .Z(G30) );
NAND3_X1 U854 ( .A1(n1143), .A2(n1178), .A3(n1161), .ZN(n1177) );
NOR2_X1 U855 ( .A1(n1147), .A2(n1179), .ZN(n1161) );
INV_X1 U856 ( .A(n1175), .ZN(n1179) );
XOR2_X1 U857 ( .A(KEYINPUT11), .B(n1023), .Z(n1178) );
AND2_X1 U858 ( .A1(n1149), .A2(n1044), .ZN(n1143) );
INV_X1 U859 ( .A(n1173), .ZN(n1044) );
XNOR2_X1 U860 ( .A(n1136), .B(n1180), .ZN(G3) );
XOR2_X1 U861 ( .A(KEYINPUT17), .B(G101), .Z(n1180) );
OR2_X1 U862 ( .A1(n1181), .A2(n1182), .ZN(n1136) );
NAND2_X1 U863 ( .A1(n1183), .A2(n1184), .ZN(G27) );
NAND2_X1 U864 ( .A1(G125), .A2(n1155), .ZN(n1184) );
XOR2_X1 U865 ( .A(KEYINPUT25), .B(n1185), .Z(n1183) );
NOR2_X1 U866 ( .A1(G125), .A2(n1155), .ZN(n1185) );
NAND3_X1 U867 ( .A1(n1041), .A2(n1023), .A3(n1170), .ZN(n1155) );
AND3_X1 U868 ( .A1(n1043), .A2(n1175), .A3(n1018), .ZN(n1170) );
INV_X1 U869 ( .A(n1186), .ZN(n1018) );
NAND2_X1 U870 ( .A1(n1011), .A2(n1187), .ZN(n1175) );
NAND4_X1 U871 ( .A1(G902), .A2(G953), .A3(n1188), .A4(n1189), .ZN(n1187) );
INV_X1 U872 ( .A(G900), .ZN(n1189) );
XOR2_X1 U873 ( .A(G122), .B(n1190), .Z(G24) );
NOR2_X1 U874 ( .A1(KEYINPUT53), .A2(n1142), .ZN(n1190) );
NAND4_X1 U875 ( .A1(n1145), .A2(n1021), .A3(n1168), .A4(n1169), .ZN(n1142) );
INV_X1 U876 ( .A(n1046), .ZN(n1168) );
NOR2_X1 U877 ( .A1(n1191), .A2(n1051), .ZN(n1021) );
XOR2_X1 U878 ( .A(G119), .B(n1192), .Z(G21) );
NOR3_X1 U879 ( .A1(n1147), .A2(n1193), .A3(n1010), .ZN(n1192) );
NAND2_X1 U880 ( .A1(n1051), .A2(n1191), .ZN(n1147) );
INV_X1 U881 ( .A(n1194), .ZN(n1051) );
XOR2_X1 U882 ( .A(G116), .B(n1140), .Z(G18) );
NOR3_X1 U883 ( .A1(n1193), .A2(n1173), .A3(n1182), .ZN(n1140) );
INV_X1 U884 ( .A(n1017), .ZN(n1182) );
NAND2_X1 U885 ( .A1(n1046), .A2(n1169), .ZN(n1173) );
NAND2_X1 U886 ( .A1(n1195), .A2(n1196), .ZN(G15) );
NAND2_X1 U887 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
INV_X1 U888 ( .A(G113), .ZN(n1198) );
NAND2_X1 U889 ( .A1(G113), .A2(n1199), .ZN(n1195) );
NAND2_X1 U890 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U891 ( .A1(n1139), .A2(n1202), .ZN(n1201) );
INV_X1 U892 ( .A(n1203), .ZN(n1139) );
OR2_X1 U893 ( .A1(n1202), .A2(n1197), .ZN(n1200) );
NOR2_X1 U894 ( .A1(KEYINPUT27), .A2(n1203), .ZN(n1197) );
NAND3_X1 U895 ( .A1(n1145), .A2(n1043), .A3(n1017), .ZN(n1203) );
NOR2_X1 U896 ( .A1(n1191), .A2(n1194), .ZN(n1017) );
NOR2_X1 U897 ( .A1(n1169), .A2(n1046), .ZN(n1043) );
INV_X1 U898 ( .A(n1193), .ZN(n1145) );
NAND2_X1 U899 ( .A1(n1041), .A2(n1148), .ZN(n1193) );
INV_X1 U900 ( .A(n1009), .ZN(n1041) );
NAND2_X1 U901 ( .A1(n1038), .A2(n1204), .ZN(n1009) );
INV_X1 U902 ( .A(KEYINPUT30), .ZN(n1202) );
XOR2_X1 U903 ( .A(G110), .B(n1205), .Z(G12) );
NOR2_X1 U904 ( .A1(n1181), .A2(n1186), .ZN(n1205) );
NAND2_X1 U905 ( .A1(n1194), .A2(n1191), .ZN(n1186) );
NAND3_X1 U906 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1191) );
INV_X1 U907 ( .A(n1061), .ZN(n1208) );
NOR2_X1 U908 ( .A1(n1059), .A2(n1058), .ZN(n1061) );
OR2_X1 U909 ( .A1(n1058), .A2(KEYINPUT49), .ZN(n1207) );
NAND3_X1 U910 ( .A1(n1058), .A2(n1059), .A3(KEYINPUT49), .ZN(n1206) );
OR2_X1 U911 ( .A1(n1097), .A2(G902), .ZN(n1059) );
XNOR2_X1 U912 ( .A(n1209), .B(n1210), .ZN(n1097) );
XOR2_X1 U913 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U914 ( .A(G128), .B(G119), .Z(n1212) );
NOR2_X1 U915 ( .A1(KEYINPUT6), .A2(G110), .ZN(n1211) );
XNOR2_X1 U916 ( .A(n1213), .B(n1214), .ZN(n1209) );
XOR2_X1 U917 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND3_X1 U918 ( .A1(G234), .A2(n1027), .A3(G221), .ZN(n1216) );
NAND2_X1 U919 ( .A1(n1217), .A2(KEYINPUT33), .ZN(n1215) );
XOR2_X1 U920 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U921 ( .A(KEYINPUT51), .B(KEYINPUT45), .Z(n1219) );
XOR2_X1 U922 ( .A(n1163), .B(n1220), .Z(n1218) );
INV_X1 U923 ( .A(n1098), .ZN(n1058) );
NAND2_X1 U924 ( .A1(G217), .A2(n1221), .ZN(n1098) );
XOR2_X1 U925 ( .A(n1222), .B(G472), .Z(n1194) );
NAND2_X1 U926 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U927 ( .A(n1225), .B(n1226), .Z(n1223) );
XNOR2_X1 U928 ( .A(n1227), .B(n1124), .ZN(n1226) );
XNOR2_X1 U929 ( .A(n1228), .B(n1229), .ZN(n1124) );
XOR2_X1 U930 ( .A(n1230), .B(n1231), .Z(n1229) );
XNOR2_X1 U931 ( .A(G116), .B(G119), .ZN(n1231) );
XOR2_X1 U932 ( .A(n1232), .B(n1233), .Z(n1228) );
NOR2_X1 U933 ( .A1(G113), .A2(KEYINPUT36), .ZN(n1233) );
NAND2_X1 U934 ( .A1(KEYINPUT28), .A2(n1234), .ZN(n1227) );
XOR2_X1 U935 ( .A(n1125), .B(n1235), .Z(n1225) );
XNOR2_X1 U936 ( .A(KEYINPUT38), .B(KEYINPUT22), .ZN(n1235) );
NAND2_X1 U937 ( .A1(G210), .A2(n1236), .ZN(n1125) );
NAND3_X1 U938 ( .A1(n1148), .A2(n1149), .A3(n1039), .ZN(n1181) );
INV_X1 U939 ( .A(n1010), .ZN(n1039) );
NAND2_X1 U940 ( .A1(n1237), .A2(n1046), .ZN(n1010) );
XOR2_X1 U941 ( .A(n1238), .B(G475), .Z(n1046) );
OR2_X1 U942 ( .A1(n1110), .A2(G902), .ZN(n1238) );
XNOR2_X1 U943 ( .A(n1239), .B(n1240), .ZN(n1110) );
XOR2_X1 U944 ( .A(G122), .B(n1241), .Z(n1240) );
NOR2_X1 U945 ( .A1(KEYINPUT0), .A2(n1242), .ZN(n1241) );
XOR2_X1 U946 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U947 ( .A(n1074), .B(n1245), .Z(n1244) );
AND2_X1 U948 ( .A1(n1236), .A2(G214), .ZN(n1245) );
NOR2_X1 U949 ( .A1(G953), .A2(G237), .ZN(n1236) );
XNOR2_X1 U950 ( .A(G131), .B(n1220), .ZN(n1074) );
XOR2_X1 U951 ( .A(G140), .B(G125), .Z(n1220) );
XOR2_X1 U952 ( .A(n1246), .B(n1247), .Z(n1243) );
XOR2_X1 U953 ( .A(KEYINPUT37), .B(G146), .Z(n1247) );
XNOR2_X1 U954 ( .A(n1248), .B(n1249), .ZN(n1239) );
NOR2_X1 U955 ( .A1(G113), .A2(KEYINPUT23), .ZN(n1249) );
NOR2_X1 U956 ( .A1(G104), .A2(KEYINPUT5), .ZN(n1248) );
INV_X1 U957 ( .A(n1169), .ZN(n1237) );
NAND3_X1 U958 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1169) );
NAND2_X1 U959 ( .A1(G478), .A2(n1067), .ZN(n1252) );
NAND2_X1 U960 ( .A1(KEYINPUT8), .A2(n1253), .ZN(n1251) );
NAND2_X1 U961 ( .A1(n1254), .A2(n1064), .ZN(n1253) );
XOR2_X1 U962 ( .A(n1067), .B(KEYINPUT50), .Z(n1254) );
INV_X1 U963 ( .A(n1101), .ZN(n1067) );
NAND2_X1 U964 ( .A1(n1255), .A2(n1256), .ZN(n1250) );
INV_X1 U965 ( .A(KEYINPUT8), .ZN(n1256) );
NAND2_X1 U966 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
OR2_X1 U967 ( .A1(n1101), .A2(KEYINPUT50), .ZN(n1258) );
NAND3_X1 U968 ( .A1(n1101), .A2(n1064), .A3(KEYINPUT50), .ZN(n1257) );
INV_X1 U969 ( .A(G478), .ZN(n1064) );
NOR2_X1 U970 ( .A1(n1104), .A2(G902), .ZN(n1101) );
XNOR2_X1 U971 ( .A(n1259), .B(n1260), .ZN(n1104) );
XOR2_X1 U972 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U973 ( .A(G122), .B(n1263), .Z(n1262) );
AND3_X1 U974 ( .A1(n1264), .A2(G234), .A3(G217), .ZN(n1263) );
XOR2_X1 U975 ( .A(KEYINPUT61), .B(n1027), .Z(n1264) );
XOR2_X1 U976 ( .A(G134), .B(G128), .Z(n1261) );
XNOR2_X1 U977 ( .A(n1265), .B(n1266), .ZN(n1259) );
XNOR2_X1 U978 ( .A(n1267), .B(n1268), .ZN(n1266) );
NOR2_X1 U979 ( .A1(G143), .A2(KEYINPUT40), .ZN(n1268) );
NAND2_X1 U980 ( .A1(n1269), .A2(KEYINPUT56), .ZN(n1267) );
XNOR2_X1 U981 ( .A(G116), .B(KEYINPUT55), .ZN(n1269) );
NOR2_X1 U982 ( .A1(n1038), .A2(n1040), .ZN(n1149) );
INV_X1 U983 ( .A(n1204), .ZN(n1040) );
NAND2_X1 U984 ( .A1(G221), .A2(n1221), .ZN(n1204) );
NAND2_X1 U985 ( .A1(G234), .A2(n1224), .ZN(n1221) );
XOR2_X1 U986 ( .A(n1270), .B(G469), .Z(n1038) );
NAND2_X1 U987 ( .A1(n1271), .A2(n1224), .ZN(n1270) );
XOR2_X1 U988 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U989 ( .A(n1131), .B(n1274), .Z(n1273) );
NOR2_X1 U990 ( .A1(KEYINPUT63), .A2(n1130), .ZN(n1274) );
INV_X1 U991 ( .A(G110), .ZN(n1130) );
XOR2_X1 U992 ( .A(n1275), .B(n1276), .Z(n1131) );
XOR2_X1 U993 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U994 ( .A(n1076), .B(n1279), .Z(n1278) );
NAND2_X1 U995 ( .A1(KEYINPUT1), .A2(n1280), .ZN(n1279) );
XOR2_X1 U996 ( .A(KEYINPUT48), .B(n1281), .Z(n1280) );
INV_X1 U997 ( .A(n1282), .ZN(n1281) );
NAND3_X1 U998 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1076) );
NAND2_X1 U999 ( .A1(n1286), .A2(n1163), .ZN(n1284) );
XOR2_X1 U1000 ( .A(n1287), .B(G128), .Z(n1286) );
NAND2_X1 U1001 ( .A1(n1288), .A2(G146), .ZN(n1283) );
NAND2_X1 U1002 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
OR2_X1 U1003 ( .A1(n1287), .A2(G128), .ZN(n1290) );
NAND2_X1 U1004 ( .A1(KEYINPUT58), .A2(G143), .ZN(n1287) );
OR2_X1 U1005 ( .A1(n1176), .A2(KEYINPUT58), .ZN(n1289) );
XOR2_X1 U1006 ( .A(KEYINPUT16), .B(G140), .Z(n1277) );
XOR2_X1 U1007 ( .A(n1291), .B(n1292), .Z(n1275) );
XOR2_X1 U1008 ( .A(n1232), .B(n1293), .Z(n1291) );
AND2_X1 U1009 ( .A1(n1027), .A2(G227), .ZN(n1293) );
XOR2_X1 U1010 ( .A(n1078), .B(G131), .Z(n1232) );
XNOR2_X1 U1011 ( .A(G134), .B(n1213), .ZN(n1078) );
XOR2_X1 U1012 ( .A(G137), .B(KEYINPUT52), .Z(n1213) );
XNOR2_X1 U1013 ( .A(KEYINPUT7), .B(KEYINPUT21), .ZN(n1272) );
AND2_X1 U1014 ( .A1(n1023), .A2(n1294), .ZN(n1148) );
NAND2_X1 U1015 ( .A1(n1011), .A2(n1295), .ZN(n1294) );
NAND4_X1 U1016 ( .A1(G902), .A2(G953), .A3(n1188), .A4(n1091), .ZN(n1295) );
INV_X1 U1017 ( .A(G898), .ZN(n1091) );
NAND3_X1 U1018 ( .A1(n1188), .A2(n1027), .A3(G952), .ZN(n1011) );
NAND2_X1 U1019 ( .A1(G237), .A2(G234), .ZN(n1188) );
AND2_X1 U1020 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1296), .ZN(n1025) );
XNOR2_X1 U1022 ( .A(n1297), .B(n1057), .ZN(n1024) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1296), .ZN(n1057) );
NAND2_X1 U1024 ( .A1(n1298), .A2(n1224), .ZN(n1296) );
INV_X1 U1025 ( .A(G237), .ZN(n1298) );
XOR2_X1 U1026 ( .A(n1063), .B(KEYINPUT26), .Z(n1297) );
NAND2_X1 U1027 ( .A1(n1299), .A2(n1224), .ZN(n1063) );
INV_X1 U1028 ( .A(G902), .ZN(n1224) );
XNOR2_X1 U1029 ( .A(n1134), .B(n1300), .ZN(n1299) );
XNOR2_X1 U1030 ( .A(KEYINPUT2), .B(KEYINPUT18), .ZN(n1300) );
XNOR2_X1 U1031 ( .A(n1301), .B(n1302), .ZN(n1134) );
XOR2_X1 U1032 ( .A(n1230), .B(n1303), .Z(n1302) );
XNOR2_X1 U1033 ( .A(G125), .B(KEYINPUT14), .ZN(n1303) );
NAND3_X1 U1034 ( .A1(n1304), .A2(n1305), .A3(n1285), .ZN(n1230) );
NAND3_X1 U1035 ( .A1(G128), .A2(n1246), .A3(G146), .ZN(n1285) );
INV_X1 U1036 ( .A(G143), .ZN(n1246) );
NAND2_X1 U1037 ( .A1(n1306), .A2(n1163), .ZN(n1305) );
INV_X1 U1038 ( .A(G146), .ZN(n1163) );
XOR2_X1 U1039 ( .A(G128), .B(n1307), .Z(n1306) );
XOR2_X1 U1040 ( .A(KEYINPUT35), .B(G143), .Z(n1307) );
NAND3_X1 U1041 ( .A1(G143), .A2(n1176), .A3(G146), .ZN(n1304) );
INV_X1 U1042 ( .A(G128), .ZN(n1176) );
XOR2_X1 U1043 ( .A(n1092), .B(n1308), .Z(n1301) );
AND2_X1 U1044 ( .A1(n1027), .A2(G224), .ZN(n1308) );
INV_X1 U1045 ( .A(G953), .ZN(n1027) );
XOR2_X1 U1046 ( .A(n1309), .B(n1310), .Z(n1092) );
XOR2_X1 U1047 ( .A(G110), .B(n1311), .Z(n1310) );
XOR2_X1 U1048 ( .A(G122), .B(G113), .Z(n1311) );
XOR2_X1 U1049 ( .A(n1312), .B(n1313), .Z(n1309) );
XOR2_X1 U1050 ( .A(n1314), .B(n1282), .Z(n1313) );
XOR2_X1 U1051 ( .A(n1234), .B(KEYINPUT12), .Z(n1282) );
INV_X1 U1052 ( .A(G101), .ZN(n1234) );
NAND2_X1 U1053 ( .A1(n1315), .A2(KEYINPUT60), .ZN(n1314) );
XNOR2_X1 U1054 ( .A(G116), .B(n1316), .ZN(n1315) );
NOR2_X1 U1055 ( .A1(G119), .A2(KEYINPUT3), .ZN(n1316) );
NAND2_X1 U1056 ( .A1(n1317), .A2(n1318), .ZN(n1312) );
NAND2_X1 U1057 ( .A1(n1292), .A2(n1319), .ZN(n1318) );
INV_X1 U1058 ( .A(KEYINPUT10), .ZN(n1319) );
XOR2_X1 U1059 ( .A(G104), .B(n1265), .Z(n1292) );
NAND3_X1 U1060 ( .A1(G104), .A2(n1265), .A3(KEYINPUT10), .ZN(n1317) );
XNOR2_X1 U1061 ( .A(n1002), .B(KEYINPUT43), .ZN(n1265) );
INV_X1 U1062 ( .A(G107), .ZN(n1002) );
endmodule


