//Key = 0101100001010000001110110100000010001011011001111011110000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315;

XNOR2_X1 U733 ( .A(G107), .B(n991), .ZN(G9) );
NOR2_X1 U734 ( .A1(n992), .A2(n993), .ZN(G75) );
NOR3_X1 U735 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n993) );
NOR2_X1 U736 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U737 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U738 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NOR2_X1 U739 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U740 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U741 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U742 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR3_X1 U743 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1009) );
AND2_X1 U744 ( .A1(n1014), .A2(KEYINPUT24), .ZN(n1013) );
NOR3_X1 U745 ( .A1(KEYINPUT24), .A2(n1015), .A3(n1014), .ZN(n1012) );
NOR2_X1 U746 ( .A1(n1016), .A2(n1017), .ZN(n1007) );
NOR2_X1 U747 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U748 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR3_X1 U749 ( .A1(n1010), .A2(n1022), .A3(n1017), .ZN(n1003) );
INV_X1 U750 ( .A(n1023), .ZN(n1017) );
NOR2_X1 U751 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U752 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
AND4_X1 U753 ( .A1(n1028), .A2(n1029), .A3(n1023), .A4(n1030), .ZN(n999) );
NAND3_X1 U754 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n994) );
NAND3_X1 U755 ( .A1(n1034), .A2(n1023), .A3(n1035), .ZN(n1033) );
NOR3_X1 U756 ( .A1(n1036), .A2(n1037), .A3(n1006), .ZN(n1035) );
XOR2_X1 U757 ( .A(n998), .B(KEYINPUT21), .Z(n1037) );
XOR2_X1 U758 ( .A(n1010), .B(KEYINPUT36), .Z(n1034) );
NOR3_X1 U759 ( .A1(n1038), .A2(G953), .A3(G952), .ZN(n992) );
INV_X1 U760 ( .A(n1031), .ZN(n1038) );
NAND2_X1 U761 ( .A1(n1039), .A2(n1040), .ZN(n1031) );
AND4_X1 U762 ( .A1(n1041), .A2(n1042), .A3(n1021), .A4(n1014), .ZN(n1040) );
NOR4_X1 U763 ( .A1(n1043), .A2(n1044), .A3(n1002), .A4(n1015), .ZN(n1039) );
NOR2_X1 U764 ( .A1(KEYINPUT18), .A2(n1045), .ZN(n1044) );
NOR3_X1 U765 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
AND2_X1 U766 ( .A1(n1006), .A2(KEYINPUT18), .ZN(n1043) );
XOR2_X1 U767 ( .A(n1049), .B(n1050), .Z(G72) );
XOR2_X1 U768 ( .A(n1051), .B(n1052), .Z(n1050) );
NOR3_X1 U769 ( .A1(n1053), .A2(KEYINPUT28), .A3(G953), .ZN(n1052) );
NOR2_X1 U770 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
XOR2_X1 U771 ( .A(n1056), .B(n1057), .Z(n1055) );
XNOR2_X1 U772 ( .A(n1058), .B(n1059), .ZN(n1057) );
XOR2_X1 U773 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR2_X1 U774 ( .A1(G134), .A2(KEYINPUT37), .ZN(n1060) );
XOR2_X1 U775 ( .A(n1062), .B(n1063), .Z(n1056) );
NOR2_X1 U776 ( .A1(KEYINPUT30), .A2(G125), .ZN(n1063) );
XOR2_X1 U777 ( .A(n1064), .B(KEYINPUT38), .Z(n1062) );
NOR2_X1 U778 ( .A1(G900), .A2(n1065), .ZN(n1054) );
XOR2_X1 U779 ( .A(KEYINPUT1), .B(G953), .Z(n1065) );
NOR2_X1 U780 ( .A1(n1066), .A2(n1032), .ZN(n1049) );
NOR2_X1 U781 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U782 ( .A(n1069), .B(n1070), .Z(G69) );
XOR2_X1 U783 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U784 ( .A1(G953), .A2(n1073), .ZN(n1072) );
NOR2_X1 U785 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U786 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U787 ( .A1(G953), .A2(n1078), .ZN(n1077) );
XOR2_X1 U788 ( .A(n1079), .B(n1080), .Z(n1076) );
NAND2_X1 U789 ( .A1(KEYINPUT39), .A2(n1081), .ZN(n1079) );
NAND2_X1 U790 ( .A1(G953), .A2(n1082), .ZN(n1069) );
NAND2_X1 U791 ( .A1(G224), .A2(G898), .ZN(n1082) );
NOR2_X1 U792 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XNOR2_X1 U793 ( .A(n1085), .B(n1086), .ZN(n1084) );
NOR2_X1 U794 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U795 ( .A1(n1083), .A2(n1089), .ZN(G63) );
XOR2_X1 U796 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U797 ( .A1(n1092), .A2(n1088), .ZN(n1090) );
INV_X1 U798 ( .A(G478), .ZN(n1092) );
NOR2_X1 U799 ( .A1(n1093), .A2(n1094), .ZN(G60) );
XOR2_X1 U800 ( .A(KEYINPUT35), .B(n1083), .Z(n1094) );
XOR2_X1 U801 ( .A(n1095), .B(n1096), .Z(n1093) );
NOR2_X1 U802 ( .A1(n1097), .A2(n1088), .ZN(n1095) );
INV_X1 U803 ( .A(G475), .ZN(n1097) );
XNOR2_X1 U804 ( .A(G104), .B(n1098), .ZN(G6) );
NOR3_X1 U805 ( .A1(n1083), .A2(n1099), .A3(n1100), .ZN(G57) );
NOR2_X1 U806 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U807 ( .A(n1103), .B(n1104), .Z(n1102) );
OR2_X1 U808 ( .A1(n1105), .A2(KEYINPUT33), .ZN(n1103) );
NOR2_X1 U809 ( .A1(G101), .A2(n1106), .ZN(n1099) );
XOR2_X1 U810 ( .A(n1107), .B(n1104), .Z(n1106) );
XOR2_X1 U811 ( .A(n1108), .B(n1109), .Z(n1104) );
XOR2_X1 U812 ( .A(n1110), .B(n1111), .Z(n1108) );
NOR2_X1 U813 ( .A1(n1048), .A2(n1088), .ZN(n1111) );
INV_X1 U814 ( .A(G472), .ZN(n1048) );
NAND2_X1 U815 ( .A1(n1112), .A2(n1105), .ZN(n1107) );
INV_X1 U816 ( .A(KEYINPUT33), .ZN(n1112) );
NOR2_X1 U817 ( .A1(n1083), .A2(n1113), .ZN(G54) );
XOR2_X1 U818 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U819 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U820 ( .A1(n1118), .A2(n1088), .ZN(n1117) );
NOR3_X1 U821 ( .A1(KEYINPUT34), .A2(n1119), .A3(n1120), .ZN(n1116) );
AND2_X1 U822 ( .A1(n1121), .A2(KEYINPUT15), .ZN(n1120) );
NOR2_X1 U823 ( .A1(KEYINPUT15), .A2(n1122), .ZN(n1119) );
XOR2_X1 U824 ( .A(n1123), .B(n1124), .Z(n1114) );
XOR2_X1 U825 ( .A(KEYINPUT8), .B(n1125), .Z(n1124) );
NOR2_X1 U826 ( .A1(KEYINPUT60), .A2(n1126), .ZN(n1123) );
XOR2_X1 U827 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U828 ( .A(n1129), .B(n1130), .Z(n1127) );
NOR2_X1 U829 ( .A1(n1083), .A2(n1131), .ZN(G51) );
XOR2_X1 U830 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U831 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR3_X1 U832 ( .A1(n1088), .A2(KEYINPUT7), .A3(n1136), .ZN(n1135) );
NAND2_X1 U833 ( .A1(G902), .A2(n996), .ZN(n1088) );
NAND3_X1 U834 ( .A1(n1137), .A2(n1138), .A3(n1053), .ZN(n996) );
AND4_X1 U835 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1053) );
AND4_X1 U836 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
AND2_X1 U837 ( .A1(n1147), .A2(n1148), .ZN(n1141) );
XOR2_X1 U838 ( .A(KEYINPUT48), .B(n1074), .Z(n1138) );
INV_X1 U839 ( .A(n1075), .ZN(n1137) );
NAND4_X1 U840 ( .A1(n1149), .A2(n1150), .A3(n1098), .A4(n1151), .ZN(n1075) );
AND4_X1 U841 ( .A1(n1152), .A2(n991), .A3(n1153), .A4(n1154), .ZN(n1151) );
NAND3_X1 U842 ( .A1(n1029), .A2(n1028), .A3(n1155), .ZN(n991) );
NAND3_X1 U843 ( .A1(n1155), .A2(n1028), .A3(n1156), .ZN(n1098) );
NOR3_X1 U844 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1134) );
AND2_X1 U845 ( .A1(n1160), .A2(KEYINPUT57), .ZN(n1159) );
NOR3_X1 U846 ( .A1(KEYINPUT57), .A2(n1161), .A3(n1162), .ZN(n1158) );
AND2_X1 U847 ( .A1(n1162), .A2(n1161), .ZN(n1157) );
XNOR2_X1 U848 ( .A(n1163), .B(KEYINPUT16), .ZN(n1161) );
OR2_X1 U849 ( .A1(KEYINPUT12), .A2(n1160), .ZN(n1162) );
XOR2_X1 U850 ( .A(n1164), .B(n1165), .Z(n1160) );
NAND2_X1 U851 ( .A1(KEYINPUT19), .A2(n1166), .ZN(n1164) );
NOR2_X1 U852 ( .A1(n1032), .A2(G952), .ZN(n1083) );
XOR2_X1 U853 ( .A(n1167), .B(n1139), .Z(G48) );
NAND3_X1 U854 ( .A1(n1156), .A2(n1019), .A3(n1168), .ZN(n1139) );
XOR2_X1 U855 ( .A(n1169), .B(n1140), .Z(G45) );
NAND4_X1 U856 ( .A1(n1170), .A2(n1019), .A3(n1171), .A4(n1172), .ZN(n1140) );
XOR2_X1 U857 ( .A(G140), .B(n1173), .Z(G42) );
NOR2_X1 U858 ( .A1(KEYINPUT14), .A2(n1148), .ZN(n1173) );
NAND3_X1 U859 ( .A1(n1174), .A2(n1011), .A3(n1030), .ZN(n1148) );
NAND2_X1 U860 ( .A1(n1175), .A2(n1176), .ZN(G39) );
OR2_X1 U861 ( .A1(n1147), .A2(G137), .ZN(n1176) );
XOR2_X1 U862 ( .A(n1177), .B(KEYINPUT17), .Z(n1175) );
NAND2_X1 U863 ( .A1(G137), .A2(n1147), .ZN(n1177) );
NAND3_X1 U864 ( .A1(n1168), .A2(n1178), .A3(n1030), .ZN(n1147) );
XOR2_X1 U865 ( .A(G134), .B(n1179), .Z(G36) );
NOR2_X1 U866 ( .A1(n1146), .A2(n1180), .ZN(n1179) );
XOR2_X1 U867 ( .A(KEYINPUT61), .B(KEYINPUT49), .Z(n1180) );
NAND3_X1 U868 ( .A1(n1170), .A2(n1029), .A3(n1030), .ZN(n1146) );
XNOR2_X1 U869 ( .A(G131), .B(n1145), .ZN(G33) );
NAND3_X1 U870 ( .A1(n1170), .A2(n1156), .A3(n1030), .ZN(n1145) );
INV_X1 U871 ( .A(n1010), .ZN(n1030) );
NAND2_X1 U872 ( .A1(n1181), .A2(n1021), .ZN(n1010) );
AND3_X1 U873 ( .A1(n1011), .A2(n1182), .A3(n1025), .ZN(n1170) );
XNOR2_X1 U874 ( .A(G128), .B(n1144), .ZN(G30) );
NAND3_X1 U875 ( .A1(n1029), .A2(n1019), .A3(n1168), .ZN(n1144) );
AND4_X1 U876 ( .A1(n1011), .A2(n1046), .A3(n1027), .A4(n1182), .ZN(n1168) );
XOR2_X1 U877 ( .A(n1074), .B(n1183), .Z(G3) );
NOR2_X1 U878 ( .A1(KEYINPUT27), .A2(n1101), .ZN(n1183) );
AND3_X1 U879 ( .A1(n1178), .A2(n1155), .A3(n1025), .ZN(n1074) );
XOR2_X1 U880 ( .A(n1166), .B(n1143), .Z(G27) );
NAND3_X1 U881 ( .A1(n1174), .A2(n1019), .A3(n1023), .ZN(n1143) );
AND4_X1 U882 ( .A1(n1184), .A2(n1156), .A3(n1046), .A4(n1182), .ZN(n1174) );
NAND2_X1 U883 ( .A1(n998), .A2(n1185), .ZN(n1182) );
NAND4_X1 U884 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1068), .ZN(n1185) );
INV_X1 U885 ( .A(G900), .ZN(n1068) );
XNOR2_X1 U886 ( .A(G122), .B(n1149), .ZN(G24) );
NAND4_X1 U887 ( .A1(n1187), .A2(n1028), .A3(n1171), .A4(n1172), .ZN(n1149) );
INV_X1 U888 ( .A(n1006), .ZN(n1028) );
NAND2_X1 U889 ( .A1(n1184), .A2(n1026), .ZN(n1006) );
XOR2_X1 U890 ( .A(n1188), .B(n1189), .Z(G21) );
XNOR2_X1 U891 ( .A(G119), .B(KEYINPUT11), .ZN(n1189) );
NAND2_X1 U892 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
OR2_X1 U893 ( .A1(n1150), .A2(KEYINPUT63), .ZN(n1191) );
NAND3_X1 U894 ( .A1(n1187), .A2(n1027), .A3(n1192), .ZN(n1150) );
NAND4_X1 U895 ( .A1(n1192), .A2(n1023), .A3(n1193), .A4(KEYINPUT63), .ZN(n1190) );
NOR3_X1 U896 ( .A1(n1184), .A2(n1194), .A3(n1019), .ZN(n1193) );
INV_X1 U897 ( .A(n1195), .ZN(n1194) );
XOR2_X1 U898 ( .A(n1196), .B(G116), .Z(G18) );
NAND2_X1 U899 ( .A1(KEYINPUT51), .A2(n1152), .ZN(n1196) );
NAND3_X1 U900 ( .A1(n1025), .A2(n1029), .A3(n1187), .ZN(n1152) );
NOR2_X1 U901 ( .A1(n1171), .A2(n1197), .ZN(n1029) );
XOR2_X1 U902 ( .A(n1154), .B(n1198), .Z(G15) );
NAND2_X1 U903 ( .A1(KEYINPUT25), .A2(G113), .ZN(n1198) );
NAND3_X1 U904 ( .A1(n1025), .A2(n1156), .A3(n1187), .ZN(n1154) );
AND3_X1 U905 ( .A1(n1019), .A2(n1195), .A3(n1023), .ZN(n1187) );
NOR2_X1 U906 ( .A1(n1199), .A2(n1015), .ZN(n1023) );
XNOR2_X1 U907 ( .A(n1014), .B(KEYINPUT55), .ZN(n1199) );
INV_X1 U908 ( .A(n1036), .ZN(n1156) );
NAND2_X1 U909 ( .A1(n1197), .A2(n1171), .ZN(n1036) );
NOR2_X1 U910 ( .A1(n1046), .A2(n1184), .ZN(n1025) );
INV_X1 U911 ( .A(n1026), .ZN(n1046) );
XOR2_X1 U912 ( .A(G110), .B(n1200), .Z(G12) );
NOR2_X1 U913 ( .A1(KEYINPUT43), .A2(n1153), .ZN(n1200) );
NAND3_X1 U914 ( .A1(n1184), .A2(n1155), .A3(n1192), .ZN(n1153) );
NOR2_X1 U915 ( .A1(n1002), .A2(n1026), .ZN(n1192) );
XNOR2_X1 U916 ( .A(n1201), .B(n1087), .ZN(n1026) );
NAND2_X1 U917 ( .A1(G217), .A2(n1202), .ZN(n1087) );
NAND2_X1 U918 ( .A1(n1085), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U919 ( .A(n1204), .B(n1205), .ZN(n1085) );
XOR2_X1 U920 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U921 ( .A(n1208), .B(n1122), .Z(n1207) );
NAND2_X1 U922 ( .A1(n1209), .A2(n1210), .ZN(n1122) );
NAND2_X1 U923 ( .A1(G140), .A2(n1211), .ZN(n1210) );
NAND2_X1 U924 ( .A1(n1212), .A2(G221), .ZN(n1208) );
NOR2_X1 U925 ( .A1(G125), .A2(KEYINPUT2), .ZN(n1206) );
XOR2_X1 U926 ( .A(n1213), .B(n1214), .Z(n1204) );
XOR2_X1 U927 ( .A(KEYINPUT4), .B(G146), .Z(n1214) );
XOR2_X1 U928 ( .A(n1215), .B(G137), .Z(n1213) );
NAND2_X1 U929 ( .A1(n1216), .A2(KEYINPUT46), .ZN(n1215) );
XNOR2_X1 U930 ( .A(G119), .B(G128), .ZN(n1216) );
INV_X1 U931 ( .A(n1178), .ZN(n1002) );
NOR2_X1 U932 ( .A1(n1172), .A2(n1171), .ZN(n1178) );
XNOR2_X1 U933 ( .A(n1217), .B(G475), .ZN(n1171) );
OR2_X1 U934 ( .A1(n1096), .A2(G902), .ZN(n1217) );
XNOR2_X1 U935 ( .A(n1218), .B(n1219), .ZN(n1096) );
XOR2_X1 U936 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U937 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U938 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U939 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U940 ( .A(n1228), .ZN(n1227) );
INV_X1 U941 ( .A(n1229), .ZN(n1224) );
NAND2_X1 U942 ( .A1(n1230), .A2(n1229), .ZN(n1222) );
XOR2_X1 U943 ( .A(n1231), .B(n1232), .Z(n1229) );
AND2_X1 U944 ( .A1(G214), .A2(n1233), .ZN(n1232) );
XOR2_X1 U945 ( .A(G146), .B(G143), .Z(n1230) );
NAND2_X1 U946 ( .A1(KEYINPUT50), .A2(n1234), .ZN(n1220) );
XOR2_X1 U947 ( .A(G140), .B(G125), .Z(n1234) );
XOR2_X1 U948 ( .A(n1235), .B(n1236), .Z(n1218) );
XOR2_X1 U949 ( .A(KEYINPUT6), .B(G131), .Z(n1236) );
INV_X1 U950 ( .A(n1197), .ZN(n1172) );
XOR2_X1 U951 ( .A(n1237), .B(G478), .Z(n1197) );
OR2_X1 U952 ( .A1(n1091), .A2(G902), .ZN(n1237) );
XNOR2_X1 U953 ( .A(n1238), .B(n1239), .ZN(n1091) );
XOR2_X1 U954 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U955 ( .A(G116), .B(n1169), .Z(n1241) );
NAND2_X1 U956 ( .A1(G217), .A2(n1212), .ZN(n1240) );
AND2_X1 U957 ( .A1(G234), .A2(n1032), .ZN(n1212) );
XNOR2_X1 U958 ( .A(n1242), .B(n1243), .ZN(n1238) );
XNOR2_X1 U959 ( .A(n1244), .B(n1245), .ZN(n1243) );
NOR2_X1 U960 ( .A1(G107), .A2(KEYINPUT59), .ZN(n1244) );
AND3_X1 U961 ( .A1(n1019), .A2(n1195), .A3(n1011), .ZN(n1155) );
AND2_X1 U962 ( .A1(n1015), .A2(n1014), .ZN(n1011) );
NAND2_X1 U963 ( .A1(G221), .A2(n1202), .ZN(n1014) );
NAND2_X1 U964 ( .A1(G234), .A2(n1246), .ZN(n1202) );
XNOR2_X1 U965 ( .A(n1118), .B(n1247), .ZN(n1015) );
NOR2_X1 U966 ( .A1(G902), .A2(n1248), .ZN(n1247) );
NOR2_X1 U967 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U968 ( .A(n1251), .B(KEYINPUT41), .Z(n1250) );
NAND2_X1 U969 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U970 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U971 ( .A(n1256), .ZN(n1252) );
AND3_X1 U972 ( .A1(n1256), .A2(n1255), .A3(n1254), .ZN(n1249) );
NAND2_X1 U973 ( .A1(n1257), .A2(n1258), .ZN(n1254) );
NAND2_X1 U974 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND2_X1 U975 ( .A1(n1261), .A2(KEYINPUT20), .ZN(n1259) );
XOR2_X1 U976 ( .A(n1262), .B(n1061), .Z(n1261) );
XOR2_X1 U977 ( .A(n1263), .B(n1264), .Z(n1257) );
NAND2_X1 U978 ( .A1(n1265), .A2(n1266), .ZN(n1255) );
NAND2_X1 U979 ( .A1(KEYINPUT20), .A2(n1267), .ZN(n1266) );
NAND2_X1 U980 ( .A1(n1268), .A2(n1260), .ZN(n1267) );
INV_X1 U981 ( .A(KEYINPUT40), .ZN(n1260) );
XOR2_X1 U982 ( .A(n1264), .B(n1128), .Z(n1268) );
INV_X1 U983 ( .A(n1263), .ZN(n1128) );
XOR2_X1 U984 ( .A(n1269), .B(n1270), .Z(n1263) );
XOR2_X1 U985 ( .A(KEYINPUT9), .B(G101), .Z(n1270) );
NAND2_X1 U986 ( .A1(KEYINPUT53), .A2(n1271), .ZN(n1269) );
XOR2_X1 U987 ( .A(G107), .B(G104), .Z(n1271) );
NOR2_X1 U988 ( .A1(KEYINPUT26), .A2(n1058), .ZN(n1264) );
XOR2_X1 U989 ( .A(n1129), .B(G128), .Z(n1058) );
NAND3_X1 U990 ( .A1(n1272), .A2(n1273), .A3(n1226), .ZN(n1129) );
OR2_X1 U991 ( .A1(n1169), .A2(KEYINPUT47), .ZN(n1273) );
INV_X1 U992 ( .A(G143), .ZN(n1169) );
NAND2_X1 U993 ( .A1(n1228), .A2(KEYINPUT47), .ZN(n1272) );
XOR2_X1 U994 ( .A(G134), .B(n1061), .Z(n1265) );
XOR2_X1 U995 ( .A(n1274), .B(n1125), .Z(n1256) );
NOR2_X1 U996 ( .A1(n1067), .A2(G953), .ZN(n1125) );
INV_X1 U997 ( .A(G227), .ZN(n1067) );
NAND2_X1 U998 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U999 ( .A1(n1277), .A2(n1211), .ZN(n1276) );
INV_X1 U1000 ( .A(G110), .ZN(n1211) );
NAND2_X1 U1001 ( .A1(KEYINPUT3), .A2(n1064), .ZN(n1277) );
NAND2_X1 U1002 ( .A1(n1121), .A2(KEYINPUT3), .ZN(n1275) );
INV_X1 U1003 ( .A(n1209), .ZN(n1121) );
NAND2_X1 U1004 ( .A1(G110), .A2(n1064), .ZN(n1209) );
INV_X1 U1005 ( .A(G140), .ZN(n1064) );
INV_X1 U1006 ( .A(G469), .ZN(n1118) );
NAND2_X1 U1007 ( .A1(n998), .A2(n1278), .ZN(n1195) );
NAND4_X1 U1008 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1186), .ZN(n1278) );
XNOR2_X1 U1009 ( .A(KEYINPUT22), .B(n1078), .ZN(n1279) );
XNOR2_X1 U1010 ( .A(G898), .B(KEYINPUT0), .ZN(n1078) );
NAND3_X1 U1011 ( .A1(n1186), .A2(n1032), .A3(G952), .ZN(n998) );
NAND2_X1 U1012 ( .A1(G237), .A2(n1280), .ZN(n1186) );
XOR2_X1 U1013 ( .A(KEYINPUT54), .B(G234), .Z(n1280) );
AND2_X1 U1014 ( .A1(n1281), .A2(n1021), .ZN(n1019) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1282), .ZN(n1021) );
XOR2_X1 U1016 ( .A(KEYINPUT32), .B(n1181), .Z(n1281) );
INV_X1 U1017 ( .A(n1020), .ZN(n1181) );
NAND2_X1 U1018 ( .A1(n1283), .A2(n1042), .ZN(n1020) );
NAND2_X1 U1019 ( .A1(n1284), .A2(n1285), .ZN(n1042) );
XNOR2_X1 U1020 ( .A(KEYINPUT42), .B(n1041), .ZN(n1283) );
OR2_X1 U1021 ( .A1(n1285), .A2(n1284), .ZN(n1041) );
INV_X1 U1022 ( .A(n1136), .ZN(n1284) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1282), .ZN(n1136) );
NAND2_X1 U1024 ( .A1(n1246), .A2(n1286), .ZN(n1282) );
INV_X1 U1025 ( .A(G237), .ZN(n1286) );
XOR2_X1 U1026 ( .A(G902), .B(KEYINPUT52), .Z(n1246) );
NAND2_X1 U1027 ( .A1(n1287), .A2(n1203), .ZN(n1285) );
XOR2_X1 U1028 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1029 ( .A(n1166), .B(n1163), .Z(n1289) );
NAND2_X1 U1030 ( .A1(G224), .A2(n1032), .ZN(n1163) );
INV_X1 U1031 ( .A(G953), .ZN(n1032) );
INV_X1 U1032 ( .A(G125), .ZN(n1166) );
XNOR2_X1 U1033 ( .A(n1132), .B(n1165), .ZN(n1288) );
XNOR2_X1 U1034 ( .A(n1290), .B(G128), .ZN(n1165) );
XOR2_X1 U1035 ( .A(n1080), .B(n1291), .Z(n1132) );
NOR2_X1 U1036 ( .A1(KEYINPUT29), .A2(n1081), .ZN(n1291) );
XOR2_X1 U1037 ( .A(n1292), .B(n1293), .Z(n1081) );
NOR2_X1 U1038 ( .A1(KEYINPUT13), .A2(n1235), .ZN(n1293) );
XNOR2_X1 U1039 ( .A(G116), .B(n1294), .ZN(n1292) );
NOR2_X1 U1040 ( .A1(G119), .A2(KEYINPUT5), .ZN(n1294) );
XNOR2_X1 U1041 ( .A(n1295), .B(n1296), .ZN(n1080) );
XOR2_X1 U1042 ( .A(G110), .B(G107), .Z(n1296) );
XOR2_X1 U1043 ( .A(n1231), .B(G101), .Z(n1295) );
XNOR2_X1 U1044 ( .A(G104), .B(n1242), .ZN(n1231) );
XOR2_X1 U1045 ( .A(G122), .B(KEYINPUT44), .Z(n1242) );
INV_X1 U1046 ( .A(n1027), .ZN(n1184) );
XOR2_X1 U1047 ( .A(n1047), .B(G472), .Z(n1027) );
AND2_X1 U1048 ( .A1(n1297), .A2(n1203), .ZN(n1047) );
INV_X1 U1049 ( .A(G902), .ZN(n1203) );
NAND2_X1 U1050 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND3_X1 U1051 ( .A1(n1109), .A2(n1300), .A3(n1301), .ZN(n1299) );
XOR2_X1 U1052 ( .A(n1302), .B(n1303), .Z(n1301) );
NAND2_X1 U1053 ( .A1(KEYINPUT23), .A2(n1304), .ZN(n1302) );
INV_X1 U1054 ( .A(n1110), .ZN(n1304) );
NAND2_X1 U1055 ( .A1(n1305), .A2(n1306), .ZN(n1298) );
NAND2_X1 U1056 ( .A1(n1109), .A2(n1300), .ZN(n1306) );
INV_X1 U1057 ( .A(KEYINPUT10), .ZN(n1300) );
XOR2_X1 U1058 ( .A(n1290), .B(n1130), .Z(n1109) );
XNOR2_X1 U1059 ( .A(n1245), .B(n1061), .ZN(n1130) );
XOR2_X1 U1060 ( .A(G131), .B(G137), .Z(n1061) );
XOR2_X1 U1061 ( .A(G128), .B(n1262), .Z(n1245) );
INV_X1 U1062 ( .A(G134), .ZN(n1262) );
NAND4_X1 U1063 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1290) );
OR3_X1 U1064 ( .A1(n1167), .A2(G143), .A3(KEYINPUT45), .ZN(n1310) );
NAND2_X1 U1065 ( .A1(KEYINPUT45), .A2(n1228), .ZN(n1309) );
NOR2_X1 U1066 ( .A1(G143), .A2(G146), .ZN(n1228) );
OR2_X1 U1067 ( .A1(n1226), .A2(KEYINPUT62), .ZN(n1308) );
NAND2_X1 U1068 ( .A1(G146), .A2(G143), .ZN(n1226) );
NAND3_X1 U1069 ( .A1(G143), .A2(n1167), .A3(KEYINPUT62), .ZN(n1307) );
INV_X1 U1070 ( .A(G146), .ZN(n1167) );
XOR2_X1 U1071 ( .A(n1311), .B(n1303), .Z(n1305) );
XNOR2_X1 U1072 ( .A(n1312), .B(n1313), .ZN(n1303) );
XNOR2_X1 U1073 ( .A(KEYINPUT56), .B(n1105), .ZN(n1313) );
NAND2_X1 U1074 ( .A1(n1233), .A2(G210), .ZN(n1105) );
NOR2_X1 U1075 ( .A1(G953), .A2(G237), .ZN(n1233) );
NAND2_X1 U1076 ( .A1(KEYINPUT58), .A2(n1101), .ZN(n1312) );
INV_X1 U1077 ( .A(G101), .ZN(n1101) );
NAND2_X1 U1078 ( .A1(n1110), .A2(KEYINPUT23), .ZN(n1311) );
XOR2_X1 U1079 ( .A(n1235), .B(n1314), .Z(n1110) );
NOR2_X1 U1080 ( .A1(KEYINPUT31), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U1081 ( .A(G116), .B(G119), .ZN(n1315) );
INV_X1 U1082 ( .A(G113), .ZN(n1235) );
endmodule


