//Key = 0111111101111001101110011110101001111001101101100010100101110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333;

XNOR2_X1 U716 ( .A(G107), .B(n1003), .ZN(G9) );
NOR2_X1 U717 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR3_X1 U718 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
NOR2_X1 U719 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NAND3_X1 U720 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1006) );
NAND3_X1 U721 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND2_X1 U722 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NAND2_X1 U723 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U724 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U725 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
OR2_X1 U726 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U727 ( .A1(n1027), .A2(n1028), .ZN(n1021) );
NAND3_X1 U728 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND2_X1 U729 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U730 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1030) );
NAND2_X1 U731 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
OR2_X1 U732 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U733 ( .A1(n1041), .A2(n1042), .ZN(n1029) );
XOR2_X1 U734 ( .A(KEYINPUT54), .B(n1033), .Z(n1042) );
NAND2_X1 U735 ( .A1(n1043), .A2(n1044), .ZN(n1014) );
XNOR2_X1 U736 ( .A(KEYINPUT61), .B(n1010), .ZN(n1043) );
NAND3_X1 U737 ( .A1(n1023), .A2(n1027), .A3(n1019), .ZN(n1010) );
INV_X1 U738 ( .A(n1045), .ZN(n1019) );
NOR3_X1 U739 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1004) );
INV_X1 U740 ( .A(n1011), .ZN(n1046) );
NAND4_X1 U741 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1011) );
NOR3_X1 U742 ( .A1(n1051), .A2(n1044), .A3(n1052), .ZN(n1050) );
NOR2_X1 U743 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U744 ( .A1(n1055), .A2(n1056), .A3(n1039), .ZN(n1051) );
NOR3_X1 U745 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1049) );
NOR2_X1 U746 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
XNOR2_X1 U747 ( .A(n1062), .B(n1063), .ZN(n1057) );
XNOR2_X1 U748 ( .A(n1064), .B(n1065), .ZN(n1048) );
NAND2_X1 U749 ( .A1(KEYINPUT10), .A2(G472), .ZN(n1064) );
XNOR2_X1 U750 ( .A(G475), .B(n1066), .ZN(n1047) );
XOR2_X1 U751 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U752 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U753 ( .A1(G953), .A2(n1071), .ZN(n1070) );
NAND2_X1 U754 ( .A1(G900), .A2(G227), .ZN(n1071) );
NAND2_X1 U755 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
NAND2_X1 U756 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XOR2_X1 U757 ( .A(n1075), .B(n1076), .Z(n1072) );
XNOR2_X1 U758 ( .A(n1077), .B(KEYINPUT58), .ZN(n1076) );
NAND2_X1 U759 ( .A1(KEYINPUT59), .A2(n1078), .ZN(n1077) );
XOR2_X1 U760 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U761 ( .A(n1081), .B(n1082), .ZN(n1080) );
INV_X1 U762 ( .A(G131), .ZN(n1082) );
NAND3_X1 U763 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
NAND2_X1 U764 ( .A1(G137), .A2(n1086), .ZN(n1085) );
OR3_X1 U765 ( .A1(n1086), .A2(G137), .A3(n1087), .ZN(n1084) );
INV_X1 U766 ( .A(KEYINPUT28), .ZN(n1086) );
NAND2_X1 U767 ( .A1(n1087), .A2(n1088), .ZN(n1083) );
NAND2_X1 U768 ( .A1(n1089), .A2(KEYINPUT28), .ZN(n1088) );
XNOR2_X1 U769 ( .A(G137), .B(KEYINPUT29), .ZN(n1089) );
NAND2_X1 U770 ( .A1(KEYINPUT5), .A2(n1090), .ZN(n1079) );
AND2_X1 U771 ( .A1(n1091), .A2(n1012), .ZN(n1067) );
XOR2_X1 U772 ( .A(n1092), .B(n1093), .Z(G69) );
NOR2_X1 U773 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U774 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U775 ( .A1(KEYINPUT16), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U776 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND3_X1 U777 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1092) );
NAND2_X1 U778 ( .A1(KEYINPUT12), .A2(n1094), .ZN(n1103) );
NAND2_X1 U779 ( .A1(G953), .A2(n1104), .ZN(n1102) );
NAND2_X1 U780 ( .A1(G224), .A2(n1105), .ZN(n1104) );
NAND2_X1 U781 ( .A1(G898), .A2(n1106), .ZN(n1105) );
INV_X1 U782 ( .A(KEYINPUT12), .ZN(n1106) );
NAND3_X1 U783 ( .A1(KEYINPUT40), .A2(n1107), .A3(n1012), .ZN(n1101) );
NOR2_X1 U784 ( .A1(n1108), .A2(n1109), .ZN(G66) );
NOR3_X1 U785 ( .A1(n1063), .A2(n1110), .A3(n1111), .ZN(n1109) );
NOR3_X1 U786 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
INV_X1 U787 ( .A(n1115), .ZN(n1112) );
NOR2_X1 U788 ( .A1(n1116), .A2(n1115), .ZN(n1110) );
NOR2_X1 U789 ( .A1(n1117), .A2(n1113), .ZN(n1116) );
XOR2_X1 U790 ( .A(G217), .B(KEYINPUT23), .Z(n1113) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1118), .ZN(G63) );
XNOR2_X1 U792 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1121), .ZN(n1120) );
XOR2_X1 U794 ( .A(KEYINPUT30), .B(G478), .Z(n1121) );
NOR3_X1 U795 ( .A1(n1122), .A2(n1108), .A3(n1123), .ZN(G60) );
NOR3_X1 U796 ( .A1(n1114), .A2(n1124), .A3(n1125), .ZN(n1123) );
NOR2_X1 U797 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
XOR2_X1 U798 ( .A(KEYINPUT24), .B(n1124), .Z(n1127) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1114), .ZN(n1126) );
INV_X1 U800 ( .A(G475), .ZN(n1125) );
XNOR2_X1 U801 ( .A(G104), .B(n1128), .ZN(G6) );
NOR2_X1 U802 ( .A1(n1108), .A2(n1129), .ZN(G57) );
XOR2_X1 U803 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U805 ( .A(KEYINPUT41), .B(n1134), .ZN(n1133) );
INV_X1 U806 ( .A(n1135), .ZN(n1132) );
NAND2_X1 U807 ( .A1(n1136), .A2(KEYINPUT34), .ZN(n1130) );
XOR2_X1 U808 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U809 ( .A1(n1139), .A2(n1114), .ZN(n1138) );
NOR2_X1 U810 ( .A1(n1108), .A2(n1140), .ZN(G54) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U812 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U813 ( .A1(n1145), .A2(KEYINPUT7), .ZN(n1143) );
XOR2_X1 U814 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U815 ( .A(n1148), .B(n1149), .ZN(n1146) );
XNOR2_X1 U816 ( .A(n1150), .B(n1151), .ZN(n1141) );
NAND3_X1 U817 ( .A1(G469), .A2(n1152), .A3(G902), .ZN(n1150) );
XNOR2_X1 U818 ( .A(KEYINPUT26), .B(n1008), .ZN(n1152) );
NOR2_X1 U819 ( .A1(n1108), .A2(n1153), .ZN(G51) );
XOR2_X1 U820 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U821 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR3_X1 U822 ( .A1(n1114), .A2(KEYINPUT37), .A3(n1158), .ZN(n1157) );
INV_X1 U823 ( .A(G210), .ZN(n1158) );
NAND2_X1 U824 ( .A1(G902), .A2(n1008), .ZN(n1114) );
INV_X1 U825 ( .A(n1117), .ZN(n1008) );
NOR2_X1 U826 ( .A1(n1107), .A2(n1091), .ZN(n1117) );
NAND4_X1 U827 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1091) );
NOR4_X1 U828 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
INV_X1 U829 ( .A(n1167), .ZN(n1166) );
NAND2_X1 U830 ( .A1(n1168), .A2(n1169), .ZN(n1161) );
NAND2_X1 U831 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U832 ( .A1(n1172), .A2(n1032), .ZN(n1171) );
XNOR2_X1 U833 ( .A(n1025), .B(KEYINPUT18), .ZN(n1172) );
NAND2_X1 U834 ( .A1(n1173), .A2(n1041), .ZN(n1170) );
XNOR2_X1 U835 ( .A(n1025), .B(KEYINPUT33), .ZN(n1173) );
NAND4_X1 U836 ( .A1(n1128), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1107) );
AND3_X1 U837 ( .A1(n1003), .A2(n1177), .A3(n1178), .ZN(n1176) );
NAND2_X1 U838 ( .A1(n1026), .A2(n1179), .ZN(n1003) );
NAND2_X1 U839 ( .A1(n1180), .A2(n1181), .ZN(n1175) );
NAND2_X1 U840 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U841 ( .A1(n1032), .A2(n1184), .ZN(n1183) );
NAND2_X1 U842 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U843 ( .A1(n1027), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U844 ( .A(KEYINPUT38), .B(n1037), .ZN(n1187) );
NAND2_X1 U845 ( .A1(n1025), .A2(n1033), .ZN(n1185) );
NAND2_X1 U846 ( .A1(n1025), .A2(n1179), .ZN(n1128) );
AND4_X1 U847 ( .A1(n1188), .A2(n1180), .A3(n1036), .A4(n1034), .ZN(n1179) );
NOR2_X1 U848 ( .A1(n1012), .A2(G952), .ZN(n1108) );
XNOR2_X1 U849 ( .A(n1189), .B(n1159), .ZN(G48) );
NAND2_X1 U850 ( .A1(n1190), .A2(n1025), .ZN(n1159) );
NAND2_X1 U851 ( .A1(KEYINPUT20), .A2(n1191), .ZN(n1189) );
XNOR2_X1 U852 ( .A(G143), .B(n1160), .ZN(G45) );
NAND3_X1 U853 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1160) );
NOR3_X1 U854 ( .A1(n1195), .A2(n1196), .A3(n1037), .ZN(n1194) );
XNOR2_X1 U855 ( .A(G140), .B(n1197), .ZN(G42) );
NAND2_X1 U856 ( .A1(n1198), .A2(n1041), .ZN(n1197) );
NAND2_X1 U857 ( .A1(n1199), .A2(n1200), .ZN(G39) );
NAND2_X1 U858 ( .A1(G137), .A2(n1167), .ZN(n1200) );
XOR2_X1 U859 ( .A(KEYINPUT3), .B(n1201), .Z(n1199) );
NOR2_X1 U860 ( .A1(G137), .A2(n1167), .ZN(n1201) );
NAND4_X1 U861 ( .A1(n1168), .A2(n1027), .A3(n1202), .A4(n1203), .ZN(n1167) );
XNOR2_X1 U862 ( .A(n1204), .B(n1165), .ZN(G36) );
AND3_X1 U863 ( .A1(n1032), .A2(n1026), .A3(n1168), .ZN(n1165) );
XNOR2_X1 U864 ( .A(G131), .B(n1205), .ZN(G33) );
NAND2_X1 U865 ( .A1(n1198), .A2(n1032), .ZN(n1205) );
AND2_X1 U866 ( .A1(n1168), .A2(n1025), .ZN(n1198) );
AND4_X1 U867 ( .A1(n1016), .A2(n1188), .A3(n1206), .A4(n1018), .ZN(n1168) );
XOR2_X1 U868 ( .A(n1207), .B(n1164), .Z(G30) );
AND2_X1 U869 ( .A1(n1190), .A2(n1026), .ZN(n1164) );
AND4_X1 U870 ( .A1(n1202), .A2(n1193), .A3(n1188), .A4(n1203), .ZN(n1190) );
XNOR2_X1 U871 ( .A(G128), .B(KEYINPUT46), .ZN(n1207) );
XNOR2_X1 U872 ( .A(n1208), .B(n1209), .ZN(G3) );
NOR2_X1 U873 ( .A1(n1195), .A2(n1210), .ZN(n1209) );
INV_X1 U874 ( .A(n1032), .ZN(n1195) );
XOR2_X1 U875 ( .A(G125), .B(n1163), .Z(G27) );
AND4_X1 U876 ( .A1(n1193), .A2(n1025), .A3(n1041), .A4(n1033), .ZN(n1163) );
INV_X1 U877 ( .A(n1211), .ZN(n1025) );
AND2_X1 U878 ( .A1(n1212), .A2(n1206), .ZN(n1193) );
NAND2_X1 U879 ( .A1(n1045), .A2(n1213), .ZN(n1206) );
NAND4_X1 U880 ( .A1(G902), .A2(G953), .A3(n1214), .A4(n1074), .ZN(n1213) );
INV_X1 U881 ( .A(G900), .ZN(n1074) );
XOR2_X1 U882 ( .A(G122), .B(n1215), .Z(G24) );
NOR3_X1 U883 ( .A1(n1182), .A2(n1216), .A3(n1217), .ZN(n1215) );
NOR2_X1 U884 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U885 ( .A(KEYINPUT17), .ZN(n1219) );
NOR2_X1 U886 ( .A1(n1212), .A2(n1220), .ZN(n1218) );
NOR2_X1 U887 ( .A1(KEYINPUT17), .A2(n1180), .ZN(n1216) );
NAND3_X1 U888 ( .A1(n1192), .A2(n1221), .A3(n1023), .ZN(n1182) );
AND3_X1 U889 ( .A1(n1036), .A2(n1034), .A3(n1033), .ZN(n1023) );
XNOR2_X1 U890 ( .A(G119), .B(n1178), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1180), .A2(n1203), .A3(n1033), .A4(n1222), .ZN(n1178) );
AND2_X1 U892 ( .A1(n1027), .A2(n1202), .ZN(n1222) );
XNOR2_X1 U893 ( .A(G116), .B(n1223), .ZN(G18) );
NOR2_X1 U894 ( .A1(n1224), .A2(KEYINPUT44), .ZN(n1223) );
INV_X1 U895 ( .A(n1177), .ZN(n1224) );
NAND4_X1 U896 ( .A1(n1032), .A2(n1033), .A3(n1026), .A4(n1180), .ZN(n1177) );
NOR2_X1 U897 ( .A1(n1225), .A2(n1196), .ZN(n1026) );
XNOR2_X1 U898 ( .A(G113), .B(n1226), .ZN(G15) );
NAND4_X1 U899 ( .A1(n1032), .A2(n1033), .A3(n1180), .A4(n1227), .ZN(n1226) );
XNOR2_X1 U900 ( .A(KEYINPUT31), .B(n1211), .ZN(n1227) );
NAND2_X1 U901 ( .A1(n1192), .A2(n1196), .ZN(n1211) );
INV_X1 U902 ( .A(n1221), .ZN(n1196) );
XOR2_X1 U903 ( .A(n1225), .B(KEYINPUT60), .Z(n1192) );
NOR2_X1 U904 ( .A1(n1040), .A2(n1228), .ZN(n1033) );
INV_X1 U905 ( .A(n1039), .ZN(n1228) );
NOR2_X1 U906 ( .A1(n1202), .A2(n1036), .ZN(n1032) );
INV_X1 U907 ( .A(n1203), .ZN(n1036) );
INV_X1 U908 ( .A(n1034), .ZN(n1202) );
XNOR2_X1 U909 ( .A(G110), .B(n1174), .ZN(G12) );
NAND2_X1 U910 ( .A1(n1041), .A2(n1229), .ZN(n1174) );
INV_X1 U911 ( .A(n1210), .ZN(n1229) );
NAND3_X1 U912 ( .A1(n1188), .A2(n1180), .A3(n1027), .ZN(n1210) );
NOR2_X1 U913 ( .A1(n1221), .A2(n1225), .ZN(n1027) );
XNOR2_X1 U914 ( .A(n1066), .B(n1230), .ZN(n1225) );
NOR2_X1 U915 ( .A1(G475), .A2(KEYINPUT62), .ZN(n1230) );
NOR2_X1 U916 ( .A1(G902), .A2(n1124), .ZN(n1066) );
AND2_X1 U917 ( .A1(n1231), .A2(n1232), .ZN(n1124) );
NAND2_X1 U918 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U919 ( .A(KEYINPUT4), .B(n1235), .Z(n1231) );
NOR2_X1 U920 ( .A1(n1234), .A2(n1233), .ZN(n1235) );
XOR2_X1 U921 ( .A(n1236), .B(n1237), .Z(n1233) );
XNOR2_X1 U922 ( .A(n1238), .B(n1239), .ZN(n1237) );
XNOR2_X1 U923 ( .A(n1191), .B(G131), .ZN(n1239) );
NAND3_X1 U924 ( .A1(n1240), .A2(n1241), .A3(G214), .ZN(n1238) );
XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n1012), .ZN(n1240) );
XOR2_X1 U926 ( .A(n1242), .B(n1243), .Z(n1236) );
NAND2_X1 U927 ( .A1(KEYINPUT50), .A2(G143), .ZN(n1242) );
XNOR2_X1 U928 ( .A(G104), .B(n1244), .ZN(n1234) );
XNOR2_X1 U929 ( .A(G122), .B(n1245), .ZN(n1244) );
NAND2_X1 U930 ( .A1(n1246), .A2(n1055), .ZN(n1221) );
NAND2_X1 U931 ( .A1(n1053), .A2(n1054), .ZN(n1055) );
NAND2_X1 U932 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
INV_X1 U933 ( .A(n1053), .ZN(n1248) );
NOR2_X1 U934 ( .A1(n1249), .A2(G902), .ZN(n1053) );
INV_X1 U935 ( .A(n1119), .ZN(n1249) );
XNOR2_X1 U936 ( .A(n1250), .B(n1251), .ZN(n1119) );
XNOR2_X1 U937 ( .A(n1252), .B(n1253), .ZN(n1251) );
XOR2_X1 U938 ( .A(n1254), .B(n1255), .Z(n1250) );
NOR2_X1 U939 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U940 ( .A(n1258), .B(KEYINPUT43), .Z(n1257) );
NAND2_X1 U941 ( .A1(n1259), .A2(n1204), .ZN(n1258) );
NOR2_X1 U942 ( .A1(n1204), .A2(n1259), .ZN(n1256) );
XOR2_X1 U943 ( .A(G143), .B(n1260), .Z(n1259) );
INV_X1 U944 ( .A(G134), .ZN(n1204) );
NAND2_X1 U945 ( .A1(G217), .A2(n1261), .ZN(n1254) );
XNOR2_X1 U946 ( .A(n1054), .B(KEYINPUT27), .ZN(n1247) );
XOR2_X1 U947 ( .A(G478), .B(KEYINPUT15), .Z(n1054) );
NOR2_X1 U948 ( .A1(n1009), .A2(n1220), .ZN(n1180) );
AND2_X1 U949 ( .A1(n1045), .A2(n1262), .ZN(n1220) );
NAND3_X1 U950 ( .A1(n1094), .A2(n1214), .A3(G902), .ZN(n1262) );
NOR2_X1 U951 ( .A1(n1012), .A2(G898), .ZN(n1094) );
NAND3_X1 U952 ( .A1(n1214), .A2(n1012), .A3(G952), .ZN(n1045) );
NAND2_X1 U953 ( .A1(G237), .A2(G234), .ZN(n1214) );
INV_X1 U954 ( .A(n1212), .ZN(n1009) );
NOR2_X1 U955 ( .A1(n1016), .A2(n1044), .ZN(n1212) );
INV_X1 U956 ( .A(n1018), .ZN(n1044) );
NAND2_X1 U957 ( .A1(G214), .A2(n1263), .ZN(n1018) );
INV_X1 U958 ( .A(n1059), .ZN(n1016) );
XNOR2_X1 U959 ( .A(n1264), .B(n1265), .ZN(n1059) );
AND2_X1 U960 ( .A1(n1263), .A2(G210), .ZN(n1265) );
NAND2_X1 U961 ( .A1(n1266), .A2(n1241), .ZN(n1263) );
NAND3_X1 U962 ( .A1(n1267), .A2(n1268), .A3(n1266), .ZN(n1264) );
NAND2_X1 U963 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
INV_X1 U964 ( .A(n1271), .ZN(n1270) );
NAND2_X1 U965 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
NAND2_X1 U966 ( .A1(KEYINPUT45), .A2(n1274), .ZN(n1273) );
NAND2_X1 U967 ( .A1(n1154), .A2(n1275), .ZN(n1274) );
NAND2_X1 U968 ( .A1(n1154), .A2(n1276), .ZN(n1272) );
INV_X1 U969 ( .A(KEYINPUT45), .ZN(n1276) );
NAND3_X1 U970 ( .A1(n1154), .A2(n1275), .A3(n1271), .ZN(n1267) );
XNOR2_X1 U971 ( .A(n1156), .B(KEYINPUT51), .ZN(n1271) );
XNOR2_X1 U972 ( .A(n1277), .B(n1090), .ZN(n1156) );
XNOR2_X1 U973 ( .A(G125), .B(n1278), .ZN(n1277) );
AND2_X1 U974 ( .A1(n1012), .A2(G224), .ZN(n1278) );
INV_X1 U975 ( .A(KEYINPUT32), .ZN(n1275) );
XOR2_X1 U976 ( .A(n1279), .B(n1097), .Z(n1154) );
XNOR2_X1 U977 ( .A(n1252), .B(n1280), .ZN(n1097) );
XOR2_X1 U978 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U979 ( .A1(KEYINPUT13), .A2(n1245), .ZN(n1281) );
XNOR2_X1 U980 ( .A(G116), .B(G122), .ZN(n1252) );
NAND2_X1 U981 ( .A1(n1283), .A2(KEYINPUT6), .ZN(n1279) );
XOR2_X1 U982 ( .A(n1099), .B(n1100), .Z(n1283) );
NAND2_X1 U983 ( .A1(KEYINPUT11), .A2(G101), .ZN(n1099) );
INV_X1 U984 ( .A(n1037), .ZN(n1188) );
NAND2_X1 U985 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND2_X1 U986 ( .A1(n1284), .A2(n1056), .ZN(n1040) );
NAND2_X1 U987 ( .A1(n1060), .A2(n1061), .ZN(n1056) );
INV_X1 U988 ( .A(G469), .ZN(n1061) );
NAND2_X1 U989 ( .A1(n1285), .A2(G469), .ZN(n1284) );
XNOR2_X1 U990 ( .A(n1060), .B(KEYINPUT0), .ZN(n1285) );
AND2_X1 U991 ( .A1(n1286), .A2(n1266), .ZN(n1060) );
XOR2_X1 U992 ( .A(n1287), .B(n1288), .Z(n1286) );
NAND2_X1 U993 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U994 ( .A1(n1291), .A2(n1151), .ZN(n1290) );
INV_X1 U995 ( .A(G140), .ZN(n1151) );
XOR2_X1 U996 ( .A(KEYINPUT52), .B(n1144), .Z(n1291) );
NAND2_X1 U997 ( .A1(n1144), .A2(G140), .ZN(n1289) );
XOR2_X1 U998 ( .A(G110), .B(n1292), .Z(n1144) );
AND2_X1 U999 ( .A1(n1012), .A2(G227), .ZN(n1292) );
NAND2_X1 U1000 ( .A1(n1293), .A2(n1294), .ZN(n1287) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U1002 ( .A(n1297), .B(n1090), .ZN(n1296) );
INV_X1 U1003 ( .A(n1298), .ZN(n1090) );
XNOR2_X1 U1004 ( .A(KEYINPUT47), .B(n1299), .ZN(n1295) );
XOR2_X1 U1005 ( .A(n1300), .B(KEYINPUT48), .Z(n1293) );
NAND2_X1 U1006 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XNOR2_X1 U1007 ( .A(n1297), .B(n1298), .ZN(n1302) );
NAND2_X1 U1008 ( .A1(KEYINPUT25), .A2(n1147), .ZN(n1297) );
XNOR2_X1 U1009 ( .A(n1208), .B(n1100), .ZN(n1147) );
XNOR2_X1 U1010 ( .A(n1303), .B(n1253), .ZN(n1100) );
XOR2_X1 U1011 ( .A(G107), .B(KEYINPUT49), .Z(n1253) );
XNOR2_X1 U1012 ( .A(G104), .B(KEYINPUT19), .ZN(n1303) );
XNOR2_X1 U1013 ( .A(n1149), .B(n1299), .ZN(n1301) );
INV_X1 U1014 ( .A(KEYINPUT47), .ZN(n1149) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1304), .ZN(n1039) );
NOR2_X1 U1016 ( .A1(n1034), .A2(n1203), .ZN(n1041) );
NAND3_X1 U1017 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1203) );
OR2_X1 U1018 ( .A1(n1139), .A2(KEYINPUT57), .ZN(n1307) );
NAND3_X1 U1019 ( .A1(KEYINPUT57), .A2(n1139), .A3(n1308), .ZN(n1306) );
INV_X1 U1020 ( .A(n1065), .ZN(n1308) );
NAND2_X1 U1021 ( .A1(n1309), .A2(n1065), .ZN(n1305) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1266), .ZN(n1065) );
XOR2_X1 U1023 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1024 ( .A1(KEYINPUT14), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1025 ( .A(n1137), .B(n1314), .Z(n1313) );
XOR2_X1 U1026 ( .A(KEYINPUT55), .B(KEYINPUT42), .Z(n1314) );
XOR2_X1 U1027 ( .A(n1315), .B(n1316), .Z(n1137) );
XOR2_X1 U1028 ( .A(G119), .B(G116), .Z(n1316) );
XNOR2_X1 U1029 ( .A(n1148), .B(n1245), .ZN(n1315) );
INV_X1 U1030 ( .A(G113), .ZN(n1245) );
XNOR2_X1 U1031 ( .A(n1298), .B(n1299), .ZN(n1148) );
XNOR2_X1 U1032 ( .A(n1317), .B(G131), .ZN(n1299) );
NAND2_X1 U1033 ( .A1(n1318), .A2(KEYINPUT2), .ZN(n1317) );
XNOR2_X1 U1034 ( .A(G137), .B(n1087), .ZN(n1318) );
XOR2_X1 U1035 ( .A(G134), .B(KEYINPUT9), .Z(n1087) );
XOR2_X1 U1036 ( .A(G143), .B(n1319), .Z(n1298) );
NAND2_X1 U1037 ( .A1(n1134), .A2(n1135), .ZN(n1311) );
NAND4_X1 U1038 ( .A1(G210), .A2(G101), .A3(n1241), .A4(n1012), .ZN(n1135) );
NAND2_X1 U1039 ( .A1(n1208), .A2(n1320), .ZN(n1134) );
NAND3_X1 U1040 ( .A1(n1241), .A2(n1012), .A3(G210), .ZN(n1320) );
INV_X1 U1041 ( .A(G237), .ZN(n1241) );
INV_X1 U1042 ( .A(G101), .ZN(n1208) );
NAND2_X1 U1043 ( .A1(KEYINPUT57), .A2(n1321), .ZN(n1309) );
XNOR2_X1 U1044 ( .A(KEYINPUT35), .B(n1139), .ZN(n1321) );
INV_X1 U1045 ( .A(G472), .ZN(n1139) );
XNOR2_X1 U1046 ( .A(n1062), .B(n1322), .ZN(n1034) );
NOR2_X1 U1047 ( .A1(KEYINPUT8), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n1324), .ZN(n1323) );
INV_X1 U1049 ( .A(n1063), .ZN(n1324) );
NOR2_X1 U1050 ( .A1(n1115), .A2(G902), .ZN(n1063) );
XNOR2_X1 U1051 ( .A(n1325), .B(n1326), .ZN(n1115) );
XOR2_X1 U1052 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1053 ( .A(n1329), .B(n1330), .ZN(n1328) );
INV_X1 U1054 ( .A(G137), .ZN(n1330) );
NAND2_X1 U1055 ( .A1(n1261), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1056 ( .A(KEYINPUT21), .B(G221), .Z(n1331) );
AND2_X1 U1057 ( .A1(G234), .A2(n1012), .ZN(n1261) );
INV_X1 U1058 ( .A(G953), .ZN(n1012) );
XNOR2_X1 U1059 ( .A(KEYINPUT56), .B(KEYINPUT1), .ZN(n1327) );
XOR2_X1 U1060 ( .A(n1332), .B(n1319), .Z(n1325) );
XNOR2_X1 U1061 ( .A(n1191), .B(n1260), .ZN(n1319) );
XOR2_X1 U1062 ( .A(G128), .B(KEYINPUT63), .Z(n1260) );
INV_X1 U1063 ( .A(G146), .ZN(n1191) );
XNOR2_X1 U1064 ( .A(n1282), .B(n1243), .ZN(n1332) );
XNOR2_X1 U1065 ( .A(n1075), .B(KEYINPUT36), .ZN(n1243) );
XNOR2_X1 U1066 ( .A(G125), .B(G140), .ZN(n1075) );
XOR2_X1 U1067 ( .A(G110), .B(G119), .Z(n1282) );
NAND2_X1 U1068 ( .A1(n1333), .A2(n1304), .ZN(n1062) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1266), .ZN(n1304) );
INV_X1 U1070 ( .A(G902), .ZN(n1266) );
XOR2_X1 U1071 ( .A(KEYINPUT22), .B(G217), .Z(n1333) );
endmodule


