//Key = 0001100110110000011010101101111100000110011010000111100000010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407;

XOR2_X1 U778 ( .A(n1075), .B(n1076), .Z(G9) );
NAND2_X1 U779 ( .A1(KEYINPUT4), .A2(G107), .ZN(n1076) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR3_X1 U781 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1078) );
NOR4_X1 U782 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1079), .ZN(n1077) );
AND4_X1 U783 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1079) );
NOR3_X1 U784 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
XOR2_X1 U785 ( .A(n1090), .B(KEYINPUT27), .Z(n1089) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1088) );
NOR2_X1 U787 ( .A1(n1093), .A2(KEYINPUT35), .ZN(n1092) );
NAND3_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1087) );
NOR3_X1 U789 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1085) );
AND3_X1 U790 ( .A1(KEYINPUT3), .A2(n1100), .A3(G475), .ZN(n1099) );
NOR2_X1 U791 ( .A1(KEYINPUT3), .A2(G475), .ZN(n1098) );
XNOR2_X1 U792 ( .A(KEYINPUT63), .B(n1101), .ZN(n1097) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1082) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR4_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
NOR3_X1 U796 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1107) );
AND2_X1 U797 ( .A1(n1113), .A2(KEYINPUT28), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1094), .ZN(n1111) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1106) );
NOR2_X1 U800 ( .A1(KEYINPUT28), .A2(n1117), .ZN(n1116) );
INV_X1 U801 ( .A(n1110), .ZN(n1115) );
NOR4_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1114), .A4(n1110), .ZN(n1104) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U804 ( .A1(n1122), .A2(n1109), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1123), .A2(n1108), .ZN(n1120) );
INV_X1 U806 ( .A(n1124), .ZN(n1108) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND3_X1 U809 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1080) );
NAND4_X1 U810 ( .A1(n1132), .A2(n1094), .A3(n1133), .A4(n1134), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1109), .A2(n1110), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NAND2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U814 ( .A(KEYINPUT32), .B(n1139), .Z(n1138) );
NAND2_X1 U815 ( .A1(n1124), .A2(n1140), .ZN(n1135) );
OR2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U817 ( .A(n1143), .ZN(n1129) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(G72) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1130), .ZN(n1145) );
AND2_X1 U820 ( .A1(G227), .A2(G900), .ZN(n1146) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1149), .A2(n1130), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1149) );
OR3_X1 U824 ( .A1(n1152), .A2(n1151), .A3(n1130), .ZN(n1147) );
XNOR2_X1 U825 ( .A(n1153), .B(n1154), .ZN(n1151) );
NOR2_X1 U826 ( .A1(KEYINPUT1), .A2(n1155), .ZN(n1154) );
XOR2_X1 U827 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U828 ( .A(G137), .B(G134), .Z(n1157) );
XOR2_X1 U829 ( .A(n1158), .B(G131), .Z(n1156) );
XOR2_X1 U830 ( .A(n1159), .B(n1160), .Z(G69) );
NOR2_X1 U831 ( .A1(n1161), .A2(n1130), .ZN(n1160) );
AND2_X1 U832 ( .A1(G224), .A2(G898), .ZN(n1161) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1130), .ZN(n1163) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND3_X1 U836 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1165) );
NOR3_X1 U837 ( .A1(n1170), .A2(n1143), .A3(n1171), .ZN(n1169) );
XOR2_X1 U838 ( .A(KEYINPUT36), .B(n1172), .Z(n1168) );
XNOR2_X1 U839 ( .A(KEYINPUT20), .B(n1173), .ZN(n1167) );
NAND3_X1 U840 ( .A1(G898), .A2(n1166), .A3(G953), .ZN(n1162) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1166) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1174) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(G66) );
XOR2_X1 U844 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U845 ( .A(n1182), .B(KEYINPUT22), .Z(n1180) );
NAND2_X1 U846 ( .A1(n1093), .A2(n1183), .ZN(n1182) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1184), .ZN(G63) );
XOR2_X1 U848 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U849 ( .A1(n1183), .A2(G478), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1187), .ZN(G60) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U852 ( .A1(n1183), .A2(G475), .ZN(n1188) );
XNOR2_X1 U853 ( .A(G104), .B(n1190), .ZN(G6) );
NOR2_X1 U854 ( .A1(n1178), .A2(n1191), .ZN(G57) );
XOR2_X1 U855 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U856 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U857 ( .A(n1196), .B(n1197), .Z(n1192) );
XOR2_X1 U858 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U859 ( .A1(G101), .A2(KEYINPUT61), .ZN(n1199) );
NAND2_X1 U860 ( .A1(n1183), .A2(G472), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1178), .A2(n1200), .ZN(G54) );
XOR2_X1 U862 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U863 ( .A(n1203), .B(n1204), .ZN(n1202) );
XOR2_X1 U864 ( .A(n1205), .B(n1206), .Z(n1201) );
NAND2_X1 U865 ( .A1(n1183), .A2(G469), .ZN(n1206) );
NAND3_X1 U866 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1205) );
NAND2_X1 U867 ( .A1(KEYINPUT54), .A2(n1210), .ZN(n1209) );
OR3_X1 U868 ( .A1(n1210), .A2(KEYINPUT54), .A3(n1211), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
INV_X1 U871 ( .A(KEYINPUT54), .ZN(n1214) );
XNOR2_X1 U872 ( .A(KEYINPUT19), .B(n1210), .ZN(n1213) );
XOR2_X1 U873 ( .A(G140), .B(n1215), .Z(n1210) );
XNOR2_X1 U874 ( .A(n1216), .B(KEYINPUT25), .ZN(n1211) );
NOR2_X1 U875 ( .A1(n1178), .A2(n1217), .ZN(G51) );
NOR2_X1 U876 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U877 ( .A(n1220), .B(KEYINPUT8), .Z(n1219) );
NAND2_X1 U878 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XNOR2_X1 U879 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U880 ( .A(KEYINPUT50), .B(KEYINPUT0), .Z(n1224) );
NOR2_X1 U881 ( .A1(n1221), .A2(n1223), .ZN(n1218) );
AND2_X1 U882 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NAND2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U884 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND3_X1 U885 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1225) );
AND2_X1 U886 ( .A1(n1183), .A2(n1232), .ZN(n1221) );
AND2_X1 U887 ( .A1(G902), .A2(n1233), .ZN(n1183) );
OR2_X1 U888 ( .A1(n1081), .A2(n1143), .ZN(n1233) );
NOR2_X1 U889 ( .A1(n1234), .A2(n1235), .ZN(n1143) );
XOR2_X1 U890 ( .A(n1084), .B(KEYINPUT17), .Z(n1234) );
NAND4_X1 U891 ( .A1(n1150), .A2(n1172), .A3(n1236), .A4(n1173), .ZN(n1081) );
NOR2_X1 U892 ( .A1(n1171), .A2(n1170), .ZN(n1236) );
AND4_X1 U893 ( .A1(n1190), .A2(n1237), .A3(n1238), .A4(n1075), .ZN(n1172) );
NAND3_X1 U894 ( .A1(n1239), .A2(n1139), .A3(n1240), .ZN(n1075) );
NAND3_X1 U895 ( .A1(n1240), .A2(n1139), .A3(n1137), .ZN(n1190) );
AND2_X1 U896 ( .A1(n1241), .A2(n1242), .ZN(n1150) );
AND4_X1 U897 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NOR4_X1 U898 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1241) );
NOR2_X1 U899 ( .A1(n1117), .A2(n1251), .ZN(n1250) );
INV_X1 U900 ( .A(n1252), .ZN(n1249) );
NOR2_X1 U901 ( .A1(n1130), .A2(G952), .ZN(n1178) );
XOR2_X1 U902 ( .A(n1253), .B(n1252), .Z(G48) );
NAND4_X1 U903 ( .A1(n1113), .A2(n1254), .A3(n1137), .A4(n1255), .ZN(n1252) );
XOR2_X1 U904 ( .A(G143), .B(n1248), .Z(G45) );
AND3_X1 U905 ( .A1(n1141), .A2(n1255), .A3(n1256), .ZN(n1248) );
XNOR2_X1 U906 ( .A(n1243), .B(n1257), .ZN(G42) );
NOR2_X1 U907 ( .A1(KEYINPUT15), .A2(n1258), .ZN(n1257) );
NAND3_X1 U908 ( .A1(n1137), .A2(n1142), .A3(n1259), .ZN(n1243) );
XOR2_X1 U909 ( .A(n1247), .B(n1260), .Z(G39) );
NOR2_X1 U910 ( .A1(KEYINPUT40), .A2(n1261), .ZN(n1260) );
AND3_X1 U911 ( .A1(n1259), .A2(n1124), .A3(n1254), .ZN(n1247) );
XOR2_X1 U912 ( .A(n1262), .B(n1246), .Z(G36) );
NAND3_X1 U913 ( .A1(n1259), .A2(n1239), .A3(n1141), .ZN(n1246) );
XOR2_X1 U914 ( .A(n1263), .B(n1245), .Z(G33) );
NAND3_X1 U915 ( .A1(n1259), .A2(n1137), .A3(n1141), .ZN(n1245) );
AND3_X1 U916 ( .A1(n1133), .A2(n1094), .A3(n1255), .ZN(n1259) );
XOR2_X1 U917 ( .A(G128), .B(n1264), .Z(G30) );
NOR2_X1 U918 ( .A1(n1265), .A2(n1117), .ZN(n1264) );
XOR2_X1 U919 ( .A(n1251), .B(KEYINPUT6), .Z(n1265) );
NAND3_X1 U920 ( .A1(n1255), .A2(n1239), .A3(n1254), .ZN(n1251) );
AND2_X1 U921 ( .A1(n1126), .A2(n1266), .ZN(n1255) );
XOR2_X1 U922 ( .A(n1237), .B(n1267), .Z(G3) );
XNOR2_X1 U923 ( .A(G101), .B(KEYINPUT12), .ZN(n1267) );
NAND3_X1 U924 ( .A1(n1240), .A2(n1124), .A3(n1141), .ZN(n1237) );
XOR2_X1 U925 ( .A(n1268), .B(n1244), .Z(G27) );
NAND3_X1 U926 ( .A1(n1113), .A2(n1084), .A3(n1269), .ZN(n1244) );
AND3_X1 U927 ( .A1(n1137), .A2(n1266), .A3(n1142), .ZN(n1269) );
NAND2_X1 U928 ( .A1(n1270), .A2(n1110), .ZN(n1266) );
NAND2_X1 U929 ( .A1(n1152), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U930 ( .A(G900), .B(KEYINPUT39), .ZN(n1152) );
XOR2_X1 U931 ( .A(n1173), .B(n1272), .Z(G24) );
XOR2_X1 U932 ( .A(KEYINPUT37), .B(G122), .Z(n1272) );
NAND4_X1 U933 ( .A1(n1256), .A2(n1084), .A3(n1139), .A4(n1273), .ZN(n1173) );
INV_X1 U934 ( .A(n1103), .ZN(n1139) );
NAND2_X1 U935 ( .A1(n1274), .A2(n1083), .ZN(n1103) );
NOR3_X1 U936 ( .A1(n1090), .A2(n1275), .A3(n1117), .ZN(n1256) );
INV_X1 U937 ( .A(n1113), .ZN(n1117) );
XOR2_X1 U938 ( .A(n1276), .B(n1277), .Z(G21) );
XOR2_X1 U939 ( .A(KEYINPUT48), .B(G119), .Z(n1277) );
NOR2_X1 U940 ( .A1(n1109), .A2(n1235), .ZN(n1276) );
NAND4_X1 U941 ( .A1(n1113), .A2(n1254), .A3(n1124), .A4(n1273), .ZN(n1235) );
NOR2_X1 U942 ( .A1(n1278), .A2(n1083), .ZN(n1254) );
XOR2_X1 U943 ( .A(G116), .B(n1170), .Z(G18) );
AND3_X1 U944 ( .A1(n1113), .A2(n1239), .A3(n1279), .ZN(n1170) );
INV_X1 U945 ( .A(n1122), .ZN(n1239) );
NAND2_X1 U946 ( .A1(n1280), .A2(n1281), .ZN(n1122) );
XOR2_X1 U947 ( .A(KEYINPUT9), .B(n1275), .Z(n1280) );
XNOR2_X1 U948 ( .A(n1282), .B(KEYINPUT42), .ZN(n1113) );
XOR2_X1 U949 ( .A(G113), .B(n1171), .Z(G15) );
AND3_X1 U950 ( .A1(n1137), .A2(n1282), .A3(n1279), .ZN(n1171) );
AND3_X1 U951 ( .A1(n1084), .A2(n1273), .A3(n1141), .ZN(n1279) );
NOR2_X1 U952 ( .A1(n1283), .A2(n1083), .ZN(n1141) );
INV_X1 U953 ( .A(n1274), .ZN(n1283) );
XNOR2_X1 U954 ( .A(n1278), .B(KEYINPUT29), .ZN(n1274) );
INV_X1 U955 ( .A(n1109), .ZN(n1084) );
NAND2_X1 U956 ( .A1(n1284), .A2(n1128), .ZN(n1109) );
XOR2_X1 U957 ( .A(n1215), .B(n1238), .Z(G12) );
NAND3_X1 U958 ( .A1(n1240), .A2(n1124), .A3(n1142), .ZN(n1238) );
AND2_X1 U959 ( .A1(n1083), .A2(n1285), .ZN(n1142) );
XOR2_X1 U960 ( .A(KEYINPUT59), .B(n1278), .Z(n1285) );
XNOR2_X1 U961 ( .A(n1091), .B(n1286), .ZN(n1278) );
NOR2_X1 U962 ( .A1(n1093), .A2(KEYINPUT23), .ZN(n1286) );
AND2_X1 U963 ( .A1(G217), .A2(n1287), .ZN(n1093) );
OR2_X1 U964 ( .A1(n1181), .A2(G902), .ZN(n1091) );
XNOR2_X1 U965 ( .A(n1288), .B(n1289), .ZN(n1181) );
XOR2_X1 U966 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U967 ( .A(n1292), .B(n1293), .ZN(n1291) );
NOR2_X1 U968 ( .A1(KEYINPUT57), .A2(n1258), .ZN(n1293) );
INV_X1 U969 ( .A(G140), .ZN(n1258) );
NOR2_X1 U970 ( .A1(KEYINPUT33), .A2(n1294), .ZN(n1292) );
XOR2_X1 U971 ( .A(n1295), .B(n1296), .Z(n1294) );
NOR2_X1 U972 ( .A1(G137), .A2(KEYINPUT14), .ZN(n1296) );
AND3_X1 U973 ( .A1(G221), .A2(n1130), .A3(G234), .ZN(n1295) );
NAND2_X1 U974 ( .A1(n1297), .A2(n1298), .ZN(n1290) );
OR2_X1 U975 ( .A1(n1299), .A2(n1215), .ZN(n1298) );
XOR2_X1 U976 ( .A(n1300), .B(KEYINPUT2), .Z(n1297) );
NAND2_X1 U977 ( .A1(n1299), .A2(n1215), .ZN(n1300) );
XNOR2_X1 U978 ( .A(n1301), .B(n1302), .ZN(n1299) );
NOR2_X1 U979 ( .A1(G119), .A2(KEYINPUT16), .ZN(n1302) );
XOR2_X1 U980 ( .A(n1268), .B(n1303), .Z(n1288) );
XOR2_X1 U981 ( .A(KEYINPUT18), .B(G146), .Z(n1303) );
XOR2_X1 U982 ( .A(n1304), .B(G472), .Z(n1083) );
NAND2_X1 U983 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U984 ( .A(n1307), .B(n1308), .Z(n1305) );
XOR2_X1 U985 ( .A(n1198), .B(G101), .Z(n1308) );
NAND3_X1 U986 ( .A1(n1309), .A2(n1310), .A3(G210), .ZN(n1198) );
XOR2_X1 U987 ( .A(KEYINPUT38), .B(G953), .Z(n1309) );
NAND2_X1 U988 ( .A1(n1311), .A2(n1312), .ZN(n1307) );
NAND2_X1 U989 ( .A1(n1195), .A2(n1194), .ZN(n1312) );
NAND2_X1 U990 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
INV_X1 U991 ( .A(n1194), .ZN(n1314) );
XNOR2_X1 U992 ( .A(KEYINPUT45), .B(n1195), .ZN(n1313) );
XOR2_X1 U993 ( .A(n1315), .B(n1316), .Z(n1195) );
NOR2_X1 U994 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
INV_X1 U995 ( .A(n1319), .ZN(n1317) );
NAND2_X1 U996 ( .A1(n1320), .A2(n1321), .ZN(n1124) );
OR3_X1 U997 ( .A1(n1322), .A2(n1281), .A3(KEYINPUT9), .ZN(n1321) );
NAND2_X1 U998 ( .A1(KEYINPUT9), .A2(n1137), .ZN(n1320) );
NOR2_X1 U999 ( .A1(n1281), .A2(n1275), .ZN(n1137) );
INV_X1 U1000 ( .A(n1322), .ZN(n1275) );
NAND2_X1 U1001 ( .A1(n1095), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1002 ( .A1(G475), .A2(n1100), .ZN(n1323) );
OR2_X1 U1003 ( .A1(n1100), .A2(G475), .ZN(n1095) );
NAND2_X1 U1004 ( .A1(n1189), .A2(n1306), .ZN(n1100) );
XNOR2_X1 U1005 ( .A(n1324), .B(n1325), .ZN(n1189) );
XOR2_X1 U1006 ( .A(G104), .B(n1326), .Z(n1325) );
NOR2_X1 U1007 ( .A1(KEYINPUT5), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1008 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1009 ( .A(n1253), .B(n1330), .Z(n1329) );
NAND3_X1 U1010 ( .A1(n1331), .A2(n1332), .A3(KEYINPUT10), .ZN(n1330) );
NAND2_X1 U1011 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
INV_X1 U1012 ( .A(KEYINPUT56), .ZN(n1334) );
XOR2_X1 U1013 ( .A(n1263), .B(n1335), .Z(n1333) );
NAND3_X1 U1014 ( .A1(n1335), .A2(n1263), .A3(KEYINPUT56), .ZN(n1331) );
XOR2_X1 U1015 ( .A(G143), .B(n1336), .Z(n1335) );
AND3_X1 U1016 ( .A1(G214), .A2(n1130), .A3(n1310), .ZN(n1336) );
NAND2_X1 U1017 ( .A1(KEYINPUT31), .A2(n1153), .ZN(n1328) );
XOR2_X1 U1018 ( .A(n1268), .B(G140), .Z(n1153) );
XNOR2_X1 U1019 ( .A(G113), .B(n1337), .ZN(n1324) );
XOR2_X1 U1020 ( .A(KEYINPUT30), .B(G122), .Z(n1337) );
INV_X1 U1021 ( .A(n1090), .ZN(n1281) );
XOR2_X1 U1022 ( .A(n1338), .B(G478), .Z(n1090) );
NAND2_X1 U1023 ( .A1(n1186), .A2(n1306), .ZN(n1338) );
XOR2_X1 U1024 ( .A(n1339), .B(n1340), .Z(n1186) );
XOR2_X1 U1025 ( .A(G107), .B(n1341), .Z(n1340) );
XOR2_X1 U1026 ( .A(G122), .B(G116), .Z(n1341) );
XOR2_X1 U1027 ( .A(n1342), .B(n1343), .Z(n1339) );
NOR2_X1 U1028 ( .A1(KEYINPUT46), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1029 ( .A(n1345), .B(n1346), .Z(n1344) );
NOR2_X1 U1030 ( .A1(KEYINPUT60), .A2(n1262), .ZN(n1345) );
INV_X1 U1031 ( .A(G134), .ZN(n1262) );
NAND3_X1 U1032 ( .A1(G234), .A2(n1130), .A3(G217), .ZN(n1342) );
AND3_X1 U1033 ( .A1(n1126), .A2(n1273), .A3(n1282), .ZN(n1240) );
NOR2_X1 U1034 ( .A1(n1133), .A2(n1118), .ZN(n1282) );
INV_X1 U1035 ( .A(n1094), .ZN(n1118) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1347), .ZN(n1094) );
INV_X1 U1037 ( .A(n1114), .ZN(n1133) );
NAND2_X1 U1038 ( .A1(n1101), .A2(n1096), .ZN(n1114) );
NAND2_X1 U1039 ( .A1(n1232), .A2(n1348), .ZN(n1096) );
NAND2_X1 U1040 ( .A1(n1349), .A2(n1306), .ZN(n1348) );
INV_X1 U1041 ( .A(n1350), .ZN(n1232) );
NAND3_X1 U1042 ( .A1(n1350), .A2(n1306), .A3(n1349), .ZN(n1101) );
XOR2_X1 U1043 ( .A(n1351), .B(n1227), .Z(n1349) );
INV_X1 U1044 ( .A(n1231), .ZN(n1227) );
XNOR2_X1 U1045 ( .A(n1175), .B(n1352), .ZN(n1231) );
NOR2_X1 U1046 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NOR2_X1 U1047 ( .A1(n1355), .A2(n1177), .ZN(n1354) );
INV_X1 U1048 ( .A(n1356), .ZN(n1177) );
NOR2_X1 U1049 ( .A1(KEYINPUT58), .A2(n1357), .ZN(n1355) );
NOR2_X1 U1050 ( .A1(KEYINPUT34), .A2(n1358), .ZN(n1357) );
NOR2_X1 U1051 ( .A1(n1359), .A2(n1360), .ZN(n1353) );
INV_X1 U1052 ( .A(n1358), .ZN(n1360) );
XOR2_X1 U1053 ( .A(n1176), .B(KEYINPUT13), .Z(n1358) );
NAND2_X1 U1054 ( .A1(n1361), .A2(n1362), .ZN(n1176) );
NAND2_X1 U1055 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1056 ( .A(KEYINPUT41), .B(n1365), .Z(n1361) );
NOR2_X1 U1057 ( .A1(n1363), .A2(n1364), .ZN(n1365) );
XNOR2_X1 U1058 ( .A(n1366), .B(KEYINPUT11), .ZN(n1364) );
XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(G101), .ZN(n1363) );
NOR2_X1 U1060 ( .A1(n1367), .A2(KEYINPUT34), .ZN(n1359) );
NOR2_X1 U1061 ( .A1(KEYINPUT58), .A2(n1356), .ZN(n1367) );
NAND3_X1 U1062 ( .A1(n1368), .A2(n1369), .A3(n1319), .ZN(n1356) );
NAND3_X1 U1063 ( .A1(G113), .A2(n1370), .A3(G116), .ZN(n1319) );
NAND2_X1 U1064 ( .A1(n1371), .A2(n1372), .ZN(n1369) );
INV_X1 U1065 ( .A(KEYINPUT44), .ZN(n1372) );
XOR2_X1 U1066 ( .A(G113), .B(n1373), .Z(n1371) );
NOR2_X1 U1067 ( .A1(G116), .A2(n1370), .ZN(n1373) );
INV_X1 U1068 ( .A(G119), .ZN(n1370) );
NAND2_X1 U1069 ( .A1(KEYINPUT44), .A2(n1318), .ZN(n1368) );
NAND2_X1 U1070 ( .A1(n1374), .A2(n1375), .ZN(n1318) );
OR3_X1 U1071 ( .A1(G113), .A2(G116), .A3(G119), .ZN(n1375) );
NAND2_X1 U1072 ( .A1(n1376), .A2(G119), .ZN(n1374) );
XOR2_X1 U1073 ( .A(G116), .B(G113), .Z(n1376) );
XOR2_X1 U1074 ( .A(n1377), .B(n1215), .Z(n1175) );
INV_X1 U1075 ( .A(G122), .ZN(n1377) );
AND2_X1 U1076 ( .A1(n1378), .A2(n1230), .ZN(n1351) );
NAND3_X1 U1077 ( .A1(G224), .A2(n1130), .A3(n1379), .ZN(n1230) );
XOR2_X1 U1078 ( .A(n1315), .B(G125), .Z(n1379) );
XNOR2_X1 U1079 ( .A(KEYINPUT51), .B(n1229), .ZN(n1378) );
NAND2_X1 U1080 ( .A1(n1380), .A2(n1381), .ZN(n1229) );
NAND2_X1 U1081 ( .A1(G224), .A2(n1130), .ZN(n1381) );
XOR2_X1 U1082 ( .A(n1268), .B(n1315), .Z(n1380) );
XOR2_X1 U1083 ( .A(n1382), .B(n1383), .Z(n1315) );
XOR2_X1 U1084 ( .A(KEYINPUT49), .B(KEYINPUT24), .Z(n1383) );
XOR2_X1 U1085 ( .A(n1253), .B(n1346), .Z(n1382) );
XOR2_X1 U1086 ( .A(G128), .B(G143), .Z(n1346) );
INV_X1 U1087 ( .A(G146), .ZN(n1253) );
INV_X1 U1088 ( .A(G125), .ZN(n1268) );
NAND2_X1 U1089 ( .A1(G210), .A2(n1347), .ZN(n1350) );
NAND2_X1 U1090 ( .A1(n1310), .A2(n1306), .ZN(n1347) );
INV_X1 U1091 ( .A(G237), .ZN(n1310) );
NAND2_X1 U1092 ( .A1(n1110), .A2(n1384), .ZN(n1273) );
NAND2_X1 U1093 ( .A1(n1271), .A2(n1385), .ZN(n1384) );
INV_X1 U1094 ( .A(G898), .ZN(n1385) );
AND3_X1 U1095 ( .A1(G902), .A2(n1386), .A3(G953), .ZN(n1271) );
NAND3_X1 U1096 ( .A1(n1386), .A2(n1130), .A3(G952), .ZN(n1110) );
NAND2_X1 U1097 ( .A1(G237), .A2(G234), .ZN(n1386) );
AND2_X1 U1098 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U1099 ( .A1(G221), .A2(n1287), .ZN(n1128) );
NAND2_X1 U1100 ( .A1(G234), .A2(n1306), .ZN(n1287) );
INV_X1 U1101 ( .A(n1284), .ZN(n1127) );
XOR2_X1 U1102 ( .A(n1387), .B(G469), .Z(n1284) );
NAND2_X1 U1103 ( .A1(n1388), .A2(n1306), .ZN(n1387) );
INV_X1 U1104 ( .A(G902), .ZN(n1306) );
XOR2_X1 U1105 ( .A(n1389), .B(n1203), .Z(n1388) );
XOR2_X1 U1106 ( .A(n1158), .B(n1194), .Z(n1203) );
XOR2_X1 U1107 ( .A(n1390), .B(n1391), .Z(n1194) );
NOR2_X1 U1108 ( .A1(KEYINPUT21), .A2(n1263), .ZN(n1391) );
INV_X1 U1109 ( .A(G131), .ZN(n1263) );
NAND3_X1 U1110 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1390) );
NAND2_X1 U1111 ( .A1(KEYINPUT47), .A2(G134), .ZN(n1394) );
NAND3_X1 U1112 ( .A1(n1395), .A2(n1396), .A3(n1261), .ZN(n1393) );
INV_X1 U1113 ( .A(KEYINPUT47), .ZN(n1396) );
OR2_X1 U1114 ( .A1(n1261), .A2(n1395), .ZN(n1392) );
NOR2_X1 U1115 ( .A1(G134), .A2(KEYINPUT43), .ZN(n1395) );
INV_X1 U1116 ( .A(G137), .ZN(n1261) );
NAND2_X1 U1117 ( .A1(n1397), .A2(n1398), .ZN(n1158) );
OR2_X1 U1118 ( .A1(n1399), .A2(n1301), .ZN(n1398) );
XOR2_X1 U1119 ( .A(n1400), .B(KEYINPUT55), .Z(n1397) );
NAND2_X1 U1120 ( .A1(n1399), .A2(n1301), .ZN(n1400) );
INV_X1 U1121 ( .A(G128), .ZN(n1301) );
XNOR2_X1 U1122 ( .A(n1401), .B(G146), .ZN(n1399) );
NAND2_X1 U1123 ( .A1(KEYINPUT7), .A2(n1402), .ZN(n1401) );
XOR2_X1 U1124 ( .A(KEYINPUT49), .B(G143), .Z(n1402) );
XOR2_X1 U1125 ( .A(n1403), .B(n1404), .Z(n1389) );
NOR2_X1 U1126 ( .A1(KEYINPUT62), .A2(n1204), .ZN(n1404) );
XOR2_X1 U1127 ( .A(G101), .B(n1366), .Z(n1204) );
XNOR2_X1 U1128 ( .A(G104), .B(G107), .ZN(n1366) );
NAND2_X1 U1129 ( .A1(KEYINPUT52), .A2(n1405), .ZN(n1403) );
XOR2_X1 U1130 ( .A(n1406), .B(n1407), .Z(n1405) );
XOR2_X1 U1131 ( .A(G110), .B(n1216), .Z(n1407) );
AND2_X1 U1132 ( .A1(G227), .A2(n1130), .ZN(n1216) );
INV_X1 U1133 ( .A(G953), .ZN(n1130) );
NOR2_X1 U1134 ( .A1(G140), .A2(KEYINPUT26), .ZN(n1406) );
INV_X1 U1135 ( .A(G110), .ZN(n1215) );
endmodule


