//Key = 1010101100111011011011000000011110000001000110000000100001001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353;

XNOR2_X1 U745 ( .A(G107), .B(n1022), .ZN(G9) );
NAND4_X1 U746 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NOR2_X1 U747 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
XOR2_X1 U748 ( .A(n1029), .B(KEYINPUT37), .Z(n1028) );
NOR2_X1 U749 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U751 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U752 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR3_X1 U754 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1039) );
NOR3_X1 U755 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
INV_X1 U756 ( .A(KEYINPUT24), .ZN(n1046) );
NOR2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1042) );
NOR3_X1 U758 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1047) );
NOR2_X1 U759 ( .A1(KEYINPUT24), .A2(n1045), .ZN(n1051) );
NAND3_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1050) );
NOR2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
XOR2_X1 U764 ( .A(n1061), .B(KEYINPUT9), .Z(n1059) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1049) );
NOR3_X1 U766 ( .A1(n1063), .A2(n1064), .A3(n1056), .ZN(n1041) );
NOR2_X1 U767 ( .A1(n1024), .A2(n1065), .ZN(n1064) );
NOR4_X1 U768 ( .A1(n1066), .A2(n1048), .A3(n1056), .A4(n1063), .ZN(n1037) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U771 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U772 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1032) );
NOR4_X1 U773 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U775 ( .A1(KEYINPUT19), .A2(n1081), .ZN(n1079) );
XOR2_X1 U776 ( .A(KEYINPUT49), .B(G472), .Z(n1081) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(n1077) );
XNOR2_X1 U778 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND2_X1 U779 ( .A1(KEYINPUT20), .A2(G478), .ZN(n1085) );
XNOR2_X1 U780 ( .A(KEYINPUT62), .B(KEYINPUT48), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1060), .A2(n1086), .ZN(n1076) );
NOR3_X1 U782 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1073) );
AND2_X1 U783 ( .A1(G472), .A2(KEYINPUT19), .ZN(n1089) );
NOR3_X1 U784 ( .A1(KEYINPUT19), .A2(G472), .A3(n1090), .ZN(n1088) );
INV_X1 U785 ( .A(n1080), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1091), .B(KEYINPUT21), .Z(n1080) );
XOR2_X1 U787 ( .A(G469), .B(n1092), .Z(n1087) );
XOR2_X1 U788 ( .A(n1093), .B(n1094), .Z(n1071) );
XOR2_X1 U789 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U790 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U791 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U792 ( .A1(G953), .A2(n1101), .ZN(n1100) );
XNOR2_X1 U793 ( .A(n1102), .B(n1103), .ZN(n1099) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND3_X1 U796 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1104) );
OR2_X1 U797 ( .A1(n1111), .A2(G131), .ZN(n1110) );
NAND2_X1 U798 ( .A1(KEYINPUT36), .A2(n1112), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1111), .ZN(n1112) );
XNOR2_X1 U800 ( .A(KEYINPUT14), .B(G131), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1114), .A2(n1115), .ZN(n1108) );
INV_X1 U802 ( .A(KEYINPUT36), .ZN(n1115) );
NAND2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
OR2_X1 U804 ( .A1(G131), .A2(KEYINPUT14), .ZN(n1117) );
NAND3_X1 U805 ( .A1(G131), .A2(n1111), .A3(KEYINPUT14), .ZN(n1116) );
NAND2_X1 U806 ( .A1(n1118), .A2(G953), .ZN(n1097) );
XOR2_X1 U807 ( .A(n1119), .B(KEYINPUT33), .Z(n1118) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1119) );
NOR2_X1 U809 ( .A1(n1120), .A2(G953), .ZN(n1095) );
NOR2_X1 U810 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND3_X1 U811 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(G69) );
NAND2_X1 U812 ( .A1(G953), .A2(n1126), .ZN(n1125) );
NAND2_X1 U813 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U815 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1127) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1131) );
NAND2_X1 U817 ( .A1(n1133), .A2(n1130), .ZN(n1124) );
INV_X1 U818 ( .A(KEYINPUT60), .ZN(n1130) );
NAND3_X1 U819 ( .A1(n1134), .A2(n1135), .A3(KEYINPUT60), .ZN(n1123) );
NAND3_X1 U820 ( .A1(n1129), .A2(n1132), .A3(G953), .ZN(n1135) );
INV_X1 U821 ( .A(KEYINPUT35), .ZN(n1132) );
INV_X1 U822 ( .A(G224), .ZN(n1129) );
INV_X1 U823 ( .A(n1133), .ZN(n1134) );
XOR2_X1 U824 ( .A(n1136), .B(n1137), .Z(n1133) );
NOR4_X1 U825 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
NOR2_X1 U826 ( .A1(G898), .A2(n1142), .ZN(n1141) );
NOR2_X1 U827 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
NOR2_X1 U828 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
INV_X1 U829 ( .A(KEYINPUT6), .ZN(n1146) );
NOR2_X1 U830 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NOR2_X1 U831 ( .A1(KEYINPUT11), .A2(n1144), .ZN(n1148) );
AND3_X1 U832 ( .A1(n1144), .A2(n1143), .A3(KEYINPUT11), .ZN(n1147) );
NOR2_X1 U833 ( .A1(KEYINPUT6), .A2(n1149), .ZN(n1138) );
NOR2_X1 U834 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
INV_X1 U835 ( .A(n1143), .ZN(n1151) );
XOR2_X1 U836 ( .A(n1152), .B(n1153), .Z(n1143) );
NOR2_X1 U837 ( .A1(KEYINPUT40), .A2(n1154), .ZN(n1153) );
XOR2_X1 U838 ( .A(n1144), .B(KEYINPUT11), .Z(n1150) );
NAND2_X1 U839 ( .A1(n1142), .A2(n1155), .ZN(n1136) );
NOR2_X1 U840 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XOR2_X1 U841 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U842 ( .A(n1160), .B(KEYINPUT51), .Z(n1158) );
NAND2_X1 U843 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U844 ( .A1(n1156), .A2(n1163), .ZN(G63) );
NOR3_X1 U845 ( .A1(n1084), .A2(n1164), .A3(n1165), .ZN(n1163) );
NOR3_X1 U846 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
AND2_X1 U847 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NAND2_X1 U848 ( .A1(n1169), .A2(G478), .ZN(n1166) );
XOR2_X1 U849 ( .A(n1034), .B(KEYINPUT26), .Z(n1169) );
NOR2_X1 U850 ( .A1(n1156), .A2(n1170), .ZN(G60) );
XOR2_X1 U851 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U852 ( .A1(KEYINPUT34), .A2(n1173), .ZN(n1172) );
NAND2_X1 U853 ( .A1(n1161), .A2(G475), .ZN(n1171) );
XNOR2_X1 U854 ( .A(G104), .B(n1174), .ZN(G6) );
NOR2_X1 U855 ( .A1(n1156), .A2(n1175), .ZN(G57) );
XOR2_X1 U856 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U857 ( .A(n1178), .B(KEYINPUT42), .ZN(n1177) );
NAND2_X1 U858 ( .A1(KEYINPUT10), .A2(n1179), .ZN(n1178) );
XOR2_X1 U859 ( .A(n1180), .B(n1181), .Z(n1176) );
NAND2_X1 U860 ( .A1(n1161), .A2(G472), .ZN(n1180) );
NOR2_X1 U861 ( .A1(n1156), .A2(n1182), .ZN(G54) );
XOR2_X1 U862 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U863 ( .A1(n1161), .A2(G469), .ZN(n1184) );
INV_X1 U864 ( .A(n1185), .ZN(n1161) );
NAND2_X1 U865 ( .A1(n1186), .A2(n1187), .ZN(n1183) );
OR2_X1 U866 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U867 ( .A(n1190), .B(KEYINPUT58), .Z(n1186) );
NAND2_X1 U868 ( .A1(n1189), .A2(n1188), .ZN(n1190) );
XNOR2_X1 U869 ( .A(n1191), .B(n1192), .ZN(n1188) );
NAND2_X1 U870 ( .A1(KEYINPUT0), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U871 ( .A(n1194), .B(n1195), .ZN(n1189) );
XOR2_X1 U872 ( .A(n1196), .B(n1197), .Z(n1194) );
NAND2_X1 U873 ( .A1(KEYINPUT43), .A2(n1198), .ZN(n1196) );
NOR2_X1 U874 ( .A1(n1156), .A2(n1199), .ZN(G51) );
XOR2_X1 U875 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U876 ( .A1(n1202), .A2(n1185), .ZN(n1201) );
NAND2_X1 U877 ( .A1(G902), .A2(n1034), .ZN(n1185) );
OR3_X1 U878 ( .A1(n1155), .A2(n1122), .A3(n1203), .ZN(n1034) );
XOR2_X1 U879 ( .A(n1121), .B(KEYINPUT22), .Z(n1203) );
INV_X1 U880 ( .A(n1204), .ZN(n1121) );
NAND4_X1 U881 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1122) );
NOR4_X1 U882 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
OR3_X1 U883 ( .A1(n1056), .A2(n1029), .A3(n1213), .ZN(n1207) );
NAND4_X1 U884 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1155) );
AND4_X1 U885 ( .A1(n1174), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1217) );
NAND3_X1 U886 ( .A1(n1221), .A2(n1026), .A3(n1065), .ZN(n1174) );
NOR3_X1 U887 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1216) );
AND4_X1 U888 ( .A1(KEYINPUT45), .A2(n1225), .A3(n1226), .A4(n1026), .ZN(n1224) );
NAND2_X1 U889 ( .A1(n1227), .A2(n1075), .ZN(n1226) );
NOR2_X1 U890 ( .A1(KEYINPUT45), .A2(n1228), .ZN(n1223) );
NAND3_X1 U891 ( .A1(n1024), .A2(n1026), .A3(n1221), .ZN(n1214) );
NAND2_X1 U892 ( .A1(n1229), .A2(KEYINPUT39), .ZN(n1200) );
XOR2_X1 U893 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U894 ( .A1(n1142), .A2(G952), .ZN(n1156) );
XNOR2_X1 U895 ( .A(G146), .B(n1205), .ZN(G48) );
NAND3_X1 U896 ( .A1(n1065), .A2(n1058), .A3(n1232), .ZN(n1205) );
XOR2_X1 U897 ( .A(n1233), .B(n1206), .Z(G45) );
NAND4_X1 U898 ( .A1(n1075), .A2(n1234), .A3(n1058), .A4(n1227), .ZN(n1206) );
XOR2_X1 U899 ( .A(G140), .B(n1235), .Z(G42) );
NOR2_X1 U900 ( .A1(KEYINPUT5), .A2(n1236), .ZN(n1235) );
INV_X1 U901 ( .A(n1212), .ZN(n1236) );
NOR3_X1 U902 ( .A1(n1063), .A2(n1062), .A3(n1213), .ZN(n1212) );
XOR2_X1 U903 ( .A(G137), .B(n1211), .Z(G39) );
AND3_X1 U904 ( .A1(n1232), .A2(n1044), .A3(n1052), .ZN(n1211) );
XOR2_X1 U905 ( .A(n1237), .B(n1204), .Z(G36) );
NAND3_X1 U906 ( .A1(n1234), .A2(n1024), .A3(n1052), .ZN(n1204) );
XOR2_X1 U907 ( .A(G131), .B(n1210), .Z(G33) );
AND3_X1 U908 ( .A1(n1234), .A2(n1065), .A3(n1052), .ZN(n1210) );
INV_X1 U909 ( .A(n1063), .ZN(n1052) );
NAND2_X1 U910 ( .A1(n1238), .A2(n1060), .ZN(n1063) );
INV_X1 U911 ( .A(n1061), .ZN(n1238) );
AND3_X1 U912 ( .A1(n1023), .A2(n1239), .A3(n1068), .ZN(n1234) );
XOR2_X1 U913 ( .A(G128), .B(n1209), .Z(G30) );
AND3_X1 U914 ( .A1(n1024), .A2(n1058), .A3(n1232), .ZN(n1209) );
AND4_X1 U915 ( .A1(n1023), .A2(n1240), .A3(n1069), .A4(n1239), .ZN(n1232) );
NAND2_X1 U916 ( .A1(n1241), .A2(n1242), .ZN(G3) );
NAND2_X1 U917 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U918 ( .A(G101), .ZN(n1244) );
XOR2_X1 U919 ( .A(n1245), .B(KEYINPUT55), .Z(n1243) );
NAND2_X1 U920 ( .A1(n1246), .A2(G101), .ZN(n1241) );
XOR2_X1 U921 ( .A(n1245), .B(KEYINPUT7), .Z(n1246) );
NAND2_X1 U922 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
NAND2_X1 U923 ( .A1(n1222), .A2(n1249), .ZN(n1248) );
INV_X1 U924 ( .A(KEYINPUT27), .ZN(n1249) );
AND3_X1 U925 ( .A1(n1044), .A2(n1221), .A3(n1068), .ZN(n1222) );
NAND4_X1 U926 ( .A1(n1068), .A2(n1044), .A3(n1250), .A4(KEYINPUT27), .ZN(n1247) );
NOR3_X1 U927 ( .A1(n1062), .A2(n1058), .A3(n1027), .ZN(n1250) );
INV_X1 U928 ( .A(n1029), .ZN(n1058) );
XOR2_X1 U929 ( .A(G125), .B(n1251), .Z(G27) );
NOR3_X1 U930 ( .A1(n1252), .A2(n1029), .A3(n1213), .ZN(n1251) );
NAND4_X1 U931 ( .A1(n1070), .A2(n1065), .A3(n1069), .A4(n1239), .ZN(n1213) );
NAND2_X1 U932 ( .A1(n1253), .A2(n1254), .ZN(n1239) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1101), .ZN(n1254) );
INV_X1 U934 ( .A(G900), .ZN(n1101) );
XNOR2_X1 U935 ( .A(KEYINPUT4), .B(n1056), .ZN(n1252) );
XOR2_X1 U936 ( .A(n1256), .B(n1228), .Z(G24) );
NAND4_X1 U937 ( .A1(n1075), .A2(n1225), .A3(n1026), .A4(n1227), .ZN(n1228) );
INV_X1 U938 ( .A(n1040), .ZN(n1026) );
NAND2_X1 U939 ( .A1(n1070), .A2(n1072), .ZN(n1040) );
XOR2_X1 U940 ( .A(n1257), .B(n1215), .Z(G21) );
NAND4_X1 U941 ( .A1(n1225), .A2(n1044), .A3(n1240), .A4(n1069), .ZN(n1215) );
XNOR2_X1 U942 ( .A(G116), .B(n1220), .ZN(G18) );
NAND3_X1 U943 ( .A1(n1068), .A2(n1024), .A3(n1225), .ZN(n1220) );
NOR2_X1 U944 ( .A1(n1075), .A2(n1258), .ZN(n1024) );
XOR2_X1 U945 ( .A(n1259), .B(n1219), .Z(G15) );
NAND3_X1 U946 ( .A1(n1068), .A2(n1065), .A3(n1225), .ZN(n1219) );
NOR3_X1 U947 ( .A1(n1029), .A2(n1027), .A3(n1056), .ZN(n1225) );
NAND2_X1 U948 ( .A1(n1053), .A2(n1086), .ZN(n1056) );
NOR2_X1 U949 ( .A1(n1227), .A2(n1260), .ZN(n1065) );
INV_X1 U950 ( .A(n1258), .ZN(n1227) );
AND2_X1 U951 ( .A1(n1072), .A2(n1240), .ZN(n1068) );
XNOR2_X1 U952 ( .A(n1070), .B(KEYINPUT41), .ZN(n1240) );
XOR2_X1 U953 ( .A(n1198), .B(n1218), .Z(G12) );
NAND4_X1 U954 ( .A1(n1044), .A2(n1221), .A3(n1070), .A4(n1069), .ZN(n1218) );
INV_X1 U955 ( .A(n1072), .ZN(n1069) );
XOR2_X1 U956 ( .A(n1261), .B(n1162), .Z(n1072) );
AND2_X1 U957 ( .A1(G217), .A2(n1262), .ZN(n1162) );
NAND2_X1 U958 ( .A1(n1159), .A2(n1168), .ZN(n1261) );
XNOR2_X1 U959 ( .A(n1263), .B(n1264), .ZN(n1159) );
XOR2_X1 U960 ( .A(G119), .B(n1265), .Z(n1264) );
XOR2_X1 U961 ( .A(G137), .B(G128), .Z(n1265) );
XOR2_X1 U962 ( .A(n1266), .B(n1267), .Z(n1263) );
AND3_X1 U963 ( .A1(G221), .A2(n1142), .A3(G234), .ZN(n1267) );
XOR2_X1 U964 ( .A(n1198), .B(n1268), .Z(n1266) );
NOR2_X1 U965 ( .A1(KEYINPUT46), .A2(n1269), .ZN(n1268) );
XOR2_X1 U966 ( .A(n1270), .B(G146), .Z(n1269) );
NAND3_X1 U967 ( .A1(n1271), .A2(n1272), .A3(n1106), .ZN(n1270) );
INV_X1 U968 ( .A(n1273), .ZN(n1106) );
OR2_X1 U969 ( .A1(n1107), .A2(KEYINPUT28), .ZN(n1272) );
NAND2_X1 U970 ( .A1(KEYINPUT28), .A2(G140), .ZN(n1271) );
XOR2_X1 U971 ( .A(n1091), .B(G472), .Z(n1070) );
NAND2_X1 U972 ( .A1(n1274), .A2(n1168), .ZN(n1091) );
XOR2_X1 U973 ( .A(n1181), .B(n1179), .Z(n1274) );
XOR2_X1 U974 ( .A(n1275), .B(n1276), .Z(n1179) );
XNOR2_X1 U975 ( .A(n1277), .B(n1278), .ZN(n1181) );
XOR2_X1 U976 ( .A(n1279), .B(n1280), .Z(n1278) );
AND3_X1 U977 ( .A1(G210), .A2(n1142), .A3(n1281), .ZN(n1279) );
XOR2_X1 U978 ( .A(n1259), .B(n1282), .Z(n1277) );
NOR2_X1 U979 ( .A1(KEYINPUT3), .A2(n1283), .ZN(n1282) );
NOR3_X1 U980 ( .A1(n1029), .A2(n1027), .A3(n1062), .ZN(n1221) );
INV_X1 U981 ( .A(n1023), .ZN(n1062) );
NOR2_X1 U982 ( .A1(n1053), .A2(n1054), .ZN(n1023) );
INV_X1 U983 ( .A(n1086), .ZN(n1054) );
NAND2_X1 U984 ( .A1(G221), .A2(n1262), .ZN(n1086) );
NAND2_X1 U985 ( .A1(n1284), .A2(n1168), .ZN(n1262) );
XOR2_X1 U986 ( .A(KEYINPUT23), .B(G234), .Z(n1284) );
XOR2_X1 U987 ( .A(G469), .B(n1285), .Z(n1053) );
NOR2_X1 U988 ( .A1(n1092), .A2(KEYINPUT38), .ZN(n1285) );
AND2_X1 U989 ( .A1(n1286), .A2(n1168), .ZN(n1092) );
XOR2_X1 U990 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U991 ( .A(n1289), .B(n1192), .Z(n1288) );
XNOR2_X1 U992 ( .A(n1275), .B(n1102), .ZN(n1192) );
XOR2_X1 U993 ( .A(n1290), .B(n1291), .Z(n1102) );
XNOR2_X1 U994 ( .A(G128), .B(KEYINPUT54), .ZN(n1290) );
XNOR2_X1 U995 ( .A(G131), .B(n1111), .ZN(n1275) );
XNOR2_X1 U996 ( .A(n1237), .B(G137), .ZN(n1111) );
XOR2_X1 U997 ( .A(n1152), .B(n1197), .Z(n1289) );
AND2_X1 U998 ( .A1(G227), .A2(n1142), .ZN(n1197) );
XOR2_X1 U999 ( .A(n1292), .B(n1293), .Z(n1287) );
NOR2_X1 U1000 ( .A1(KEYINPUT61), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1001 ( .A(G110), .B(n1195), .Z(n1294) );
XOR2_X1 U1002 ( .A(G140), .B(KEYINPUT15), .Z(n1195) );
XNOR2_X1 U1003 ( .A(KEYINPUT50), .B(KEYINPUT30), .ZN(n1292) );
AND2_X1 U1004 ( .A1(n1295), .A2(n1253), .ZN(n1027) );
NAND3_X1 U1005 ( .A1(n1255), .A2(n1142), .A3(n1296), .ZN(n1253) );
XNOR2_X1 U1006 ( .A(G952), .B(KEYINPUT32), .ZN(n1296) );
XOR2_X1 U1007 ( .A(n1297), .B(KEYINPUT53), .Z(n1295) );
OR4_X1 U1008 ( .A1(n1142), .A2(n1168), .A3(n1035), .A4(G898), .ZN(n1297) );
INV_X1 U1009 ( .A(n1255), .ZN(n1035) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1255) );
NAND2_X1 U1011 ( .A1(n1061), .A2(n1060), .ZN(n1029) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1298), .ZN(n1060) );
XOR2_X1 U1013 ( .A(n1093), .B(n1299), .Z(n1061) );
NOR2_X1 U1014 ( .A1(n1094), .A2(KEYINPUT16), .ZN(n1299) );
INV_X1 U1015 ( .A(n1202), .ZN(n1094) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1298), .ZN(n1202) );
NAND2_X1 U1017 ( .A1(n1281), .A2(n1168), .ZN(n1298) );
NAND3_X1 U1018 ( .A1(n1300), .A2(n1168), .A3(n1301), .ZN(n1093) );
NAND3_X1 U1019 ( .A1(n1302), .A2(n1303), .A3(KEYINPUT31), .ZN(n1301) );
NAND2_X1 U1020 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
INV_X1 U1021 ( .A(n1230), .ZN(n1304) );
NAND2_X1 U1022 ( .A1(n1230), .A2(n1306), .ZN(n1302) );
NAND2_X1 U1023 ( .A1(n1231), .A2(n1305), .ZN(n1306) );
INV_X1 U1024 ( .A(KEYINPUT25), .ZN(n1305) );
INV_X1 U1025 ( .A(n1307), .ZN(n1231) );
NAND2_X1 U1026 ( .A1(n1307), .A2(n1308), .ZN(n1300) );
NAND2_X1 U1027 ( .A1(n1230), .A2(n1309), .ZN(n1308) );
OR2_X1 U1028 ( .A1(KEYINPUT25), .A2(KEYINPUT31), .ZN(n1309) );
XOR2_X1 U1029 ( .A(n1310), .B(n1276), .Z(n1230) );
XNOR2_X1 U1030 ( .A(n1291), .B(n1311), .ZN(n1276) );
NOR2_X1 U1031 ( .A1(G128), .A2(KEYINPUT13), .ZN(n1311) );
XNOR2_X1 U1032 ( .A(G143), .B(G146), .ZN(n1291) );
XOR2_X1 U1033 ( .A(n1312), .B(n1313), .Z(n1310) );
NAND2_X1 U1034 ( .A1(G224), .A2(n1142), .ZN(n1312) );
XOR2_X1 U1035 ( .A(n1314), .B(n1193), .Z(n1307) );
INV_X1 U1036 ( .A(n1152), .ZN(n1193) );
XOR2_X1 U1037 ( .A(n1315), .B(n1316), .Z(n1152) );
XOR2_X1 U1038 ( .A(KEYINPUT57), .B(G107), .Z(n1316) );
XNOR2_X1 U1039 ( .A(G104), .B(n1280), .ZN(n1315) );
XOR2_X1 U1040 ( .A(G101), .B(KEYINPUT56), .Z(n1280) );
XOR2_X1 U1041 ( .A(n1154), .B(n1317), .Z(n1314) );
NOR2_X1 U1042 ( .A1(KEYINPUT63), .A2(n1144), .ZN(n1317) );
NAND3_X1 U1043 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1144) );
NAND2_X1 U1044 ( .A1(G110), .A2(n1256), .ZN(n1320) );
NAND2_X1 U1045 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
INV_X1 U1046 ( .A(KEYINPUT17), .ZN(n1322) );
NAND2_X1 U1047 ( .A1(n1323), .A2(n1198), .ZN(n1321) );
XOR2_X1 U1048 ( .A(KEYINPUT47), .B(G122), .Z(n1323) );
NAND2_X1 U1049 ( .A1(KEYINPUT17), .A2(n1324), .ZN(n1318) );
NAND2_X1 U1050 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
OR3_X1 U1051 ( .A1(n1256), .A2(G110), .A3(KEYINPUT47), .ZN(n1326) );
NAND2_X1 U1052 ( .A1(KEYINPUT47), .A2(n1256), .ZN(n1325) );
XNOR2_X1 U1053 ( .A(n1327), .B(n1283), .ZN(n1154) );
XOR2_X1 U1054 ( .A(G116), .B(n1257), .Z(n1283) );
INV_X1 U1055 ( .A(G119), .ZN(n1257) );
NAND2_X1 U1056 ( .A1(KEYINPUT2), .A2(n1259), .ZN(n1327) );
INV_X1 U1057 ( .A(G113), .ZN(n1259) );
INV_X1 U1058 ( .A(n1048), .ZN(n1044) );
NAND2_X1 U1059 ( .A1(n1258), .A2(n1260), .ZN(n1048) );
INV_X1 U1060 ( .A(n1075), .ZN(n1260) );
XOR2_X1 U1061 ( .A(n1328), .B(n1329), .Z(n1075) );
XOR2_X1 U1062 ( .A(KEYINPUT12), .B(G475), .Z(n1329) );
OR2_X1 U1063 ( .A1(n1173), .A2(G902), .ZN(n1328) );
XNOR2_X1 U1064 ( .A(n1330), .B(n1331), .ZN(n1173) );
XOR2_X1 U1065 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1066 ( .A(n1334), .B(n1335), .Z(n1333) );
NOR3_X1 U1067 ( .A1(n1273), .A2(n1336), .A3(n1337), .ZN(n1335) );
AND2_X1 U1068 ( .A1(G140), .A2(KEYINPUT59), .ZN(n1337) );
NOR2_X1 U1069 ( .A1(KEYINPUT59), .A2(n1107), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(n1313), .A2(n1338), .ZN(n1107) );
NOR2_X1 U1071 ( .A1(n1313), .A2(n1338), .ZN(n1273) );
INV_X1 U1072 ( .A(G140), .ZN(n1338) );
XOR2_X1 U1073 ( .A(G125), .B(KEYINPUT44), .Z(n1313) );
NAND2_X1 U1074 ( .A1(n1339), .A2(n1340), .ZN(n1334) );
NAND2_X1 U1075 ( .A1(n1341), .A2(n1233), .ZN(n1340) );
XOR2_X1 U1076 ( .A(n1342), .B(KEYINPUT8), .Z(n1339) );
OR2_X1 U1077 ( .A1(n1341), .A2(n1233), .ZN(n1342) );
INV_X1 U1078 ( .A(G143), .ZN(n1233) );
NAND3_X1 U1079 ( .A1(n1281), .A2(n1142), .A3(G214), .ZN(n1341) );
INV_X1 U1080 ( .A(G237), .ZN(n1281) );
NAND2_X1 U1081 ( .A1(KEYINPUT29), .A2(G146), .ZN(n1332) );
XOR2_X1 U1082 ( .A(n1343), .B(n1344), .Z(n1330) );
XOR2_X1 U1083 ( .A(G113), .B(n1345), .Z(n1344) );
NOR2_X1 U1084 ( .A1(G104), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(KEYINPUT1), .ZN(n1346) );
XOR2_X1 U1086 ( .A(n1256), .B(G131), .Z(n1343) );
INV_X1 U1087 ( .A(G122), .ZN(n1256) );
XNOR2_X1 U1088 ( .A(n1084), .B(G478), .ZN(n1258) );
AND2_X1 U1089 ( .A1(n1167), .A2(n1168), .ZN(n1084) );
INV_X1 U1090 ( .A(G902), .ZN(n1168) );
XOR2_X1 U1091 ( .A(n1347), .B(n1348), .Z(n1167) );
XOR2_X1 U1092 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1093 ( .A(G122), .B(G116), .Z(n1350) );
XOR2_X1 U1094 ( .A(G143), .B(G128), .Z(n1349) );
XOR2_X1 U1095 ( .A(n1351), .B(n1352), .Z(n1347) );
AND3_X1 U1096 ( .A1(G217), .A2(n1142), .A3(G234), .ZN(n1352) );
INV_X1 U1097 ( .A(G953), .ZN(n1142) );
XOR2_X1 U1098 ( .A(n1353), .B(G107), .Z(n1351) );
NAND2_X1 U1099 ( .A1(KEYINPUT18), .A2(n1237), .ZN(n1353) );
INV_X1 U1100 ( .A(G134), .ZN(n1237) );
INV_X1 U1101 ( .A(G110), .ZN(n1198) );
endmodule


