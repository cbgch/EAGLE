//Key = 0100001010111001001010011010110000111000001101110110011100111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273;

XOR2_X1 U709 ( .A(n970), .B(n971), .Z(G9) );
XOR2_X1 U710 ( .A(KEYINPUT8), .B(G107), .Z(n971) );
NAND4_X1 U711 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(G75) );
NAND4_X1 U712 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n974) );
NOR4_X1 U713 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n979) );
XOR2_X1 U714 ( .A(n984), .B(n985), .Z(n983) );
XNOR2_X1 U715 ( .A(KEYINPUT4), .B(n986), .ZN(n982) );
NOR2_X1 U716 ( .A1(n987), .A2(n988), .ZN(n981) );
XOR2_X1 U717 ( .A(KEYINPUT3), .B(G478), .Z(n987) );
NOR2_X1 U718 ( .A1(n989), .A2(n990), .ZN(n980) );
XNOR2_X1 U719 ( .A(G478), .B(KEYINPUT7), .ZN(n990) );
AND2_X1 U720 ( .A1(n991), .A2(n992), .ZN(n978) );
XOR2_X1 U721 ( .A(n993), .B(n994), .Z(n976) );
XOR2_X1 U722 ( .A(n995), .B(KEYINPUT35), .Z(n994) );
NAND2_X1 U723 ( .A1(n996), .A2(n997), .ZN(n973) );
NAND2_X1 U724 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND3_X1 U725 ( .A1(n991), .A2(n1000), .A3(n1001), .ZN(n999) );
NAND2_X1 U726 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NAND2_X1 U727 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
OR2_X1 U728 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U729 ( .A1(n1008), .A2(n1009), .ZN(n1002) );
NAND2_X1 U730 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U731 ( .A1(n1004), .A2(n1012), .A3(n1008), .ZN(n998) );
NAND2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U733 ( .A1(n1001), .A2(n1015), .ZN(n1014) );
NAND2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U736 ( .A1(n991), .A2(n1020), .ZN(n1013) );
NAND3_X1 U737 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
OR3_X1 U738 ( .A1(n977), .A2(n1024), .A3(KEYINPUT62), .ZN(n1022) );
NAND2_X1 U739 ( .A1(KEYINPUT62), .A2(n977), .ZN(n1021) );
INV_X1 U740 ( .A(n1025), .ZN(n996) );
NAND2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(G72) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U743 ( .A1(G953), .A2(n1030), .ZN(n1029) );
NAND2_X1 U744 ( .A1(G900), .A2(G227), .ZN(n1030) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1026) );
INV_X1 U746 ( .A(n1028), .ZN(n1032) );
NOR2_X1 U747 ( .A1(KEYINPUT5), .A2(n1033), .ZN(n1028) );
XOR2_X1 U748 ( .A(n1034), .B(n1035), .Z(n1033) );
NOR2_X1 U749 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U750 ( .A(n1038), .B(n1039), .Z(n1037) );
XOR2_X1 U751 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U752 ( .A1(KEYINPUT41), .A2(n1042), .ZN(n1040) );
XOR2_X1 U753 ( .A(n1043), .B(n1044), .Z(n1038) );
NOR2_X1 U754 ( .A1(KEYINPUT27), .A2(n1045), .ZN(n1044) );
XOR2_X1 U755 ( .A(n1046), .B(G134), .Z(n1043) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1034) );
XOR2_X1 U757 ( .A(n975), .B(KEYINPUT52), .Z(n1047) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1031) );
NAND2_X1 U759 ( .A1(G953), .A2(n1051), .ZN(n1050) );
INV_X1 U760 ( .A(n1036), .ZN(n1049) );
XOR2_X1 U761 ( .A(n1052), .B(n1053), .Z(G69) );
NAND2_X1 U762 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND2_X1 U764 ( .A1(G898), .A2(G953), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1059), .A2(n975), .ZN(n1056) );
NAND2_X1 U766 ( .A1(KEYINPUT36), .A2(n1060), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1060), .A2(n975), .ZN(n1062) );
XNOR2_X1 U769 ( .A(n1063), .B(KEYINPUT47), .ZN(n1060) );
NAND2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U771 ( .A(n970), .B(KEYINPUT33), .Z(n1064) );
NAND2_X1 U772 ( .A1(KEYINPUT36), .A2(n1058), .ZN(n1061) );
XNOR2_X1 U773 ( .A(n1066), .B(n1067), .ZN(n1058) );
XOR2_X1 U774 ( .A(KEYINPUT32), .B(KEYINPUT28), .Z(n1067) );
XNOR2_X1 U775 ( .A(n1068), .B(KEYINPUT15), .ZN(n1066) );
NAND3_X1 U776 ( .A1(G953), .A2(n1069), .A3(KEYINPUT6), .ZN(n1052) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1069) );
NOR2_X1 U778 ( .A1(n1070), .A2(n1071), .ZN(G66) );
XOR2_X1 U779 ( .A(n1072), .B(n1073), .Z(n1071) );
NAND4_X1 U780 ( .A1(KEYINPUT55), .A2(n1074), .A3(G902), .A4(n1075), .ZN(n1072) );
XOR2_X1 U781 ( .A(KEYINPUT42), .B(n972), .Z(n1075) );
INV_X1 U782 ( .A(n1076), .ZN(n972) );
INV_X1 U783 ( .A(n995), .ZN(n1074) );
NOR2_X1 U784 ( .A1(n1070), .A2(n1077), .ZN(G63) );
NOR3_X1 U785 ( .A1(n989), .A2(n1078), .A3(n1079), .ZN(n1077) );
NOR3_X1 U786 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
AND2_X1 U787 ( .A1(n1080), .A2(n1082), .ZN(n1078) );
NAND3_X1 U788 ( .A1(KEYINPUT60), .A2(G478), .A3(n1083), .ZN(n1082) );
XOR2_X1 U789 ( .A(n1076), .B(KEYINPUT16), .Z(n1083) );
INV_X1 U790 ( .A(n988), .ZN(n989) );
NOR2_X1 U791 ( .A1(n1070), .A2(n1084), .ZN(G60) );
XOR2_X1 U792 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U793 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
INV_X1 U794 ( .A(G475), .ZN(n1087) );
XNOR2_X1 U795 ( .A(G104), .B(n1089), .ZN(G6) );
NOR2_X1 U796 ( .A1(n1070), .A2(n1090), .ZN(G57) );
XOR2_X1 U797 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U798 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U799 ( .A(n1095), .B(n1096), .Z(n1091) );
XOR2_X1 U800 ( .A(KEYINPUT44), .B(n1097), .Z(n1096) );
NOR2_X1 U801 ( .A1(n984), .A2(n1088), .ZN(n1097) );
INV_X1 U802 ( .A(G472), .ZN(n984) );
NOR2_X1 U803 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
XOR2_X1 U804 ( .A(n1100), .B(KEYINPUT10), .Z(n1099) );
NOR2_X1 U805 ( .A1(n1070), .A2(n1101), .ZN(G54) );
XOR2_X1 U806 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U807 ( .A1(n1104), .A2(n1088), .ZN(n1102) );
INV_X1 U808 ( .A(G469), .ZN(n1104) );
NOR2_X1 U809 ( .A1(n1070), .A2(n1105), .ZN(G51) );
XOR2_X1 U810 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U811 ( .A(n1042), .B(n1068), .Z(n1107) );
XOR2_X1 U812 ( .A(n1108), .B(n1109), .Z(n1106) );
NOR2_X1 U813 ( .A1(G125), .A2(KEYINPUT13), .ZN(n1109) );
XOR2_X1 U814 ( .A(n1110), .B(n1111), .Z(n1108) );
NOR2_X1 U815 ( .A1(n1112), .A2(n1088), .ZN(n1111) );
NAND2_X1 U816 ( .A1(G902), .A2(n1076), .ZN(n1088) );
NAND3_X1 U817 ( .A1(n1065), .A2(n970), .A3(n1113), .ZN(n1076) );
INV_X1 U818 ( .A(n1048), .ZN(n1113) );
NAND2_X1 U819 ( .A1(n1114), .A2(n1115), .ZN(n1048) );
AND4_X1 U820 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
NOR4_X1 U821 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1114) );
NOR2_X1 U822 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR3_X1 U823 ( .A1(n1126), .A2(n1016), .A3(n1127), .ZN(n1122) );
INV_X1 U824 ( .A(n1128), .ZN(n1121) );
INV_X1 U825 ( .A(n1129), .ZN(n1120) );
NAND3_X1 U826 ( .A1(n1004), .A2(n1007), .A3(n1130), .ZN(n970) );
AND4_X1 U827 ( .A1(n1131), .A2(n1089), .A3(n1132), .A4(n1133), .ZN(n1065) );
AND4_X1 U828 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
NAND2_X1 U829 ( .A1(n1138), .A2(n1139), .ZN(n1132) );
NAND2_X1 U830 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U831 ( .A1(KEYINPUT26), .A2(n1142), .ZN(n1141) );
NAND2_X1 U832 ( .A1(n1143), .A2(n1006), .ZN(n1140) );
XOR2_X1 U833 ( .A(n1010), .B(KEYINPUT58), .Z(n1143) );
NAND3_X1 U834 ( .A1(n1130), .A2(n1004), .A3(n1006), .ZN(n1089) );
NAND3_X1 U835 ( .A1(n1001), .A2(n1142), .A3(n1144), .ZN(n1131) );
NOR3_X1 U836 ( .A1(n1145), .A2(KEYINPUT26), .A3(n1146), .ZN(n1144) );
NOR2_X1 U837 ( .A1(n975), .A2(G952), .ZN(n1070) );
XNOR2_X1 U838 ( .A(G146), .B(n1118), .ZN(G48) );
NAND3_X1 U839 ( .A1(n1147), .A2(n1146), .A3(n1006), .ZN(n1118) );
XOR2_X1 U840 ( .A(n1148), .B(n1128), .Z(G45) );
NAND4_X1 U841 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1128) );
NOR2_X1 U842 ( .A1(n992), .A2(n1016), .ZN(n1151) );
NAND2_X1 U843 ( .A1(n1153), .A2(n1154), .ZN(G42) );
OR2_X1 U844 ( .A1(n1129), .A2(G140), .ZN(n1154) );
XOR2_X1 U845 ( .A(n1155), .B(KEYINPUT19), .Z(n1153) );
NAND2_X1 U846 ( .A1(G140), .A2(n1129), .ZN(n1155) );
NAND2_X1 U847 ( .A1(n1156), .A2(n1157), .ZN(n1129) );
XOR2_X1 U848 ( .A(n1045), .B(n1117), .Z(G39) );
NAND3_X1 U849 ( .A1(n1147), .A2(n991), .A3(n1008), .ZN(n1117) );
INV_X1 U850 ( .A(G137), .ZN(n1045) );
XNOR2_X1 U851 ( .A(G134), .B(n1116), .ZN(G36) );
NAND3_X1 U852 ( .A1(n1142), .A2(n1149), .A3(n991), .ZN(n1116) );
XOR2_X1 U853 ( .A(n1046), .B(n1119), .Z(G33) );
NAND2_X1 U854 ( .A1(n1157), .A2(n1150), .ZN(n1119) );
AND3_X1 U855 ( .A1(n991), .A2(n1149), .A3(n1006), .ZN(n1157) );
NOR2_X1 U856 ( .A1(n1158), .A2(n1018), .ZN(n991) );
INV_X1 U857 ( .A(n1019), .ZN(n1158) );
XNOR2_X1 U858 ( .A(G128), .B(n1159), .ZN(G30) );
NAND3_X1 U859 ( .A1(n1147), .A2(n1007), .A3(n1160), .ZN(n1159) );
XOR2_X1 U860 ( .A(n1016), .B(KEYINPUT23), .Z(n1160) );
INV_X1 U861 ( .A(n1127), .ZN(n1007) );
INV_X1 U862 ( .A(n1126), .ZN(n1147) );
NAND3_X1 U863 ( .A1(n1149), .A2(n1161), .A3(n1162), .ZN(n1126) );
NOR2_X1 U864 ( .A1(n1023), .A2(n1124), .ZN(n1149) );
XOR2_X1 U865 ( .A(n1163), .B(n1137), .Z(G3) );
NAND3_X1 U866 ( .A1(n1150), .A2(n1130), .A3(n1008), .ZN(n1137) );
XOR2_X1 U867 ( .A(n1164), .B(n1165), .Z(G27) );
NOR2_X1 U868 ( .A1(KEYINPUT56), .A2(n1166), .ZN(n1165) );
NOR2_X1 U869 ( .A1(n1167), .A2(n1125), .ZN(n1164) );
NAND4_X1 U870 ( .A1(n1001), .A2(n1156), .A3(n1006), .A4(n1146), .ZN(n1125) );
INV_X1 U871 ( .A(n1168), .ZN(n1001) );
XNOR2_X1 U872 ( .A(n1124), .B(KEYINPUT29), .ZN(n1167) );
AND2_X1 U873 ( .A1(n1025), .A2(n1169), .ZN(n1124) );
NAND3_X1 U874 ( .A1(G902), .A2(n1170), .A3(n1036), .ZN(n1169) );
NOR2_X1 U875 ( .A1(n975), .A2(G900), .ZN(n1036) );
XOR2_X1 U876 ( .A(n1171), .B(n1136), .Z(G24) );
NAND4_X1 U877 ( .A1(n1138), .A2(n1004), .A3(n1152), .A4(n1172), .ZN(n1136) );
NOR2_X1 U878 ( .A1(n1173), .A2(n1161), .ZN(n1004) );
XNOR2_X1 U879 ( .A(G119), .B(n1135), .ZN(G21) );
NAND4_X1 U880 ( .A1(n1138), .A2(n1008), .A3(n1162), .A4(n1161), .ZN(n1135) );
INV_X1 U881 ( .A(n1174), .ZN(n1161) );
XOR2_X1 U882 ( .A(n1175), .B(G116), .Z(G18) );
NAND2_X1 U883 ( .A1(KEYINPUT18), .A2(n1176), .ZN(n1175) );
NAND3_X1 U884 ( .A1(n1177), .A2(n1178), .A3(n1142), .ZN(n1176) );
NOR2_X1 U885 ( .A1(n1010), .A2(n1127), .ZN(n1142) );
NAND2_X1 U886 ( .A1(n1152), .A2(n992), .ZN(n1127) );
INV_X1 U887 ( .A(n1150), .ZN(n1010) );
OR2_X1 U888 ( .A1(n1138), .A2(KEYINPUT22), .ZN(n1178) );
NAND2_X1 U889 ( .A1(KEYINPUT22), .A2(n1179), .ZN(n1177) );
NAND3_X1 U890 ( .A1(n1180), .A2(n1168), .A3(n1146), .ZN(n1179) );
XOR2_X1 U891 ( .A(n1181), .B(n1182), .Z(G15) );
NAND3_X1 U892 ( .A1(n1006), .A2(n1150), .A3(n1138), .ZN(n1182) );
NOR3_X1 U893 ( .A1(n1016), .A2(n1145), .A3(n1168), .ZN(n1138) );
NAND2_X1 U894 ( .A1(n986), .A2(n977), .ZN(n1168) );
INV_X1 U895 ( .A(n1024), .ZN(n986) );
NOR2_X1 U896 ( .A1(n1173), .A2(n1174), .ZN(n1150) );
NOR2_X1 U897 ( .A1(n992), .A2(n1152), .ZN(n1006) );
XNOR2_X1 U898 ( .A(G110), .B(n1134), .ZN(G12) );
NAND3_X1 U899 ( .A1(n1008), .A2(n1130), .A3(n1156), .ZN(n1134) );
INV_X1 U900 ( .A(n1011), .ZN(n1156) );
NAND2_X1 U901 ( .A1(n1162), .A2(n1174), .ZN(n1011) );
XNOR2_X1 U902 ( .A(n1183), .B(n985), .ZN(n1174) );
NAND2_X1 U903 ( .A1(n1184), .A2(n1081), .ZN(n985) );
XOR2_X1 U904 ( .A(n1185), .B(n1093), .Z(n1184) );
XOR2_X1 U905 ( .A(n1186), .B(n1163), .Z(n1093) );
NAND2_X1 U906 ( .A1(n1187), .A2(G210), .ZN(n1186) );
NAND2_X1 U907 ( .A1(KEYINPUT54), .A2(n1188), .ZN(n1185) );
XNOR2_X1 U908 ( .A(n1189), .B(n1094), .ZN(n1188) );
XNOR2_X1 U909 ( .A(n1190), .B(n1191), .ZN(n1094) );
NOR2_X1 U910 ( .A1(G119), .A2(KEYINPUT39), .ZN(n1191) );
XOR2_X1 U911 ( .A(n1181), .B(G116), .Z(n1190) );
INV_X1 U912 ( .A(G113), .ZN(n1181) );
NAND2_X1 U913 ( .A1(KEYINPUT11), .A2(G472), .ZN(n1183) );
XOR2_X1 U914 ( .A(n1173), .B(KEYINPUT40), .Z(n1162) );
NAND2_X1 U915 ( .A1(n1192), .A2(n1193), .ZN(n1173) );
NAND2_X1 U916 ( .A1(n1194), .A2(n995), .ZN(n1193) );
XOR2_X1 U917 ( .A(KEYINPUT63), .B(n1195), .Z(n1192) );
NOR2_X1 U918 ( .A1(n995), .A2(n1194), .ZN(n1195) );
XNOR2_X1 U919 ( .A(KEYINPUT31), .B(n993), .ZN(n1194) );
NAND2_X1 U920 ( .A1(n1196), .A2(n1073), .ZN(n993) );
XNOR2_X1 U921 ( .A(n1197), .B(n1198), .ZN(n1073) );
XOR2_X1 U922 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U923 ( .A(G119), .B(n1201), .Z(n1200) );
AND3_X1 U924 ( .A1(G221), .A2(n975), .A3(G234), .ZN(n1201) );
XOR2_X1 U925 ( .A(KEYINPUT51), .B(G137), .Z(n1199) );
XOR2_X1 U926 ( .A(n1202), .B(n1203), .Z(n1197) );
XNOR2_X1 U927 ( .A(n1041), .B(n1204), .ZN(n1202) );
XNOR2_X1 U928 ( .A(n1166), .B(n1205), .ZN(n1041) );
XOR2_X1 U929 ( .A(KEYINPUT46), .B(G902), .Z(n1196) );
NAND2_X1 U930 ( .A1(G217), .A2(n1206), .ZN(n995) );
NOR3_X1 U931 ( .A1(n1016), .A2(n1145), .A3(n1023), .ZN(n1130) );
NAND2_X1 U932 ( .A1(n1024), .A2(n977), .ZN(n1023) );
NAND2_X1 U933 ( .A1(G221), .A2(n1206), .ZN(n977) );
NAND2_X1 U934 ( .A1(G234), .A2(n1081), .ZN(n1206) );
XNOR2_X1 U935 ( .A(n1207), .B(G469), .ZN(n1024) );
OR2_X1 U936 ( .A1(n1103), .A2(G902), .ZN(n1207) );
XNOR2_X1 U937 ( .A(n1208), .B(n1209), .ZN(n1103) );
XOR2_X1 U938 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U939 ( .A(n1189), .B(n1212), .Z(n1211) );
NOR2_X1 U940 ( .A1(G953), .A2(n1051), .ZN(n1212) );
INV_X1 U941 ( .A(G227), .ZN(n1051) );
NAND2_X1 U942 ( .A1(n1213), .A2(n1100), .ZN(n1189) );
NAND2_X1 U943 ( .A1(n1214), .A2(n1215), .ZN(n1100) );
INV_X1 U944 ( .A(n1098), .ZN(n1213) );
NOR2_X1 U945 ( .A1(n1215), .A2(n1214), .ZN(n1098) );
XNOR2_X1 U946 ( .A(n1216), .B(n1217), .ZN(n1215) );
XOR2_X1 U947 ( .A(G137), .B(G134), .Z(n1217) );
NAND2_X1 U948 ( .A1(KEYINPUT43), .A2(n1046), .ZN(n1216) );
INV_X1 U949 ( .A(G131), .ZN(n1046) );
XNOR2_X1 U950 ( .A(KEYINPUT25), .B(G107), .ZN(n1210) );
XOR2_X1 U951 ( .A(n1218), .B(n1203), .Z(n1208) );
XOR2_X1 U952 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND2_X1 U953 ( .A1(KEYINPUT24), .A2(n1163), .ZN(n1219) );
INV_X1 U954 ( .A(G101), .ZN(n1163) );
INV_X1 U955 ( .A(n1180), .ZN(n1145) );
NAND2_X1 U956 ( .A1(n1025), .A2(n1221), .ZN(n1180) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1170), .A4(n1222), .ZN(n1221) );
INV_X1 U958 ( .A(G898), .ZN(n1222) );
NAND3_X1 U959 ( .A1(n1170), .A2(n975), .A3(G952), .ZN(n1025) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1170) );
INV_X1 U961 ( .A(n1146), .ZN(n1016) );
NOR2_X1 U962 ( .A1(n1019), .A2(n1018), .ZN(n1146) );
AND2_X1 U963 ( .A1(G214), .A2(n1223), .ZN(n1018) );
XNOR2_X1 U964 ( .A(n1224), .B(n1112), .ZN(n1019) );
NAND2_X1 U965 ( .A1(G210), .A2(n1223), .ZN(n1112) );
NAND2_X1 U966 ( .A1(n1081), .A2(n1225), .ZN(n1223) );
INV_X1 U967 ( .A(G237), .ZN(n1225) );
NAND2_X1 U968 ( .A1(n1226), .A2(n1081), .ZN(n1224) );
XOR2_X1 U969 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U970 ( .A(n1229), .B(n1230), .ZN(n1228) );
NOR2_X1 U971 ( .A1(KEYINPUT30), .A2(n1068), .ZN(n1230) );
XNOR2_X1 U972 ( .A(n1231), .B(n1232), .ZN(n1068) );
XOR2_X1 U973 ( .A(n1233), .B(n1203), .Z(n1232) );
XOR2_X1 U974 ( .A(G110), .B(KEYINPUT57), .Z(n1203) );
XOR2_X1 U975 ( .A(n1234), .B(n1235), .Z(n1231) );
XOR2_X1 U976 ( .A(G101), .B(n1236), .Z(n1235) );
NOR2_X1 U977 ( .A1(KEYINPUT0), .A2(n1237), .ZN(n1236) );
XOR2_X1 U978 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U979 ( .A(G119), .B(G116), .Z(n1239) );
XNOR2_X1 U980 ( .A(KEYINPUT50), .B(KEYINPUT2), .ZN(n1238) );
NAND2_X1 U981 ( .A1(KEYINPUT45), .A2(n1240), .ZN(n1234) );
XOR2_X1 U982 ( .A(G107), .B(n1241), .Z(n1240) );
NOR2_X1 U983 ( .A1(KEYINPUT38), .A2(n1242), .ZN(n1241) );
XNOR2_X1 U984 ( .A(G104), .B(n1243), .ZN(n1242) );
XOR2_X1 U985 ( .A(KEYINPUT25), .B(KEYINPUT14), .Z(n1243) );
NAND2_X1 U986 ( .A1(n1244), .A2(n1245), .ZN(n1229) );
NAND2_X1 U987 ( .A1(KEYINPUT61), .A2(n1246), .ZN(n1245) );
NAND2_X1 U988 ( .A1(KEYINPUT49), .A2(n1247), .ZN(n1244) );
INV_X1 U989 ( .A(n1246), .ZN(n1247) );
XOR2_X1 U990 ( .A(n1248), .B(n1042), .Z(n1246) );
INV_X1 U991 ( .A(n1214), .ZN(n1042) );
XOR2_X1 U992 ( .A(n1148), .B(n1204), .Z(n1214) );
XOR2_X1 U993 ( .A(G146), .B(G128), .Z(n1204) );
INV_X1 U994 ( .A(G143), .ZN(n1148) );
XOR2_X1 U995 ( .A(n1166), .B(KEYINPUT48), .Z(n1248) );
XNOR2_X1 U996 ( .A(KEYINPUT1), .B(n1110), .ZN(n1227) );
NAND2_X1 U997 ( .A1(G224), .A2(n975), .ZN(n1110) );
NOR2_X1 U998 ( .A1(n1172), .A2(n1152), .ZN(n1008) );
XOR2_X1 U999 ( .A(n988), .B(n1249), .Z(n1152) );
NOR2_X1 U1000 ( .A1(G478), .A2(KEYINPUT21), .ZN(n1249) );
NAND2_X1 U1001 ( .A1(n1081), .A2(n1080), .ZN(n988) );
NAND2_X1 U1002 ( .A1(n1250), .A2(n1251), .ZN(n1080) );
NAND4_X1 U1003 ( .A1(n1252), .A2(G217), .A3(G234), .A4(n975), .ZN(n1251) );
XOR2_X1 U1004 ( .A(n1253), .B(KEYINPUT20), .Z(n1252) );
XOR2_X1 U1005 ( .A(n1254), .B(KEYINPUT37), .Z(n1250) );
NAND2_X1 U1006 ( .A1(n1253), .A2(n1255), .ZN(n1254) );
NAND3_X1 U1007 ( .A1(G234), .A2(n975), .A3(G217), .ZN(n1255) );
INV_X1 U1008 ( .A(G953), .ZN(n975) );
XOR2_X1 U1009 ( .A(n1256), .B(n1257), .Z(n1253) );
XOR2_X1 U1010 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U1011 ( .A1(KEYINPUT59), .A2(G107), .ZN(n1259) );
NAND2_X1 U1012 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NAND2_X1 U1013 ( .A1(G134), .A2(n1262), .ZN(n1261) );
XOR2_X1 U1014 ( .A(KEYINPUT34), .B(n1263), .Z(n1260) );
NOR2_X1 U1015 ( .A1(G134), .A2(n1262), .ZN(n1263) );
XOR2_X1 U1016 ( .A(G143), .B(G128), .Z(n1262) );
XOR2_X1 U1017 ( .A(n1264), .B(G116), .Z(n1256) );
NAND2_X1 U1018 ( .A1(KEYINPUT12), .A2(n1171), .ZN(n1264) );
INV_X1 U1019 ( .A(G122), .ZN(n1171) );
INV_X1 U1020 ( .A(G902), .ZN(n1081) );
INV_X1 U1021 ( .A(n992), .ZN(n1172) );
XOR2_X1 U1022 ( .A(n1265), .B(G475), .Z(n992) );
OR2_X1 U1023 ( .A1(n1086), .A2(G902), .ZN(n1265) );
XNOR2_X1 U1024 ( .A(n1266), .B(n1267), .ZN(n1086) );
XOR2_X1 U1025 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U1026 ( .A(G143), .B(G131), .Z(n1269) );
XOR2_X1 U1027 ( .A(KEYINPUT9), .B(G146), .Z(n1268) );
XOR2_X1 U1028 ( .A(n1270), .B(n1271), .Z(n1266) );
XOR2_X1 U1029 ( .A(n1272), .B(n1273), .Z(n1271) );
NAND2_X1 U1030 ( .A1(n1187), .A2(G214), .ZN(n1273) );
NOR2_X1 U1031 ( .A1(G953), .A2(G237), .ZN(n1187) );
NAND2_X1 U1032 ( .A1(KEYINPUT53), .A2(n1166), .ZN(n1272) );
INV_X1 U1033 ( .A(G125), .ZN(n1166) );
XNOR2_X1 U1034 ( .A(n1220), .B(n1233), .ZN(n1270) );
XOR2_X1 U1035 ( .A(G113), .B(G122), .Z(n1233) );
XOR2_X1 U1036 ( .A(G104), .B(n1205), .Z(n1220) );
XOR2_X1 U1037 ( .A(G140), .B(KEYINPUT17), .Z(n1205) );
endmodule


