//Key = 1101101101111110010111100001101101011011101111000110111000001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U729 ( .A(n1014), .B(n1015), .ZN(G9) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U731 ( .A1(G953), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1017) );
NOR2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U738 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U739 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U740 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1035) );
NOR2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U743 ( .A1(n1041), .A2(n1044), .A3(n1034), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U745 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR4_X1 U746 ( .A1(n1049), .A2(n1034), .A3(n1041), .A4(n1030), .ZN(n1023) );
NOR2_X1 U747 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR3_X1 U748 ( .A1(n1018), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U749 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1018) );
NOR4_X1 U750 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
INV_X1 U751 ( .A(n1060), .ZN(n1059) );
AND2_X1 U752 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
NOR2_X1 U753 ( .A1(n1030), .A2(n1063), .ZN(n1054) );
XNOR2_X1 U754 ( .A(G472), .B(n1064), .ZN(n1063) );
INV_X1 U755 ( .A(n1065), .ZN(n1030) );
XOR2_X1 U756 ( .A(n1066), .B(n1067), .Z(G72) );
XOR2_X1 U757 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U758 ( .A1(G953), .A2(n1070), .ZN(n1069) );
NAND2_X1 U759 ( .A1(G900), .A2(G227), .ZN(n1070) );
NAND2_X1 U760 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NAND2_X1 U761 ( .A1(G953), .A2(n1073), .ZN(n1072) );
XOR2_X1 U762 ( .A(n1074), .B(n1075), .Z(n1071) );
XNOR2_X1 U763 ( .A(n1076), .B(G125), .ZN(n1075) );
NAND2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
NAND2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U766 ( .A(KEYINPUT14), .B(n1081), .Z(n1077) );
NOR2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1081) );
XNOR2_X1 U768 ( .A(n1082), .B(n1083), .ZN(n1080) );
NAND2_X1 U769 ( .A1(KEYINPUT36), .A2(n1084), .ZN(n1082) );
NOR2_X1 U770 ( .A1(n1085), .A2(G953), .ZN(n1066) );
XOR2_X1 U771 ( .A(n1086), .B(n1087), .Z(G69) );
NOR2_X1 U772 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NAND2_X1 U774 ( .A1(n1092), .A2(KEYINPUT35), .ZN(n1086) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U776 ( .A1(n1095), .A2(G953), .ZN(n1094) );
NOR3_X1 U777 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
XOR2_X1 U778 ( .A(n1099), .B(KEYINPUT38), .Z(n1098) );
NAND3_X1 U779 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1093) );
XOR2_X1 U780 ( .A(n1103), .B(KEYINPUT58), .Z(n1102) );
NAND2_X1 U781 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
OR2_X1 U782 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
XOR2_X1 U783 ( .A(n1106), .B(n1107), .Z(n1104) );
NAND2_X1 U784 ( .A1(G953), .A2(n1091), .ZN(n1100) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U786 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U787 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U788 ( .A1(n1061), .A2(n1114), .ZN(n1112) );
XOR2_X1 U789 ( .A(KEYINPUT25), .B(KEYINPUT18), .Z(n1110) );
NOR2_X1 U790 ( .A1(n1115), .A2(n1116), .ZN(G63) );
XOR2_X1 U791 ( .A(KEYINPUT8), .B(n1108), .Z(n1116) );
XNOR2_X1 U792 ( .A(n1117), .B(n1118), .ZN(n1115) );
NOR2_X1 U793 ( .A1(n1119), .A2(n1114), .ZN(n1118) );
INV_X1 U794 ( .A(G478), .ZN(n1119) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1120), .ZN(G60) );
XNOR2_X1 U796 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U797 ( .A1(n1123), .A2(n1114), .ZN(n1122) );
XNOR2_X1 U798 ( .A(G104), .B(n1124), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1108), .A2(n1125), .ZN(G57) );
XOR2_X1 U800 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U801 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U802 ( .A(n1130), .B(n1131), .Z(n1126) );
NOR2_X1 U803 ( .A1(n1132), .A2(n1114), .ZN(n1130) );
NOR2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(G54) );
XOR2_X1 U805 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U806 ( .A1(n1137), .A2(n1114), .ZN(n1136) );
XNOR2_X1 U807 ( .A(G469), .B(KEYINPUT32), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
XOR2_X1 U809 ( .A(n1140), .B(KEYINPUT1), .Z(n1139) );
NAND2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1142), .A2(n1141), .ZN(n1138) );
XNOR2_X1 U812 ( .A(n1143), .B(n1144), .ZN(n1141) );
XNOR2_X1 U813 ( .A(n1145), .B(n1129), .ZN(n1142) );
XNOR2_X1 U814 ( .A(n1079), .B(n1146), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1147), .B(KEYINPUT57), .Z(n1145) );
XNOR2_X1 U816 ( .A(n1108), .B(KEYINPUT53), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1108), .A2(n1148), .ZN(G51) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U819 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1114), .ZN(n1151) );
NAND2_X1 U821 ( .A1(G902), .A2(n1020), .ZN(n1114) );
NAND4_X1 U822 ( .A1(n1085), .A2(n1154), .A3(n1155), .A4(n1099), .ZN(n1020) );
XOR2_X1 U823 ( .A(KEYINPUT4), .B(n1097), .Z(n1155) );
INV_X1 U824 ( .A(n1096), .ZN(n1154) );
NAND4_X1 U825 ( .A1(n1156), .A2(n1157), .A3(n1124), .A4(n1158), .ZN(n1096) );
NOR3_X1 U826 ( .A1(n1159), .A2(n1015), .A3(n1160), .ZN(n1158) );
AND3_X1 U827 ( .A1(n1161), .A2(n1050), .A3(n1162), .ZN(n1015) );
NAND3_X1 U828 ( .A1(n1162), .A2(n1161), .A3(n1051), .ZN(n1124) );
AND4_X1 U829 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1085) );
NOR4_X1 U830 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U831 ( .A(n1171), .ZN(n1169) );
NOR3_X1 U832 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1168) );
XOR2_X1 U833 ( .A(KEYINPUT42), .B(n1051), .Z(n1172) );
NOR4_X1 U834 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1165) );
AND4_X1 U835 ( .A1(KEYINPUT37), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1178) );
NOR2_X1 U836 ( .A1(KEYINPUT37), .A2(n1182), .ZN(n1177) );
NOR4_X1 U837 ( .A1(n1183), .A2(n1184), .A3(n1053), .A4(n1185), .ZN(n1176) );
AND2_X1 U838 ( .A1(n1183), .A2(n1186), .ZN(n1175) );
INV_X1 U839 ( .A(KEYINPUT41), .ZN(n1183) );
XNOR2_X1 U840 ( .A(KEYINPUT63), .B(KEYINPUT44), .ZN(n1149) );
NOR2_X1 U841 ( .A1(n1089), .A2(G952), .ZN(n1108) );
XNOR2_X1 U842 ( .A(G146), .B(n1163), .ZN(G48) );
NAND2_X1 U843 ( .A1(n1187), .A2(n1051), .ZN(n1163) );
XNOR2_X1 U844 ( .A(G143), .B(n1182), .ZN(G45) );
NAND3_X1 U845 ( .A1(n1043), .A2(n1181), .A3(n1179), .ZN(n1182) );
INV_X1 U846 ( .A(n1185), .ZN(n1181) );
XNOR2_X1 U847 ( .A(G140), .B(n1188), .ZN(G42) );
NAND2_X1 U848 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U849 ( .A(n1167), .B(n1191), .Z(G39) );
NOR2_X1 U850 ( .A1(KEYINPUT2), .A2(n1192), .ZN(n1191) );
AND2_X1 U851 ( .A1(n1193), .A2(n1190), .ZN(n1167) );
NAND2_X1 U852 ( .A1(n1194), .A2(n1195), .ZN(G36) );
NAND2_X1 U853 ( .A1(n1186), .A2(n1196), .ZN(n1195) );
XOR2_X1 U854 ( .A(KEYINPUT39), .B(n1197), .Z(n1194) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1196), .ZN(n1197) );
XOR2_X1 U856 ( .A(KEYINPUT3), .B(G134), .Z(n1196) );
NOR2_X1 U857 ( .A1(n1184), .A2(n1173), .ZN(n1186) );
INV_X1 U858 ( .A(n1190), .ZN(n1173) );
XNOR2_X1 U859 ( .A(G131), .B(n1164), .ZN(G33) );
NAND3_X1 U860 ( .A1(n1190), .A2(n1051), .A3(n1043), .ZN(n1164) );
NOR2_X1 U861 ( .A1(n1185), .A2(n1041), .ZN(n1190) );
INV_X1 U862 ( .A(n1053), .ZN(n1041) );
NOR2_X1 U863 ( .A1(n1037), .A2(n1198), .ZN(n1053) );
NOR2_X1 U864 ( .A1(n1039), .A2(n1038), .ZN(n1198) );
INV_X1 U865 ( .A(G214), .ZN(n1039) );
XOR2_X1 U866 ( .A(G128), .B(n1170), .Z(G30) );
AND2_X1 U867 ( .A1(n1187), .A2(n1050), .ZN(n1170) );
NOR4_X1 U868 ( .A1(n1199), .A2(n1185), .A3(n1200), .A4(n1201), .ZN(n1187) );
NAND2_X1 U869 ( .A1(n1046), .A2(n1202), .ZN(n1185) );
XOR2_X1 U870 ( .A(n1203), .B(n1097), .Z(G3) );
AND3_X1 U871 ( .A1(n1162), .A2(n1204), .A3(n1043), .ZN(n1097) );
NAND2_X1 U872 ( .A1(KEYINPUT0), .A2(n1205), .ZN(n1203) );
INV_X1 U873 ( .A(G101), .ZN(n1205) );
NAND2_X1 U874 ( .A1(n1206), .A2(n1207), .ZN(G27) );
NAND2_X1 U875 ( .A1(G125), .A2(n1171), .ZN(n1207) );
XOR2_X1 U876 ( .A(KEYINPUT10), .B(n1208), .Z(n1206) );
NOR2_X1 U877 ( .A1(G125), .A2(n1171), .ZN(n1208) );
NAND4_X1 U878 ( .A1(n1189), .A2(n1065), .A3(n1036), .A4(n1202), .ZN(n1171) );
NAND2_X1 U879 ( .A1(n1022), .A2(n1209), .ZN(n1202) );
NAND4_X1 U880 ( .A1(G953), .A2(G902), .A3(n1210), .A4(n1073), .ZN(n1209) );
INV_X1 U881 ( .A(G900), .ZN(n1073) );
AND2_X1 U882 ( .A1(n1042), .A2(n1051), .ZN(n1189) );
XOR2_X1 U883 ( .A(G122), .B(n1159), .Z(G24) );
AND3_X1 U884 ( .A1(n1179), .A2(n1161), .A3(n1211), .ZN(n1159) );
INV_X1 U885 ( .A(n1034), .ZN(n1161) );
NAND2_X1 U886 ( .A1(n1201), .A2(n1199), .ZN(n1034) );
AND3_X1 U887 ( .A1(n1036), .A2(n1212), .A3(n1213), .ZN(n1179) );
NAND2_X1 U888 ( .A1(n1214), .A2(n1215), .ZN(G21) );
OR2_X1 U889 ( .A1(n1216), .A2(G119), .ZN(n1215) );
NAND2_X1 U890 ( .A1(n1217), .A2(G119), .ZN(n1214) );
NAND2_X1 U891 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
OR2_X1 U892 ( .A1(n1156), .A2(KEYINPUT28), .ZN(n1219) );
NAND2_X1 U893 ( .A1(KEYINPUT28), .A2(n1216), .ZN(n1218) );
NAND2_X1 U894 ( .A1(KEYINPUT30), .A2(n1220), .ZN(n1216) );
INV_X1 U895 ( .A(n1156), .ZN(n1220) );
NAND3_X1 U896 ( .A1(n1193), .A2(n1036), .A3(n1211), .ZN(n1156) );
NOR3_X1 U897 ( .A1(n1026), .A2(n1201), .A3(n1199), .ZN(n1193) );
INV_X1 U898 ( .A(n1204), .ZN(n1026) );
XNOR2_X1 U899 ( .A(G116), .B(n1221), .ZN(G18) );
NOR2_X1 U900 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U901 ( .A1(n1224), .A2(n1099), .ZN(n1223) );
NAND2_X1 U902 ( .A1(n1225), .A2(n1036), .ZN(n1099) );
INV_X1 U903 ( .A(KEYINPUT50), .ZN(n1224) );
NOR3_X1 U904 ( .A1(KEYINPUT50), .A2(n1225), .A3(n1200), .ZN(n1222) );
NOR2_X1 U905 ( .A1(n1226), .A2(n1184), .ZN(n1225) );
NAND2_X1 U906 ( .A1(n1043), .A2(n1050), .ZN(n1184) );
AND2_X1 U907 ( .A1(n1227), .A2(n1228), .ZN(n1050) );
XOR2_X1 U908 ( .A(n1212), .B(KEYINPUT46), .Z(n1227) );
XNOR2_X1 U909 ( .A(G113), .B(n1157), .ZN(G15) );
NAND4_X1 U910 ( .A1(n1211), .A2(n1043), .A3(n1229), .A4(n1051), .ZN(n1157) );
INV_X1 U911 ( .A(n1180), .ZN(n1043) );
NAND2_X1 U912 ( .A1(n1230), .A2(n1201), .ZN(n1180) );
INV_X1 U913 ( .A(n1199), .ZN(n1230) );
INV_X1 U914 ( .A(n1226), .ZN(n1211) );
NAND2_X1 U915 ( .A1(n1065), .A2(n1231), .ZN(n1226) );
NOR2_X1 U916 ( .A1(n1048), .A2(n1232), .ZN(n1065) );
INV_X1 U917 ( .A(n1047), .ZN(n1232) );
XNOR2_X1 U918 ( .A(n1233), .B(n1160), .ZN(G12) );
AND3_X1 U919 ( .A1(n1162), .A2(n1204), .A3(n1042), .ZN(n1160) );
INV_X1 U920 ( .A(n1174), .ZN(n1042) );
NAND2_X1 U921 ( .A1(n1234), .A2(n1199), .ZN(n1174) );
XOR2_X1 U922 ( .A(n1235), .B(n1064), .Z(n1199) );
NAND2_X1 U923 ( .A1(n1236), .A2(n1237), .ZN(n1064) );
XOR2_X1 U924 ( .A(n1238), .B(n1131), .Z(n1236) );
XNOR2_X1 U925 ( .A(n1239), .B(n1240), .ZN(n1131) );
NAND2_X1 U926 ( .A1(n1241), .A2(G210), .ZN(n1239) );
NAND2_X1 U927 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
OR2_X1 U928 ( .A1(n1128), .A2(n1244), .ZN(n1243) );
XOR2_X1 U929 ( .A(n1245), .B(KEYINPUT16), .Z(n1242) );
NAND2_X1 U930 ( .A1(n1244), .A2(n1128), .ZN(n1245) );
XNOR2_X1 U931 ( .A(n1246), .B(n1247), .ZN(n1128) );
NOR2_X1 U932 ( .A1(KEYINPUT51), .A2(G116), .ZN(n1247) );
XNOR2_X1 U933 ( .A(G113), .B(G119), .ZN(n1246) );
XOR2_X1 U934 ( .A(n1248), .B(n1249), .Z(n1244) );
NOR2_X1 U935 ( .A1(KEYINPUT24), .A2(n1250), .ZN(n1249) );
INV_X1 U936 ( .A(n1146), .ZN(n1250) );
NAND2_X1 U937 ( .A1(KEYINPUT22), .A2(n1132), .ZN(n1235) );
INV_X1 U938 ( .A(G472), .ZN(n1132) );
XOR2_X1 U939 ( .A(KEYINPUT61), .B(n1201), .Z(n1234) );
NOR2_X1 U940 ( .A1(n1251), .A2(n1056), .ZN(n1201) );
NOR2_X1 U941 ( .A1(n1061), .A2(n1062), .ZN(n1056) );
AND2_X1 U942 ( .A1(n1252), .A2(n1062), .ZN(n1251) );
NOR2_X1 U943 ( .A1(n1113), .A2(G902), .ZN(n1062) );
XNOR2_X1 U944 ( .A(n1253), .B(n1254), .ZN(n1113) );
XOR2_X1 U945 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U946 ( .A(n1257), .B(n1258), .ZN(n1256) );
NAND2_X1 U947 ( .A1(KEYINPUT52), .A2(n1233), .ZN(n1258) );
NAND2_X1 U948 ( .A1(KEYINPUT19), .A2(n1259), .ZN(n1257) );
XNOR2_X1 U949 ( .A(n1260), .B(n1261), .ZN(n1259) );
XNOR2_X1 U950 ( .A(n1262), .B(n1263), .ZN(n1261) );
NAND2_X1 U951 ( .A1(KEYINPUT7), .A2(n1264), .ZN(n1262) );
NAND3_X1 U952 ( .A1(n1265), .A2(G221), .A3(KEYINPUT20), .ZN(n1255) );
XNOR2_X1 U953 ( .A(G119), .B(n1266), .ZN(n1253) );
XNOR2_X1 U954 ( .A(n1192), .B(G128), .ZN(n1266) );
XOR2_X1 U955 ( .A(n1061), .B(KEYINPUT34), .Z(n1252) );
NAND2_X1 U956 ( .A1(G217), .A2(n1267), .ZN(n1061) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1269), .ZN(n1204) );
OR3_X1 U958 ( .A1(n1212), .A2(n1213), .A3(KEYINPUT29), .ZN(n1269) );
INV_X1 U959 ( .A(n1228), .ZN(n1213) );
NAND2_X1 U960 ( .A1(KEYINPUT29), .A2(n1051), .ZN(n1268) );
NOR2_X1 U961 ( .A1(n1228), .A2(n1212), .ZN(n1051) );
NAND2_X1 U962 ( .A1(n1270), .A2(n1060), .ZN(n1212) );
NAND2_X1 U963 ( .A1(G478), .A2(n1271), .ZN(n1060) );
NAND2_X1 U964 ( .A1(n1117), .A2(n1237), .ZN(n1271) );
XNOR2_X1 U965 ( .A(n1057), .B(KEYINPUT26), .ZN(n1270) );
NOR3_X1 U966 ( .A1(G478), .A2(G902), .A3(n1272), .ZN(n1057) );
INV_X1 U967 ( .A(n1117), .ZN(n1272) );
XNOR2_X1 U968 ( .A(n1273), .B(n1274), .ZN(n1117) );
XNOR2_X1 U969 ( .A(n1014), .B(n1275), .ZN(n1274) );
XOR2_X1 U970 ( .A(G122), .B(G116), .Z(n1275) );
XOR2_X1 U971 ( .A(n1276), .B(n1277), .Z(n1273) );
AND2_X1 U972 ( .A1(G217), .A2(n1265), .ZN(n1277) );
AND2_X1 U973 ( .A1(G234), .A2(n1089), .ZN(n1265) );
NAND3_X1 U974 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1276) );
OR2_X1 U975 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U976 ( .A1(n1283), .A2(n1284), .ZN(n1279) );
INV_X1 U977 ( .A(KEYINPUT33), .ZN(n1284) );
NAND2_X1 U978 ( .A1(n1285), .A2(n1281), .ZN(n1283) );
XNOR2_X1 U979 ( .A(KEYINPUT9), .B(n1282), .ZN(n1285) );
NAND2_X1 U980 ( .A1(KEYINPUT33), .A2(n1286), .ZN(n1278) );
NAND2_X1 U981 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND3_X1 U982 ( .A1(KEYINPUT9), .A2(n1281), .A3(n1282), .ZN(n1288) );
XOR2_X1 U983 ( .A(n1084), .B(KEYINPUT48), .Z(n1281) );
OR2_X1 U984 ( .A1(n1282), .A2(KEYINPUT9), .ZN(n1287) );
XNOR2_X1 U985 ( .A(n1052), .B(KEYINPUT12), .ZN(n1228) );
XNOR2_X1 U986 ( .A(n1289), .B(n1123), .ZN(n1052) );
INV_X1 U987 ( .A(G475), .ZN(n1123) );
NAND2_X1 U988 ( .A1(n1121), .A2(n1237), .ZN(n1289) );
XNOR2_X1 U989 ( .A(n1290), .B(n1291), .ZN(n1121) );
XOR2_X1 U990 ( .A(n1260), .B(n1292), .Z(n1291) );
XOR2_X1 U991 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U992 ( .A1(KEYINPUT55), .A2(n1295), .ZN(n1294) );
XNOR2_X1 U993 ( .A(n1296), .B(n1297), .ZN(n1295) );
XOR2_X1 U994 ( .A(G122), .B(G113), .Z(n1297) );
NOR2_X1 U995 ( .A1(n1298), .A2(n1299), .ZN(n1293) );
XOR2_X1 U996 ( .A(n1300), .B(KEYINPUT31), .Z(n1299) );
NAND2_X1 U997 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U998 ( .A1(n1241), .A2(G214), .ZN(n1302) );
INV_X1 U999 ( .A(G143), .ZN(n1301) );
AND3_X1 U1000 ( .A1(n1241), .A2(G143), .A3(G214), .ZN(n1298) );
NOR2_X1 U1001 ( .A1(G953), .A2(G237), .ZN(n1241) );
XOR2_X1 U1002 ( .A(G140), .B(KEYINPUT40), .Z(n1260) );
XNOR2_X1 U1003 ( .A(G125), .B(n1303), .ZN(n1290) );
XNOR2_X1 U1004 ( .A(n1263), .B(G131), .ZN(n1303) );
INV_X1 U1005 ( .A(G146), .ZN(n1263) );
AND3_X1 U1006 ( .A1(n1229), .A2(n1231), .A3(n1046), .ZN(n1162) );
AND2_X1 U1007 ( .A1(n1304), .A2(n1048), .ZN(n1046) );
XNOR2_X1 U1008 ( .A(n1305), .B(G469), .ZN(n1048) );
NAND2_X1 U1009 ( .A1(n1306), .A2(n1237), .ZN(n1305) );
XOR2_X1 U1010 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1011 ( .A(n1248), .B(n1309), .ZN(n1308) );
XOR2_X1 U1012 ( .A(n1147), .B(n1310), .Z(n1309) );
NOR2_X1 U1013 ( .A1(KEYINPUT15), .A2(n1144), .ZN(n1310) );
XNOR2_X1 U1014 ( .A(n1233), .B(n1076), .ZN(n1144) );
INV_X1 U1015 ( .A(G140), .ZN(n1076) );
NAND2_X1 U1016 ( .A1(n1311), .A2(n1312), .ZN(n1147) );
NAND2_X1 U1017 ( .A1(n1313), .A2(n1240), .ZN(n1312) );
XOR2_X1 U1018 ( .A(n1314), .B(KEYINPUT47), .Z(n1311) );
OR2_X1 U1019 ( .A1(n1240), .A2(n1313), .ZN(n1314) );
XOR2_X1 U1020 ( .A(n1315), .B(n1296), .Z(n1313) );
INV_X1 U1021 ( .A(G104), .ZN(n1296) );
NAND2_X1 U1022 ( .A1(KEYINPUT60), .A2(n1014), .ZN(n1315) );
INV_X1 U1023 ( .A(n1079), .ZN(n1248) );
XOR2_X1 U1024 ( .A(n1316), .B(n1143), .Z(n1307) );
AND2_X1 U1025 ( .A1(G227), .A2(n1089), .ZN(n1143) );
XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n1317), .ZN(n1316) );
NOR2_X1 U1027 ( .A1(KEYINPUT5), .A2(n1146), .ZN(n1317) );
XNOR2_X1 U1028 ( .A(n1318), .B(n1083), .ZN(n1146) );
XNOR2_X1 U1029 ( .A(G131), .B(n1192), .ZN(n1083) );
INV_X1 U1030 ( .A(G137), .ZN(n1192) );
XNOR2_X1 U1031 ( .A(KEYINPUT45), .B(n1319), .ZN(n1318) );
NOR2_X1 U1032 ( .A1(KEYINPUT59), .A2(n1084), .ZN(n1319) );
XOR2_X1 U1033 ( .A(G134), .B(KEYINPUT54), .Z(n1084) );
XOR2_X1 U1034 ( .A(n1047), .B(KEYINPUT56), .Z(n1304) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1267), .ZN(n1047) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1320), .ZN(n1267) );
NAND2_X1 U1037 ( .A1(n1022), .A2(n1321), .ZN(n1231) );
NAND4_X1 U1038 ( .A1(G953), .A2(G902), .A3(n1210), .A4(n1091), .ZN(n1321) );
INV_X1 U1039 ( .A(G898), .ZN(n1091) );
NAND3_X1 U1040 ( .A1(n1210), .A2(n1089), .A3(G952), .ZN(n1022) );
INV_X1 U1041 ( .A(G953), .ZN(n1089) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1210) );
XNOR2_X1 U1043 ( .A(n1036), .B(KEYINPUT11), .ZN(n1229) );
INV_X1 U1044 ( .A(n1200), .ZN(n1036) );
NAND2_X1 U1045 ( .A1(n1037), .A2(n1322), .ZN(n1200) );
NAND2_X1 U1046 ( .A1(G214), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1047 ( .A(n1324), .B(n1153), .Z(n1037) );
NAND2_X1 U1048 ( .A1(G210), .A2(n1323), .ZN(n1153) );
INV_X1 U1049 ( .A(n1038), .ZN(n1323) );
NOR2_X1 U1050 ( .A1(n1325), .A2(G237), .ZN(n1038) );
INV_X1 U1051 ( .A(n1320), .ZN(n1325) );
XNOR2_X1 U1052 ( .A(n1237), .B(KEYINPUT27), .ZN(n1320) );
NAND2_X1 U1053 ( .A1(n1326), .A2(n1237), .ZN(n1324) );
INV_X1 U1054 ( .A(G902), .ZN(n1237) );
XOR2_X1 U1055 ( .A(KEYINPUT62), .B(n1152), .Z(n1326) );
XNOR2_X1 U1056 ( .A(n1327), .B(n1328), .ZN(n1152) );
XOR2_X1 U1057 ( .A(n1106), .B(n1329), .Z(n1328) );
XNOR2_X1 U1058 ( .A(n1105), .B(n1079), .ZN(n1329) );
XOR2_X1 U1059 ( .A(G146), .B(n1282), .Z(n1079) );
XNOR2_X1 U1060 ( .A(G128), .B(G143), .ZN(n1282) );
XNOR2_X1 U1061 ( .A(n1330), .B(n1233), .ZN(n1105) );
NAND2_X1 U1062 ( .A1(KEYINPUT43), .A2(G122), .ZN(n1330) );
NAND2_X1 U1063 ( .A1(n1331), .A2(n1332), .ZN(n1106) );
NAND2_X1 U1064 ( .A1(n1333), .A2(n1014), .ZN(n1332) );
INV_X1 U1065 ( .A(G107), .ZN(n1014) );
XNOR2_X1 U1066 ( .A(n1334), .B(KEYINPUT17), .ZN(n1333) );
NAND2_X1 U1067 ( .A1(n1335), .A2(G107), .ZN(n1331) );
XOR2_X1 U1068 ( .A(KEYINPUT13), .B(n1334), .Z(n1335) );
XOR2_X1 U1069 ( .A(G104), .B(n1240), .Z(n1334) );
XOR2_X1 U1070 ( .A(G101), .B(KEYINPUT6), .Z(n1240) );
XOR2_X1 U1071 ( .A(n1336), .B(n1337), .Z(n1327) );
XNOR2_X1 U1072 ( .A(n1264), .B(n1338), .ZN(n1337) );
NOR2_X1 U1073 ( .A1(G953), .A2(n1090), .ZN(n1338) );
INV_X1 U1074 ( .A(G224), .ZN(n1090) );
INV_X1 U1075 ( .A(G125), .ZN(n1264) );
NAND2_X1 U1076 ( .A1(KEYINPUT21), .A2(n1107), .ZN(n1336) );
XOR2_X1 U1077 ( .A(n1339), .B(n1340), .Z(n1107) );
NOR2_X1 U1078 ( .A1(KEYINPUT23), .A2(n1341), .ZN(n1340) );
INV_X1 U1079 ( .A(G119), .ZN(n1341) );
XNOR2_X1 U1080 ( .A(G113), .B(G116), .ZN(n1339) );
INV_X1 U1081 ( .A(G110), .ZN(n1233) );
endmodule


