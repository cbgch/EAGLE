//Key = 0101110000011110000110111011110011100110110101001111100100000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;

XNOR2_X1 U747 ( .A(G107), .B(n1033), .ZN(G9) );
NOR2_X1 U748 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U749 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U750 ( .A1(KEYINPUT49), .A2(n1039), .ZN(n1037) );
NOR4_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND3_X1 U752 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1040) );
NAND3_X1 U753 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1036) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND4_X1 U756 ( .A1(n1054), .A2(n1044), .A3(n1055), .A4(n1045), .ZN(n1053) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U761 ( .A(n1064), .ZN(n1060) );
NAND2_X1 U762 ( .A1(n1046), .A2(n1065), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
OR2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U765 ( .A1(n1046), .A2(n1070), .A3(n1058), .ZN(n1052) );
NAND2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1044), .ZN(n1072) );
OR2_X1 U768 ( .A1(n1045), .A2(n1054), .ZN(n1074) );
NAND3_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1045), .ZN(n1073) );
NAND2_X1 U770 ( .A1(KEYINPUT49), .A2(n1077), .ZN(n1075) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1054), .ZN(n1071) );
INV_X1 U772 ( .A(n1041), .ZN(n1050) );
NOR3_X1 U773 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1034) );
INV_X1 U774 ( .A(n1047), .ZN(n1079) );
NAND4_X1 U775 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1047) );
AND3_X1 U776 ( .A1(n1045), .A2(n1084), .A3(n1068), .ZN(n1083) );
NOR3_X1 U777 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1082) );
NOR2_X1 U778 ( .A1(G478), .A2(n1088), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
XOR2_X1 U780 ( .A(n1091), .B(KEYINPUT9), .Z(n1085) );
NAND3_X1 U781 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U783 ( .A1(KEYINPUT0), .A2(n1097), .ZN(n1093) );
NAND2_X1 U784 ( .A1(n1098), .A2(G472), .ZN(n1097) );
XNOR2_X1 U785 ( .A(n1095), .B(KEYINPUT60), .ZN(n1098) );
NAND2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1092) );
INV_X1 U787 ( .A(KEYINPUT0), .ZN(n1100) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
OR3_X1 U789 ( .A1(n1096), .A2(n1095), .A3(KEYINPUT60), .ZN(n1102) );
NAND2_X1 U790 ( .A1(KEYINPUT60), .A2(n1095), .ZN(n1101) );
NOR3_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1081) );
XNOR2_X1 U792 ( .A(n1106), .B(n1107), .ZN(n1105) );
XOR2_X1 U793 ( .A(KEYINPUT40), .B(G469), .Z(n1107) );
XOR2_X1 U794 ( .A(n1108), .B(KEYINPUT34), .Z(n1104) );
NAND2_X1 U795 ( .A1(G478), .A2(n1088), .ZN(n1108) );
NOR2_X1 U796 ( .A1(KEYINPUT27), .A2(n1109), .ZN(n1103) );
NOR3_X1 U797 ( .A1(n1063), .A2(n1110), .A3(n1111), .ZN(n1080) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U800 ( .A(n1109), .B(KEYINPUT23), .Z(n1114) );
INV_X1 U801 ( .A(n1116), .ZN(n1112) );
NOR3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1115), .ZN(n1110) );
INV_X1 U803 ( .A(KEYINPUT27), .ZN(n1115) );
INV_X1 U804 ( .A(n1109), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(G72) );
NOR3_X1 U806 ( .A1(n1048), .A2(KEYINPUT17), .A3(n1120), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1118) );
NOR2_X1 U809 ( .A1(n1125), .A2(KEYINPUT15), .ZN(n1124) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U813 ( .A(n1132), .B(n1133), .Z(n1128) );
XOR2_X1 U814 ( .A(KEYINPUT26), .B(G131), .Z(n1133) );
NAND2_X1 U815 ( .A1(KEYINPUT1), .A2(n1134), .ZN(n1132) );
NOR2_X1 U816 ( .A1(G900), .A2(n1135), .ZN(n1126) );
XOR2_X1 U817 ( .A(KEYINPUT63), .B(G953), .Z(n1135) );
NAND2_X1 U818 ( .A1(n1048), .A2(n1136), .ZN(n1123) );
NAND2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U820 ( .A(KEYINPUT18), .B(n1139), .Z(n1138) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(G69) );
NOR2_X1 U822 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U823 ( .A(n1144), .B(n1145), .ZN(n1143) );
XOR2_X1 U824 ( .A(n1146), .B(KEYINPUT30), .Z(n1144) );
NAND3_X1 U825 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1140) );
INV_X1 U826 ( .A(n1142), .ZN(n1149) );
OR2_X1 U827 ( .A1(n1048), .A2(G224), .ZN(n1148) );
NAND2_X1 U828 ( .A1(n1150), .A2(n1048), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XNOR2_X1 U831 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U832 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U833 ( .A1(n1153), .A2(n1159), .ZN(G63) );
NOR3_X1 U834 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1159) );
NOR4_X1 U835 ( .A1(n1163), .A2(n1158), .A3(KEYINPUT46), .A4(n1164), .ZN(n1162) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1161) );
INV_X1 U837 ( .A(n1163), .ZN(n1166) );
NOR3_X1 U838 ( .A1(n1164), .A2(KEYINPUT46), .A3(n1167), .ZN(n1165) );
INV_X1 U839 ( .A(n1038), .ZN(n1167) );
INV_X1 U840 ( .A(G478), .ZN(n1164) );
INV_X1 U841 ( .A(n1088), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1153), .A2(n1168), .ZN(G60) );
XOR2_X1 U843 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U844 ( .A(KEYINPUT3), .B(n1171), .Z(n1170) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1158), .ZN(n1171) );
XNOR2_X1 U846 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(G57) );
XOR2_X1 U848 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U849 ( .A(KEYINPUT5), .B(n1178), .Z(n1177) );
NOR2_X1 U850 ( .A1(KEYINPUT2), .A2(n1179), .ZN(n1178) );
XOR2_X1 U851 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U852 ( .A(KEYINPUT59), .B(n1182), .ZN(n1181) );
NOR2_X1 U853 ( .A1(KEYINPUT31), .A2(n1183), .ZN(n1182) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1176) );
NOR2_X1 U855 ( .A1(n1096), .A2(n1158), .ZN(n1185) );
INV_X1 U856 ( .A(G472), .ZN(n1096) );
XNOR2_X1 U857 ( .A(n1153), .B(KEYINPUT38), .ZN(n1174) );
NOR2_X1 U858 ( .A1(n1153), .A2(n1186), .ZN(G54) );
XOR2_X1 U859 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U860 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U861 ( .A(n1191), .B(n1192), .Z(n1190) );
XNOR2_X1 U862 ( .A(G140), .B(n1183), .ZN(n1192) );
XOR2_X1 U863 ( .A(KEYINPUT45), .B(KEYINPUT24), .Z(n1191) );
XOR2_X1 U864 ( .A(n1193), .B(n1194), .Z(n1189) );
XOR2_X1 U865 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U866 ( .A1(n1197), .A2(n1158), .ZN(n1196) );
NOR2_X1 U867 ( .A1(KEYINPUT21), .A2(n1198), .ZN(n1195) );
XNOR2_X1 U868 ( .A(n1199), .B(n1134), .ZN(n1193) );
NAND2_X1 U869 ( .A1(G227), .A2(n1048), .ZN(n1199) );
NOR2_X1 U870 ( .A1(n1153), .A2(n1200), .ZN(G51) );
XOR2_X1 U871 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U872 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U873 ( .A1(n1116), .A2(n1158), .ZN(n1204) );
NAND2_X1 U874 ( .A1(G902), .A2(n1038), .ZN(n1158) );
NAND4_X1 U875 ( .A1(n1205), .A2(n1139), .A3(n1151), .A4(n1137), .ZN(n1038) );
AND4_X1 U876 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1137) );
AND4_X1 U877 ( .A1(n1210), .A2(n1211), .A3(n1173), .A4(n1212), .ZN(n1151) );
AND4_X1 U878 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1033), .ZN(n1212) );
NAND3_X1 U879 ( .A1(n1046), .A2(n1216), .A3(n1217), .ZN(n1033) );
NAND3_X1 U880 ( .A1(n1046), .A2(n1216), .A3(n1077), .ZN(n1173) );
AND4_X1 U881 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1139) );
XOR2_X1 U882 ( .A(n1152), .B(KEYINPUT8), .Z(n1205) );
NAND2_X1 U883 ( .A1(n1222), .A2(n1223), .ZN(n1152) );
XOR2_X1 U884 ( .A(n1224), .B(KEYINPUT61), .Z(n1222) );
NOR2_X1 U885 ( .A1(n1048), .A2(G952), .ZN(n1153) );
XOR2_X1 U886 ( .A(n1225), .B(n1218), .Z(G48) );
NAND3_X1 U887 ( .A1(n1077), .A2(n1223), .A3(n1226), .ZN(n1218) );
XNOR2_X1 U888 ( .A(G143), .B(n1219), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1078), .A2(n1223), .A3(n1064), .A4(n1227), .ZN(n1219) );
AND3_X1 U890 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
XOR2_X1 U891 ( .A(n1231), .B(G140), .Z(G42) );
NAND2_X1 U892 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
OR2_X1 U893 ( .A1(n1220), .A2(KEYINPUT10), .ZN(n1233) );
NAND3_X1 U894 ( .A1(n1058), .A2(n1078), .A3(n1234), .ZN(n1220) );
NAND3_X1 U895 ( .A1(n1058), .A2(n1235), .A3(KEYINPUT10), .ZN(n1232) );
NAND2_X1 U896 ( .A1(n1234), .A2(n1078), .ZN(n1235) );
XOR2_X1 U897 ( .A(n1236), .B(n1221), .Z(G39) );
NAND3_X1 U898 ( .A1(n1058), .A2(n1054), .A3(n1226), .ZN(n1221) );
XNOR2_X1 U899 ( .A(n1206), .B(n1237), .ZN(G36) );
NOR2_X1 U900 ( .A1(KEYINPUT16), .A2(n1238), .ZN(n1237) );
NAND2_X1 U901 ( .A1(n1239), .A2(n1217), .ZN(n1206) );
NAND2_X1 U902 ( .A1(n1240), .A2(n1241), .ZN(G33) );
NAND2_X1 U903 ( .A1(G131), .A2(n1207), .ZN(n1241) );
XOR2_X1 U904 ( .A(KEYINPUT48), .B(n1242), .Z(n1240) );
NOR2_X1 U905 ( .A1(G131), .A2(n1207), .ZN(n1242) );
NAND2_X1 U906 ( .A1(n1239), .A2(n1077), .ZN(n1207) );
AND4_X1 U907 ( .A1(n1064), .A2(n1058), .A3(n1078), .A4(n1229), .ZN(n1239) );
INV_X1 U908 ( .A(n1043), .ZN(n1058) );
NAND2_X1 U909 ( .A1(n1243), .A2(n1068), .ZN(n1043) );
INV_X1 U910 ( .A(n1069), .ZN(n1243) );
XOR2_X1 U911 ( .A(G128), .B(n1244), .Z(G30) );
NOR2_X1 U912 ( .A1(KEYINPUT47), .A2(n1208), .ZN(n1244) );
NAND3_X1 U913 ( .A1(n1217), .A2(n1223), .A3(n1226), .ZN(n1208) );
AND4_X1 U914 ( .A1(n1245), .A2(n1078), .A3(n1063), .A4(n1229), .ZN(n1226) );
XNOR2_X1 U915 ( .A(G101), .B(n1210), .ZN(G3) );
NAND3_X1 U916 ( .A1(n1216), .A2(n1054), .A3(n1064), .ZN(n1210) );
AND3_X1 U917 ( .A1(n1223), .A2(n1246), .A3(n1078), .ZN(n1216) );
XOR2_X1 U918 ( .A(n1209), .B(n1247), .Z(G27) );
NAND2_X1 U919 ( .A1(KEYINPUT28), .A2(G125), .ZN(n1247) );
NAND2_X1 U920 ( .A1(n1248), .A2(n1234), .ZN(n1209) );
AND4_X1 U921 ( .A1(n1077), .A2(n1062), .A3(n1063), .A4(n1229), .ZN(n1234) );
NAND2_X1 U922 ( .A1(n1249), .A2(n1041), .ZN(n1229) );
NAND4_X1 U923 ( .A1(G902), .A2(G953), .A3(n1250), .A4(n1122), .ZN(n1249) );
INV_X1 U924 ( .A(G900), .ZN(n1122) );
XOR2_X1 U925 ( .A(n1251), .B(n1211), .Z(G24) );
NAND4_X1 U926 ( .A1(n1252), .A2(n1046), .A3(n1228), .A4(n1230), .ZN(n1211) );
NOR2_X1 U927 ( .A1(n1063), .A2(n1253), .ZN(n1046) );
XNOR2_X1 U928 ( .A(G119), .B(n1215), .ZN(G21) );
NAND4_X1 U929 ( .A1(n1245), .A2(n1252), .A3(n1054), .A4(n1063), .ZN(n1215) );
XOR2_X1 U930 ( .A(n1253), .B(KEYINPUT25), .Z(n1245) );
XNOR2_X1 U931 ( .A(G116), .B(n1214), .ZN(G18) );
NAND3_X1 U932 ( .A1(n1064), .A2(n1217), .A3(n1252), .ZN(n1214) );
INV_X1 U933 ( .A(n1076), .ZN(n1217) );
NAND2_X1 U934 ( .A1(n1254), .A2(n1228), .ZN(n1076) );
INV_X1 U935 ( .A(n1255), .ZN(n1228) );
XNOR2_X1 U936 ( .A(G113), .B(n1213), .ZN(G15) );
NAND3_X1 U937 ( .A1(n1064), .A2(n1077), .A3(n1252), .ZN(n1213) );
AND2_X1 U938 ( .A1(n1248), .A2(n1246), .ZN(n1252) );
AND3_X1 U939 ( .A1(n1044), .A2(n1045), .A3(n1223), .ZN(n1248) );
INV_X1 U940 ( .A(n1066), .ZN(n1223) );
INV_X1 U941 ( .A(n1042), .ZN(n1077) );
NOR2_X1 U942 ( .A1(n1062), .A2(n1063), .ZN(n1064) );
XOR2_X1 U943 ( .A(G110), .B(n1256), .Z(G12) );
NOR2_X1 U944 ( .A1(n1066), .A2(n1224), .ZN(n1256) );
NAND3_X1 U945 ( .A1(n1078), .A2(n1054), .A3(n1257), .ZN(n1224) );
AND3_X1 U946 ( .A1(n1062), .A2(n1246), .A3(n1063), .ZN(n1257) );
XOR2_X1 U947 ( .A(n1258), .B(n1157), .Z(n1063) );
NAND2_X1 U948 ( .A1(G217), .A2(n1259), .ZN(n1157) );
NAND2_X1 U949 ( .A1(n1155), .A2(n1260), .ZN(n1258) );
XNOR2_X1 U950 ( .A(n1261), .B(n1262), .ZN(n1155) );
XOR2_X1 U951 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U952 ( .A(n1198), .B(n1265), .Z(n1264) );
NAND2_X1 U953 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND4_X1 U954 ( .A1(n1268), .A2(G221), .A3(G234), .A4(n1048), .ZN(n1267) );
XOR2_X1 U955 ( .A(n1236), .B(KEYINPUT12), .Z(n1268) );
NAND2_X1 U956 ( .A1(n1269), .A2(n1270), .ZN(n1266) );
NAND3_X1 U957 ( .A1(G234), .A2(n1048), .A3(G221), .ZN(n1270) );
XOR2_X1 U958 ( .A(KEYINPUT20), .B(G137), .Z(n1269) );
XOR2_X1 U959 ( .A(n1271), .B(n1272), .Z(n1261) );
NAND2_X1 U960 ( .A1(n1041), .A2(n1273), .ZN(n1246) );
NAND3_X1 U961 ( .A1(n1142), .A2(n1250), .A3(G902), .ZN(n1273) );
NOR2_X1 U962 ( .A1(G898), .A2(n1048), .ZN(n1142) );
NAND3_X1 U963 ( .A1(n1250), .A2(n1048), .A3(G952), .ZN(n1041) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1250) );
INV_X1 U965 ( .A(n1253), .ZN(n1062) );
XNOR2_X1 U966 ( .A(n1095), .B(n1274), .ZN(n1253) );
NOR2_X1 U967 ( .A1(G472), .A2(KEYINPUT35), .ZN(n1274) );
AND2_X1 U968 ( .A1(n1275), .A2(n1260), .ZN(n1095) );
XOR2_X1 U969 ( .A(n1180), .B(n1276), .Z(n1275) );
XNOR2_X1 U970 ( .A(n1184), .B(n1183), .ZN(n1276) );
XOR2_X1 U971 ( .A(n1277), .B(n1278), .Z(n1184) );
XOR2_X1 U972 ( .A(n1263), .B(n1279), .Z(n1278) );
XOR2_X1 U973 ( .A(n1280), .B(G101), .Z(n1277) );
NAND2_X1 U974 ( .A1(G210), .A2(n1281), .ZN(n1280) );
NAND2_X1 U975 ( .A1(n1282), .A2(n1283), .ZN(n1054) );
OR2_X1 U976 ( .A1(n1042), .A2(KEYINPUT14), .ZN(n1283) );
NAND2_X1 U977 ( .A1(n1255), .A2(n1230), .ZN(n1042) );
NAND3_X1 U978 ( .A1(n1254), .A2(n1255), .A3(KEYINPUT14), .ZN(n1282) );
XOR2_X1 U979 ( .A(n1284), .B(n1285), .Z(n1255) );
XOR2_X1 U980 ( .A(KEYINPUT29), .B(G478), .Z(n1285) );
NAND2_X1 U981 ( .A1(n1286), .A2(KEYINPUT32), .ZN(n1284) );
XOR2_X1 U982 ( .A(n1088), .B(KEYINPUT57), .Z(n1286) );
NAND2_X1 U983 ( .A1(n1163), .A2(n1260), .ZN(n1088) );
XOR2_X1 U984 ( .A(n1287), .B(n1288), .Z(n1163) );
AND3_X1 U985 ( .A1(G234), .A2(n1048), .A3(G217), .ZN(n1288) );
NAND2_X1 U986 ( .A1(n1289), .A2(KEYINPUT37), .ZN(n1287) );
XOR2_X1 U987 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U988 ( .A(n1292), .B(n1272), .Z(n1291) );
INV_X1 U989 ( .A(n1293), .ZN(n1272) );
NOR2_X1 U990 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1292) );
XOR2_X1 U991 ( .A(n1294), .B(G143), .Z(n1290) );
NAND2_X1 U992 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U993 ( .A1(G107), .A2(n1297), .ZN(n1296) );
XOR2_X1 U994 ( .A(KEYINPUT4), .B(n1298), .Z(n1295) );
NOR2_X1 U995 ( .A1(G107), .A2(n1297), .ZN(n1298) );
XOR2_X1 U996 ( .A(G122), .B(G116), .Z(n1297) );
INV_X1 U997 ( .A(n1230), .ZN(n1254) );
NAND3_X1 U998 ( .A1(n1299), .A2(n1300), .A3(n1084), .ZN(n1230) );
NAND2_X1 U999 ( .A1(n1089), .A2(n1090), .ZN(n1084) );
NAND2_X1 U1000 ( .A1(n1090), .A2(n1301), .ZN(n1300) );
OR3_X1 U1001 ( .A1(n1090), .A2(n1089), .A3(n1301), .ZN(n1299) );
INV_X1 U1002 ( .A(KEYINPUT11), .ZN(n1301) );
AND2_X1 U1003 ( .A1(n1169), .A2(n1260), .ZN(n1089) );
XOR2_X1 U1004 ( .A(n1302), .B(KEYINPUT39), .Z(n1169) );
XOR2_X1 U1005 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1006 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1007 ( .A(G131), .B(G122), .Z(n1306) );
XOR2_X1 U1008 ( .A(KEYINPUT42), .B(G143), .Z(n1305) );
XOR2_X1 U1009 ( .A(n1307), .B(n1308), .Z(n1303) );
XOR2_X1 U1010 ( .A(G113), .B(n1309), .Z(n1308) );
NOR2_X1 U1011 ( .A1(G104), .A2(KEYINPUT53), .ZN(n1309) );
XOR2_X1 U1012 ( .A(n1271), .B(n1310), .Z(n1307) );
AND2_X1 U1013 ( .A1(n1281), .A2(G214), .ZN(n1310) );
NOR2_X1 U1014 ( .A1(G953), .A2(G237), .ZN(n1281) );
XOR2_X1 U1015 ( .A(n1225), .B(n1131), .Z(n1271) );
XOR2_X1 U1016 ( .A(G125), .B(G140), .Z(n1131) );
XNOR2_X1 U1017 ( .A(n1172), .B(KEYINPUT41), .ZN(n1090) );
INV_X1 U1018 ( .A(G475), .ZN(n1172) );
NOR2_X1 U1019 ( .A1(n1044), .A2(n1311), .ZN(n1078) );
INV_X1 U1020 ( .A(n1045), .ZN(n1311) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1259), .ZN(n1045) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U1023 ( .A(n1197), .B(n1312), .ZN(n1044) );
NOR2_X1 U1024 ( .A1(n1106), .A2(KEYINPUT36), .ZN(n1312) );
AND2_X1 U1025 ( .A1(n1313), .A2(n1260), .ZN(n1106) );
XOR2_X1 U1026 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1027 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND2_X1 U1028 ( .A1(KEYINPUT50), .A2(G140), .ZN(n1317) );
NAND2_X1 U1029 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
NAND2_X1 U1030 ( .A1(n1320), .A2(n1134), .ZN(n1319) );
XOR2_X1 U1031 ( .A(KEYINPUT19), .B(n1321), .Z(n1318) );
NOR2_X1 U1032 ( .A1(n1134), .A2(n1320), .ZN(n1321) );
XOR2_X1 U1033 ( .A(n1187), .B(KEYINPUT55), .Z(n1320) );
XNOR2_X1 U1034 ( .A(n1322), .B(n1293), .ZN(n1134) );
NAND2_X1 U1035 ( .A1(KEYINPUT43), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1036 ( .A(n1183), .B(n1324), .Z(n1314) );
XOR2_X1 U1037 ( .A(n1198), .B(n1325), .Z(n1324) );
NOR2_X1 U1038 ( .A1(KEYINPUT7), .A2(n1121), .ZN(n1325) );
INV_X1 U1039 ( .A(G227), .ZN(n1121) );
INV_X1 U1040 ( .A(G110), .ZN(n1198) );
NAND2_X1 U1041 ( .A1(n1326), .A2(n1327), .ZN(n1183) );
NAND2_X1 U1042 ( .A1(G131), .A2(n1130), .ZN(n1327) );
XOR2_X1 U1043 ( .A(n1328), .B(KEYINPUT58), .Z(n1326) );
OR2_X1 U1044 ( .A1(n1130), .A2(G131), .ZN(n1328) );
XOR2_X1 U1045 ( .A(n1238), .B(n1236), .Z(n1130) );
INV_X1 U1046 ( .A(G137), .ZN(n1236) );
INV_X1 U1047 ( .A(G134), .ZN(n1238) );
INV_X1 U1048 ( .A(G469), .ZN(n1197) );
NAND2_X1 U1049 ( .A1(n1069), .A2(n1068), .ZN(n1066) );
NAND2_X1 U1050 ( .A1(G214), .A2(n1329), .ZN(n1068) );
XOR2_X1 U1051 ( .A(n1109), .B(n1116), .Z(n1069) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1329), .ZN(n1116) );
NAND2_X1 U1053 ( .A1(n1330), .A2(n1260), .ZN(n1329) );
INV_X1 U1054 ( .A(G237), .ZN(n1330) );
NAND2_X1 U1055 ( .A1(n1331), .A2(n1260), .ZN(n1109) );
INV_X1 U1056 ( .A(G902), .ZN(n1260) );
XOR2_X1 U1057 ( .A(n1332), .B(n1203), .Z(n1331) );
XOR2_X1 U1058 ( .A(n1146), .B(n1333), .Z(n1203) );
XOR2_X1 U1059 ( .A(n1334), .B(n1335), .Z(n1333) );
NAND2_X1 U1060 ( .A1(KEYINPUT51), .A2(n1145), .ZN(n1335) );
NAND2_X1 U1061 ( .A1(n1336), .A2(n1337), .ZN(n1145) );
NAND2_X1 U1062 ( .A1(n1279), .A2(n1338), .ZN(n1337) );
NAND2_X1 U1063 ( .A1(n1263), .A2(n1339), .ZN(n1336) );
XNOR2_X1 U1064 ( .A(n1279), .B(KEYINPUT62), .ZN(n1339) );
XOR2_X1 U1065 ( .A(G113), .B(G116), .Z(n1279) );
INV_X1 U1066 ( .A(n1338), .ZN(n1263) );
XNOR2_X1 U1067 ( .A(G119), .B(KEYINPUT13), .ZN(n1338) );
NAND2_X1 U1068 ( .A1(G224), .A2(n1048), .ZN(n1334) );
INV_X1 U1069 ( .A(G953), .ZN(n1048) );
XOR2_X1 U1070 ( .A(n1340), .B(n1341), .Z(n1146) );
XOR2_X1 U1071 ( .A(n1251), .B(n1342), .Z(n1341) );
XNOR2_X1 U1072 ( .A(KEYINPUT54), .B(KEYINPUT22), .ZN(n1342) );
INV_X1 U1073 ( .A(G122), .ZN(n1251) );
XOR2_X1 U1074 ( .A(n1187), .B(G110), .Z(n1340) );
XNOR2_X1 U1075 ( .A(G101), .B(n1343), .ZN(n1187) );
XOR2_X1 U1076 ( .A(G107), .B(G104), .Z(n1343) );
NAND2_X1 U1077 ( .A1(KEYINPUT33), .A2(n1201), .ZN(n1332) );
XOR2_X1 U1078 ( .A(n1180), .B(G125), .Z(n1201) );
NAND2_X1 U1079 ( .A1(n1344), .A2(n1345), .ZN(n1180) );
NAND2_X1 U1080 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
INV_X1 U1081 ( .A(KEYINPUT6), .ZN(n1347) );
XOR2_X1 U1082 ( .A(n1323), .B(n1293), .Z(n1346) );
XNOR2_X1 U1083 ( .A(n1225), .B(n1348), .ZN(n1323) );
NAND2_X1 U1084 ( .A1(n1349), .A2(KEYINPUT6), .ZN(n1344) );
XOR2_X1 U1085 ( .A(n1350), .B(n1293), .Z(n1349) );
XNOR2_X1 U1086 ( .A(G128), .B(KEYINPUT52), .ZN(n1293) );
NAND2_X1 U1087 ( .A1(n1348), .A2(n1225), .ZN(n1350) );
INV_X1 U1088 ( .A(G146), .ZN(n1225) );
XOR2_X1 U1089 ( .A(G143), .B(KEYINPUT56), .Z(n1348) );
endmodule


