//Key = 1011101110111111110011000101101110011001110100011111010111001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416;

NAND2_X1 U784 ( .A1(n1080), .A2(n1081), .ZN(G9) );
NAND2_X1 U785 ( .A1(G107), .A2(n1082), .ZN(n1081) );
XOR2_X1 U786 ( .A(KEYINPUT20), .B(n1083), .Z(n1080) );
NOR2_X1 U787 ( .A1(G107), .A2(n1082), .ZN(n1083) );
NAND2_X1 U788 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
XNOR2_X1 U789 ( .A(KEYINPUT18), .B(n1086), .ZN(n1085) );
INV_X1 U790 ( .A(n1087), .ZN(n1084) );
NAND3_X1 U791 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(G75) );
NAND2_X1 U792 ( .A1(G952), .A2(n1091), .ZN(n1090) );
NAND4_X1 U793 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
NAND3_X1 U794 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
NAND2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
NAND3_X1 U796 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NAND2_X1 U797 ( .A1(n1098), .A2(n1104), .ZN(n1103) );
INV_X1 U798 ( .A(n1105), .ZN(n1098) );
NAND4_X1 U799 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1102) );
NAND2_X1 U800 ( .A1(KEYINPUT27), .A2(n1105), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
NAND2_X1 U802 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
INV_X1 U803 ( .A(KEYINPUT27), .ZN(n1113) );
NAND2_X1 U804 ( .A1(n1110), .A2(n1114), .ZN(n1112) );
NAND3_X1 U805 ( .A1(n1115), .A2(n1111), .A3(n1096), .ZN(n1101) );
NAND2_X1 U806 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND3_X1 U807 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NAND3_X1 U809 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1118) );
INV_X1 U810 ( .A(n1126), .ZN(n1124) );
NAND2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
NAND2_X1 U812 ( .A1(n1129), .A2(n1130), .ZN(n1116) );
NAND4_X1 U813 ( .A1(n1130), .A2(n1106), .A3(n1131), .A4(n1132), .ZN(n1088) );
NOR4_X1 U814 ( .A1(n1107), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1132) );
XOR2_X1 U815 ( .A(n1136), .B(n1137), .Z(n1133) );
NAND2_X1 U816 ( .A1(KEYINPUT36), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U817 ( .A(n1139), .B(n1140), .ZN(n1131) );
XOR2_X1 U818 ( .A(n1141), .B(n1142), .Z(G72) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U821 ( .A1(G953), .A2(n1147), .ZN(n1146) );
XNOR2_X1 U822 ( .A(KEYINPUT57), .B(n1148), .ZN(n1147) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1145) );
XNOR2_X1 U824 ( .A(n1151), .B(n1152), .ZN(n1150) );
XNOR2_X1 U825 ( .A(n1153), .B(G134), .ZN(n1152) );
XNOR2_X1 U826 ( .A(n1154), .B(n1155), .ZN(n1149) );
XOR2_X1 U827 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U828 ( .A1(KEYINPUT7), .A2(n1158), .ZN(n1157) );
NAND2_X1 U829 ( .A1(n1089), .A2(n1159), .ZN(n1143) );
NAND4_X1 U830 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1164), .A2(n1089), .ZN(n1141) );
NOR2_X1 U832 ( .A1(n1165), .A2(n1148), .ZN(n1164) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(G69) );
XOR2_X1 U834 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U835 ( .A1(G953), .A2(n1170), .ZN(n1169) );
NAND2_X1 U836 ( .A1(G898), .A2(G224), .ZN(n1170) );
NAND2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
NAND2_X1 U838 ( .A1(G953), .A2(n1173), .ZN(n1172) );
XOR2_X1 U839 ( .A(n1174), .B(n1175), .Z(n1171) );
XOR2_X1 U840 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U841 ( .A1(KEYINPUT60), .A2(n1178), .ZN(n1177) );
XOR2_X1 U842 ( .A(G113), .B(n1179), .Z(n1174) );
NOR2_X1 U843 ( .A1(KEYINPUT52), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U844 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U845 ( .A1(n1093), .A2(G953), .ZN(n1166) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1184), .ZN(G66) );
NOR3_X1 U847 ( .A1(n1139), .A2(n1185), .A3(n1186), .ZN(n1184) );
NOR3_X1 U848 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NOR2_X1 U849 ( .A1(n1190), .A2(n1191), .ZN(n1185) );
AND2_X1 U850 ( .A1(n1192), .A2(n1140), .ZN(n1190) );
NOR2_X1 U851 ( .A1(n1183), .A2(n1193), .ZN(G63) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U853 ( .A1(n1189), .A2(n1138), .ZN(n1195) );
NAND2_X1 U854 ( .A1(KEYINPUT47), .A2(n1196), .ZN(n1194) );
NOR2_X1 U855 ( .A1(n1183), .A2(n1197), .ZN(G60) );
XNOR2_X1 U856 ( .A(n1198), .B(n1199), .ZN(n1197) );
NOR2_X1 U857 ( .A1(n1189), .A2(n1200), .ZN(n1199) );
XOR2_X1 U858 ( .A(KEYINPUT50), .B(G475), .Z(n1200) );
XOR2_X1 U859 ( .A(G104), .B(n1201), .Z(G6) );
NOR3_X1 U860 ( .A1(n1202), .A2(KEYINPUT46), .A3(n1087), .ZN(n1201) );
NOR2_X1 U861 ( .A1(n1183), .A2(n1203), .ZN(G57) );
XOR2_X1 U862 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U863 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U864 ( .A(KEYINPUT3), .B(n1208), .Z(n1207) );
NOR2_X1 U865 ( .A1(n1209), .A2(n1189), .ZN(n1206) );
XOR2_X1 U866 ( .A(n1210), .B(n1211), .Z(n1204) );
XNOR2_X1 U867 ( .A(n1212), .B(n1213), .ZN(n1211) );
NOR2_X1 U868 ( .A1(n1183), .A2(n1214), .ZN(G54) );
XOR2_X1 U869 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U870 ( .A(n1217), .B(n1218), .ZN(n1216) );
NOR2_X1 U871 ( .A1(n1219), .A2(n1189), .ZN(n1217) );
XOR2_X1 U872 ( .A(n1220), .B(n1221), .Z(n1215) );
NAND2_X1 U873 ( .A1(n1222), .A2(KEYINPUT41), .ZN(n1221) );
XOR2_X1 U874 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U875 ( .A(n1156), .B(KEYINPUT32), .Z(n1223) );
NAND2_X1 U876 ( .A1(n1225), .A2(KEYINPUT17), .ZN(n1220) );
XOR2_X1 U877 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U878 ( .A1(KEYINPUT61), .A2(n1153), .ZN(n1227) );
XNOR2_X1 U879 ( .A(G110), .B(n1228), .ZN(n1226) );
NOR2_X1 U880 ( .A1(n1183), .A2(n1229), .ZN(G51) );
XOR2_X1 U881 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U882 ( .A1(n1232), .A2(n1189), .ZN(n1230) );
NAND2_X1 U883 ( .A1(G902), .A2(n1192), .ZN(n1189) );
NAND2_X1 U884 ( .A1(n1092), .A2(n1233), .ZN(n1192) );
XOR2_X1 U885 ( .A(KEYINPUT23), .B(n1093), .Z(n1233) );
AND4_X1 U886 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1093) );
NOR2_X1 U887 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
NAND2_X1 U888 ( .A1(n1097), .A2(n1240), .ZN(n1234) );
NAND2_X1 U889 ( .A1(n1241), .A2(n1087), .ZN(n1240) );
NAND2_X1 U890 ( .A1(n1242), .A2(n1125), .ZN(n1087) );
NAND2_X1 U891 ( .A1(n1202), .A2(n1086), .ZN(n1097) );
INV_X1 U892 ( .A(n1243), .ZN(n1202) );
AND4_X1 U893 ( .A1(n1244), .A2(n1160), .A3(n1162), .A4(n1163), .ZN(n1092) );
NAND2_X1 U894 ( .A1(n1245), .A2(n1126), .ZN(n1162) );
AND3_X1 U895 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1160) );
NOR3_X1 U896 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1248) );
XOR2_X1 U897 ( .A(n1161), .B(KEYINPUT33), .Z(n1244) );
NAND3_X1 U898 ( .A1(n1126), .A2(n1252), .A3(n1253), .ZN(n1161) );
INV_X1 U899 ( .A(n1254), .ZN(n1253) );
XNOR2_X1 U900 ( .A(KEYINPUT1), .B(n1255), .ZN(n1252) );
NOR2_X1 U901 ( .A1(n1089), .A2(G952), .ZN(n1183) );
XNOR2_X1 U902 ( .A(G146), .B(n1246), .ZN(G48) );
NAND3_X1 U903 ( .A1(n1256), .A2(n1104), .A3(n1243), .ZN(n1246) );
XOR2_X1 U904 ( .A(G143), .B(n1257), .Z(G45) );
NOR3_X1 U905 ( .A1(n1254), .A2(n1258), .A3(n1255), .ZN(n1257) );
XNOR2_X1 U906 ( .A(n1126), .B(KEYINPUT59), .ZN(n1258) );
NAND4_X1 U907 ( .A1(n1259), .A2(n1129), .A3(n1260), .A4(n1261), .ZN(n1254) );
XNOR2_X1 U908 ( .A(G140), .B(n1247), .ZN(G42) );
NAND3_X1 U909 ( .A1(n1096), .A2(n1126), .A3(n1262), .ZN(n1247) );
XNOR2_X1 U910 ( .A(n1158), .B(n1249), .ZN(G39) );
AND3_X1 U911 ( .A1(n1096), .A2(n1256), .A3(n1099), .ZN(n1249) );
INV_X1 U912 ( .A(G137), .ZN(n1158) );
XOR2_X1 U913 ( .A(G134), .B(n1251), .Z(G36) );
AND4_X1 U914 ( .A1(n1126), .A2(n1261), .A3(n1263), .A4(n1264), .ZN(n1251) );
AND2_X1 U915 ( .A1(n1096), .A2(n1129), .ZN(n1264) );
NAND3_X1 U916 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(G33) );
OR2_X1 U917 ( .A1(n1268), .A2(G131), .ZN(n1267) );
NAND2_X1 U918 ( .A1(KEYINPUT37), .A2(n1269), .ZN(n1266) );
NAND2_X1 U919 ( .A1(n1270), .A2(n1268), .ZN(n1269) );
XNOR2_X1 U920 ( .A(KEYINPUT39), .B(G131), .ZN(n1270) );
NAND2_X1 U921 ( .A1(n1271), .A2(n1272), .ZN(n1265) );
INV_X1 U922 ( .A(KEYINPUT37), .ZN(n1272) );
NAND2_X1 U923 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
OR2_X1 U924 ( .A1(G131), .A2(KEYINPUT39), .ZN(n1274) );
NAND3_X1 U925 ( .A1(G131), .A2(n1268), .A3(KEYINPUT39), .ZN(n1273) );
NAND2_X1 U926 ( .A1(n1275), .A2(n1245), .ZN(n1268) );
AND4_X1 U927 ( .A1(n1243), .A2(n1129), .A3(n1096), .A4(n1261), .ZN(n1245) );
AND2_X1 U928 ( .A1(n1276), .A2(n1277), .ZN(n1096) );
XNOR2_X1 U929 ( .A(n1106), .B(KEYINPUT0), .ZN(n1276) );
INV_X1 U930 ( .A(n1278), .ZN(n1106) );
XNOR2_X1 U931 ( .A(n1126), .B(KEYINPUT43), .ZN(n1275) );
XNOR2_X1 U932 ( .A(n1279), .B(n1250), .ZN(G30) );
AND3_X1 U933 ( .A1(n1263), .A2(n1104), .A3(n1256), .ZN(n1250) );
AND4_X1 U934 ( .A1(n1126), .A2(n1121), .A3(n1135), .A4(n1261), .ZN(n1256) );
INV_X1 U935 ( .A(n1086), .ZN(n1263) );
XNOR2_X1 U936 ( .A(G101), .B(n1235), .ZN(G3) );
NAND4_X1 U937 ( .A1(n1099), .A2(n1129), .A3(n1126), .A4(n1280), .ZN(n1235) );
XNOR2_X1 U938 ( .A(n1281), .B(n1151), .ZN(G27) );
NAND2_X1 U939 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
OR2_X1 U940 ( .A1(n1163), .A2(KEYINPUT24), .ZN(n1283) );
NAND3_X1 U941 ( .A1(n1130), .A2(n1104), .A3(n1262), .ZN(n1163) );
NAND4_X1 U942 ( .A1(n1130), .A2(n1255), .A3(n1262), .A4(KEYINPUT24), .ZN(n1282) );
AND4_X1 U943 ( .A1(n1120), .A2(n1243), .A3(n1121), .A4(n1261), .ZN(n1262) );
NAND2_X1 U944 ( .A1(n1284), .A2(n1285), .ZN(n1261) );
NAND2_X1 U945 ( .A1(n1286), .A2(n1148), .ZN(n1285) );
INV_X1 U946 ( .A(G900), .ZN(n1148) );
NAND2_X1 U947 ( .A1(n1287), .A2(n1288), .ZN(G24) );
NAND2_X1 U948 ( .A1(n1238), .A2(n1289), .ZN(n1288) );
XOR2_X1 U949 ( .A(KEYINPUT8), .B(n1290), .Z(n1287) );
NOR2_X1 U950 ( .A1(n1238), .A2(n1289), .ZN(n1290) );
AND4_X1 U951 ( .A1(n1259), .A2(n1110), .A3(n1280), .A4(n1260), .ZN(n1238) );
NOR3_X1 U952 ( .A1(n1135), .A2(n1121), .A3(n1122), .ZN(n1110) );
XOR2_X1 U953 ( .A(n1291), .B(G119), .Z(G21) );
NAND2_X1 U954 ( .A1(KEYINPUT28), .A2(n1237), .ZN(n1291) );
NAND4_X1 U955 ( .A1(n1099), .A2(n1130), .A3(n1292), .A4(n1280), .ZN(n1237) );
NOR2_X1 U956 ( .A1(n1120), .A2(n1125), .ZN(n1292) );
INV_X1 U957 ( .A(n1121), .ZN(n1125) );
XNOR2_X1 U958 ( .A(n1293), .B(n1294), .ZN(G18) );
NOR2_X1 U959 ( .A1(n1086), .A2(n1241), .ZN(n1294) );
NAND2_X1 U960 ( .A1(n1259), .A2(n1295), .ZN(n1086) );
XOR2_X1 U961 ( .A(G113), .B(n1296), .Z(G15) );
NOR2_X1 U962 ( .A1(n1297), .A2(n1241), .ZN(n1296) );
NAND3_X1 U963 ( .A1(n1130), .A2(n1280), .A3(n1129), .ZN(n1241) );
NOR2_X1 U964 ( .A1(n1121), .A2(n1120), .ZN(n1129) );
INV_X1 U965 ( .A(n1122), .ZN(n1130) );
NAND2_X1 U966 ( .A1(n1128), .A2(n1298), .ZN(n1122) );
XNOR2_X1 U967 ( .A(n1243), .B(KEYINPUT45), .ZN(n1297) );
NOR2_X1 U968 ( .A1(n1295), .A2(n1259), .ZN(n1243) );
INV_X1 U969 ( .A(n1260), .ZN(n1295) );
NAND2_X1 U970 ( .A1(n1299), .A2(n1300), .ZN(G12) );
NAND2_X1 U971 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
INV_X1 U972 ( .A(G110), .ZN(n1302) );
NAND2_X1 U973 ( .A1(G110), .A2(n1303), .ZN(n1299) );
NAND2_X1 U974 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U975 ( .A1(n1239), .A2(n1306), .ZN(n1305) );
INV_X1 U976 ( .A(n1307), .ZN(n1239) );
OR2_X1 U977 ( .A1(n1306), .A2(n1301), .ZN(n1304) );
NOR2_X1 U978 ( .A1(KEYINPUT9), .A2(n1307), .ZN(n1301) );
NAND3_X1 U979 ( .A1(n1242), .A2(n1121), .A3(n1099), .ZN(n1307) );
NOR2_X1 U980 ( .A1(n1260), .A2(n1259), .ZN(n1099) );
XOR2_X1 U981 ( .A(n1308), .B(n1137), .Z(n1259) );
AND2_X1 U982 ( .A1(n1196), .A2(n1309), .ZN(n1137) );
XOR2_X1 U983 ( .A(n1310), .B(n1311), .Z(n1196) );
XNOR2_X1 U984 ( .A(n1279), .B(G122), .ZN(n1311) );
XNOR2_X1 U985 ( .A(n1312), .B(n1293), .ZN(n1310) );
XOR2_X1 U986 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U987 ( .A(G143), .B(n1315), .ZN(n1314) );
XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT19), .ZN(n1315) );
XOR2_X1 U989 ( .A(n1316), .B(n1317), .Z(n1313) );
XOR2_X1 U990 ( .A(G134), .B(G107), .Z(n1317) );
NAND3_X1 U991 ( .A1(G234), .A2(n1089), .A3(G217), .ZN(n1316) );
NAND2_X1 U992 ( .A1(KEYINPUT51), .A2(n1138), .ZN(n1308) );
INV_X1 U993 ( .A(G478), .ZN(n1138) );
XOR2_X1 U994 ( .A(n1134), .B(KEYINPUT63), .Z(n1260) );
XNOR2_X1 U995 ( .A(n1318), .B(G475), .ZN(n1134) );
NAND2_X1 U996 ( .A1(n1198), .A2(n1309), .ZN(n1318) );
XNOR2_X1 U997 ( .A(n1319), .B(n1320), .ZN(n1198) );
XOR2_X1 U998 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U999 ( .A(G113), .B(G104), .Z(n1322) );
XNOR2_X1 U1000 ( .A(KEYINPUT11), .B(n1289), .ZN(n1321) );
INV_X1 U1001 ( .A(G122), .ZN(n1289) );
XOR2_X1 U1002 ( .A(n1323), .B(n1324), .Z(n1319) );
XOR2_X1 U1003 ( .A(n1325), .B(n1326), .Z(n1324) );
NAND2_X1 U1004 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1005 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XNOR2_X1 U1006 ( .A(KEYINPUT12), .B(n1153), .ZN(n1330) );
INV_X1 U1007 ( .A(G140), .ZN(n1153) );
XNOR2_X1 U1008 ( .A(G125), .B(KEYINPUT29), .ZN(n1329) );
NAND2_X1 U1009 ( .A1(n1331), .A2(n1332), .ZN(n1327) );
XNOR2_X1 U1010 ( .A(G125), .B(KEYINPUT49), .ZN(n1332) );
XNOR2_X1 U1011 ( .A(KEYINPUT12), .B(G140), .ZN(n1331) );
NAND3_X1 U1012 ( .A1(n1333), .A2(n1089), .A3(G214), .ZN(n1325) );
XNOR2_X1 U1013 ( .A(n1334), .B(n1154), .ZN(n1323) );
XOR2_X1 U1014 ( .A(n1335), .B(n1336), .Z(n1121) );
INV_X1 U1015 ( .A(n1139), .ZN(n1336) );
NOR2_X1 U1016 ( .A1(n1191), .A2(G902), .ZN(n1139) );
INV_X1 U1017 ( .A(n1187), .ZN(n1191) );
XNOR2_X1 U1018 ( .A(n1337), .B(n1338), .ZN(n1187) );
XOR2_X1 U1019 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1020 ( .A(n1341), .B(n1342), .Z(n1340) );
NOR2_X1 U1021 ( .A1(KEYINPUT26), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1022 ( .A(KEYINPUT11), .B(n1344), .Z(n1343) );
NAND3_X1 U1023 ( .A1(G234), .A2(n1089), .A3(G221), .ZN(n1341) );
XOR2_X1 U1024 ( .A(n1345), .B(n1346), .Z(n1337) );
XNOR2_X1 U1025 ( .A(n1151), .B(G119), .ZN(n1346) );
XNOR2_X1 U1026 ( .A(G137), .B(G128), .ZN(n1345) );
NAND2_X1 U1027 ( .A1(KEYINPUT53), .A2(n1140), .ZN(n1335) );
INV_X1 U1028 ( .A(n1188), .ZN(n1140) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1347), .ZN(n1188) );
AND3_X1 U1030 ( .A1(n1120), .A2(n1280), .A3(n1126), .ZN(n1242) );
NOR2_X1 U1031 ( .A1(n1128), .A2(n1127), .ZN(n1126) );
INV_X1 U1032 ( .A(n1298), .ZN(n1127) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1347), .ZN(n1298) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1309), .ZN(n1347) );
XNOR2_X1 U1035 ( .A(n1348), .B(n1219), .ZN(n1128) );
INV_X1 U1036 ( .A(G469), .ZN(n1219) );
NAND2_X1 U1037 ( .A1(n1349), .A2(n1309), .ZN(n1348) );
XOR2_X1 U1038 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1039 ( .A(n1352), .B(n1218), .ZN(n1351) );
NAND2_X1 U1040 ( .A1(KEYINPUT30), .A2(n1224), .ZN(n1352) );
XNOR2_X1 U1041 ( .A(n1353), .B(n1181), .ZN(n1224) );
NAND2_X1 U1042 ( .A1(KEYINPUT25), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1043 ( .A(n1355), .B(n1356), .Z(n1350) );
NOR2_X1 U1044 ( .A1(KEYINPUT54), .A2(n1339), .ZN(n1356) );
XNOR2_X1 U1045 ( .A(G110), .B(G140), .ZN(n1339) );
XOR2_X1 U1046 ( .A(n1156), .B(n1228), .Z(n1355) );
NOR2_X1 U1047 ( .A1(n1165), .A2(G953), .ZN(n1228) );
INV_X1 U1048 ( .A(G227), .ZN(n1165) );
NAND3_X1 U1049 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1156) );
NAND2_X1 U1050 ( .A1(n1360), .A2(n1279), .ZN(n1359) );
NAND2_X1 U1051 ( .A1(KEYINPUT22), .A2(n1361), .ZN(n1358) );
NAND2_X1 U1052 ( .A1(n1362), .A2(n1334), .ZN(n1361) );
XNOR2_X1 U1053 ( .A(KEYINPUT62), .B(n1279), .ZN(n1362) );
NAND2_X1 U1054 ( .A1(n1363), .A2(n1364), .ZN(n1357) );
INV_X1 U1055 ( .A(KEYINPUT22), .ZN(n1364) );
NAND2_X1 U1056 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
OR3_X1 U1057 ( .A1(n1279), .A2(n1360), .A3(KEYINPUT62), .ZN(n1366) );
INV_X1 U1058 ( .A(n1334), .ZN(n1360) );
NAND2_X1 U1059 ( .A1(KEYINPUT62), .A2(n1279), .ZN(n1365) );
INV_X1 U1060 ( .A(G128), .ZN(n1279) );
AND2_X1 U1061 ( .A1(n1104), .A2(n1367), .ZN(n1280) );
NAND2_X1 U1062 ( .A1(n1284), .A2(n1368), .ZN(n1367) );
NAND2_X1 U1063 ( .A1(n1286), .A2(n1173), .ZN(n1368) );
INV_X1 U1064 ( .A(G898), .ZN(n1173) );
NOR3_X1 U1065 ( .A1(n1309), .A2(n1114), .A3(n1089), .ZN(n1286) );
INV_X1 U1066 ( .A(n1111), .ZN(n1114) );
NAND3_X1 U1067 ( .A1(n1369), .A2(n1089), .A3(G952), .ZN(n1284) );
XNOR2_X1 U1068 ( .A(KEYINPUT55), .B(n1111), .ZN(n1369) );
NAND2_X1 U1069 ( .A1(G237), .A2(G234), .ZN(n1111) );
INV_X1 U1070 ( .A(n1255), .ZN(n1104) );
NAND2_X1 U1071 ( .A1(n1277), .A2(n1278), .ZN(n1255) );
NAND2_X1 U1072 ( .A1(n1370), .A2(n1371), .ZN(n1278) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1372), .ZN(n1371) );
NAND2_X1 U1074 ( .A1(n1309), .A2(n1373), .ZN(n1372) );
OR2_X1 U1075 ( .A1(n1333), .A2(n1374), .ZN(n1373) );
NAND3_X1 U1076 ( .A1(n1375), .A2(n1309), .A3(n1374), .ZN(n1370) );
XOR2_X1 U1077 ( .A(n1231), .B(KEYINPUT2), .Z(n1374) );
XNOR2_X1 U1078 ( .A(n1376), .B(n1377), .ZN(n1231) );
XOR2_X1 U1079 ( .A(n1378), .B(n1379), .Z(n1377) );
XOR2_X1 U1080 ( .A(n1176), .B(n1380), .Z(n1379) );
NAND2_X1 U1081 ( .A1(G224), .A2(n1089), .ZN(n1380) );
INV_X1 U1082 ( .A(G953), .ZN(n1089) );
NAND3_X1 U1083 ( .A1(n1381), .A2(n1382), .A3(KEYINPUT21), .ZN(n1176) );
NAND2_X1 U1084 ( .A1(G119), .A2(n1293), .ZN(n1382) );
XOR2_X1 U1085 ( .A(KEYINPUT4), .B(n1383), .Z(n1381) );
NOR2_X1 U1086 ( .A1(G119), .A2(n1293), .ZN(n1383) );
XNOR2_X1 U1087 ( .A(KEYINPUT56), .B(n1151), .ZN(n1378) );
INV_X1 U1088 ( .A(G125), .ZN(n1151) );
XOR2_X1 U1089 ( .A(n1384), .B(n1385), .Z(n1376) );
NOR2_X1 U1090 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
AND2_X1 U1091 ( .A1(KEYINPUT40), .A2(n1178), .ZN(n1387) );
NOR2_X1 U1092 ( .A1(KEYINPUT6), .A2(n1178), .ZN(n1386) );
XNOR2_X1 U1093 ( .A(G110), .B(n1388), .ZN(n1178) );
NOR2_X1 U1094 ( .A1(G122), .A2(KEYINPUT38), .ZN(n1388) );
XNOR2_X1 U1095 ( .A(n1210), .B(n1389), .ZN(n1384) );
INV_X1 U1096 ( .A(n1181), .ZN(n1389) );
XOR2_X1 U1097 ( .A(G104), .B(G107), .Z(n1181) );
XNOR2_X1 U1098 ( .A(n1390), .B(n1354), .ZN(n1210) );
INV_X1 U1099 ( .A(n1182), .ZN(n1354) );
XOR2_X1 U1100 ( .A(n1391), .B(G113), .Z(n1390) );
NAND2_X1 U1101 ( .A1(G210), .A2(G237), .ZN(n1375) );
XOR2_X1 U1102 ( .A(KEYINPUT31), .B(n1107), .Z(n1277) );
AND2_X1 U1103 ( .A1(G214), .A2(n1392), .ZN(n1107) );
NAND2_X1 U1104 ( .A1(n1309), .A2(n1333), .ZN(n1392) );
INV_X1 U1105 ( .A(G237), .ZN(n1333) );
INV_X1 U1106 ( .A(n1135), .ZN(n1120) );
XOR2_X1 U1107 ( .A(n1393), .B(n1209), .Z(n1135) );
INV_X1 U1108 ( .A(G472), .ZN(n1209) );
NAND2_X1 U1109 ( .A1(n1394), .A2(n1309), .ZN(n1393) );
INV_X1 U1110 ( .A(G902), .ZN(n1309) );
XOR2_X1 U1111 ( .A(n1395), .B(n1396), .Z(n1394) );
XNOR2_X1 U1112 ( .A(n1208), .B(n1397), .ZN(n1396) );
NAND2_X1 U1113 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
NAND2_X1 U1114 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
NAND2_X1 U1115 ( .A1(KEYINPUT13), .A2(n1402), .ZN(n1401) );
NAND2_X1 U1116 ( .A1(KEYINPUT16), .A2(n1403), .ZN(n1402) );
INV_X1 U1117 ( .A(n1404), .ZN(n1403) );
INV_X1 U1118 ( .A(n1405), .ZN(n1400) );
NAND2_X1 U1119 ( .A1(n1404), .A2(n1406), .ZN(n1398) );
NAND2_X1 U1120 ( .A1(KEYINPUT16), .A2(n1407), .ZN(n1406) );
NAND2_X1 U1121 ( .A1(KEYINPUT13), .A2(n1405), .ZN(n1407) );
XNOR2_X1 U1122 ( .A(n1213), .B(G113), .ZN(n1405) );
XOR2_X1 U1123 ( .A(n1408), .B(KEYINPUT35), .Z(n1213) );
NAND3_X1 U1124 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(n1408) );
NAND2_X1 U1125 ( .A1(G116), .A2(n1412), .ZN(n1411) );
NAND2_X1 U1126 ( .A1(KEYINPUT10), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1127 ( .A(KEYINPUT44), .B(G119), .Z(n1413) );
NAND3_X1 U1128 ( .A1(KEYINPUT10), .A2(n1293), .A3(G119), .ZN(n1410) );
INV_X1 U1129 ( .A(G116), .ZN(n1293) );
OR2_X1 U1130 ( .A1(G119), .A2(KEYINPUT10), .ZN(n1409) );
XNOR2_X1 U1131 ( .A(n1391), .B(n1414), .ZN(n1404) );
XNOR2_X1 U1132 ( .A(KEYINPUT34), .B(n1218), .ZN(n1414) );
INV_X1 U1133 ( .A(n1212), .ZN(n1218) );
XOR2_X1 U1134 ( .A(n1415), .B(n1416), .Z(n1212) );
INV_X1 U1135 ( .A(n1154), .ZN(n1416) );
XOR2_X1 U1136 ( .A(G131), .B(KEYINPUT14), .Z(n1154) );
XNOR2_X1 U1137 ( .A(G134), .B(G137), .ZN(n1415) );
XNOR2_X1 U1138 ( .A(G128), .B(n1334), .ZN(n1391) );
XOR2_X1 U1139 ( .A(G143), .B(n1344), .Z(n1334) );
XOR2_X1 U1140 ( .A(G146), .B(KEYINPUT5), .Z(n1344) );
NOR3_X1 U1141 ( .A1(G237), .A2(G953), .A3(n1232), .ZN(n1208) );
INV_X1 U1142 ( .A(G210), .ZN(n1232) );
NOR2_X1 U1143 ( .A1(KEYINPUT42), .A2(n1182), .ZN(n1395) );
XOR2_X1 U1144 ( .A(G101), .B(KEYINPUT58), .Z(n1182) );
INV_X1 U1145 ( .A(KEYINPUT15), .ZN(n1306) );
endmodule


