//Key = 0010000001101110111011111010000000001010011010110110011011001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305;

XNOR2_X1 U721 ( .A(G107), .B(n991), .ZN(G9) );
NOR2_X1 U722 ( .A1(n992), .A2(KEYINPUT8), .ZN(n991) );
NOR2_X1 U723 ( .A1(n993), .A2(n994), .ZN(G75) );
NOR4_X1 U724 ( .A1(n995), .A2(n996), .A3(G953), .A4(n997), .ZN(n994) );
NOR2_X1 U725 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR2_X1 U726 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NOR2_X1 U727 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U728 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR2_X1 U729 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U732 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U733 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1008) );
NOR2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR3_X1 U736 ( .A1(n1017), .A2(n1020), .A3(n1011), .ZN(n1004) );
NOR2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR4_X1 U739 ( .A1(n1025), .A2(n1011), .A3(n1007), .A4(n1017), .ZN(n1000) );
NOR2_X1 U740 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND3_X1 U741 ( .A1(n1028), .A2(n1029), .A3(KEYINPUT41), .ZN(n995) );
XNOR2_X1 U742 ( .A(KEYINPUT1), .B(n1030), .ZN(n1029) );
NOR3_X1 U743 ( .A1(n997), .A2(G953), .A3(G952), .ZN(n993) );
AND4_X1 U744 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n997) );
NOR4_X1 U745 ( .A1(n1035), .A2(n1036), .A3(n1007), .A4(n1037), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1038), .B(n1039), .Z(n1036) );
NOR2_X1 U747 ( .A1(n1040), .A2(KEYINPUT15), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1035) );
XNOR2_X1 U749 ( .A(n1043), .B(KEYINPUT3), .ZN(n1042) );
INV_X1 U750 ( .A(n1044), .ZN(n1041) );
NOR3_X1 U751 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1033) );
NAND3_X1 U752 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1031) );
OR2_X1 U753 ( .A1(n1051), .A2(KEYINPUT9), .ZN(n1050) );
NAND3_X1 U754 ( .A1(KEYINPUT9), .A2(n1052), .A3(n1053), .ZN(n1049) );
INV_X1 U755 ( .A(n1054), .ZN(n1052) );
NAND2_X1 U756 ( .A1(G475), .A2(n1054), .ZN(n1048) );
NAND2_X1 U757 ( .A1(KEYINPUT24), .A2(n1051), .ZN(n1054) );
XOR2_X1 U758 ( .A(n1055), .B(KEYINPUT16), .Z(n1051) );
XOR2_X1 U759 ( .A(n1056), .B(n1057), .Z(G72) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NAND2_X1 U764 ( .A1(G953), .A2(n1063), .ZN(n1065) );
XOR2_X1 U765 ( .A(n1066), .B(n1067), .Z(n1064) );
XNOR2_X1 U766 ( .A(n1068), .B(KEYINPUT13), .ZN(n1067) );
NAND2_X1 U767 ( .A1(KEYINPUT10), .A2(n1069), .ZN(n1068) );
XOR2_X1 U768 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U769 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U770 ( .A1(G137), .A2(KEYINPUT25), .ZN(n1073) );
XOR2_X1 U771 ( .A(G131), .B(n1074), .Z(n1070) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
XOR2_X1 U773 ( .A(n1077), .B(KEYINPUT60), .Z(n1076) );
NAND2_X1 U774 ( .A1(G125), .A2(n1078), .ZN(n1077) );
NOR2_X1 U775 ( .A1(G125), .A2(n1078), .ZN(n1075) );
NAND2_X1 U776 ( .A1(n1061), .A2(n1030), .ZN(n1056) );
XOR2_X1 U777 ( .A(n1079), .B(n1080), .Z(G69) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U780 ( .A(KEYINPUT35), .B(n1085), .Z(n1084) );
NOR2_X1 U781 ( .A1(n1028), .A2(G953), .ZN(n1085) );
XNOR2_X1 U782 ( .A(n1086), .B(KEYINPUT51), .ZN(n1083) );
NOR3_X1 U783 ( .A1(n1086), .A2(G953), .A3(n1028), .ZN(n1081) );
INV_X1 U784 ( .A(n1087), .ZN(n1028) );
AND3_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1086) );
XOR2_X1 U786 ( .A(n1091), .B(KEYINPUT11), .Z(n1090) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U789 ( .A(n1096), .B(G122), .Z(n1092) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1089) );
XOR2_X1 U791 ( .A(G122), .B(G110), .Z(n1098) );
XOR2_X1 U792 ( .A(n1099), .B(n1094), .Z(n1097) );
NOR2_X1 U793 ( .A1(KEYINPUT48), .A2(n1100), .ZN(n1094) );
NAND2_X1 U794 ( .A1(G953), .A2(n1101), .ZN(n1088) );
NAND2_X1 U795 ( .A1(n1102), .A2(G953), .ZN(n1079) );
XOR2_X1 U796 ( .A(n1103), .B(KEYINPUT62), .Z(n1102) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1103) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U799 ( .A(KEYINPUT37), .B(n1106), .Z(n1105) );
NOR2_X1 U800 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
XOR2_X1 U801 ( .A(n1109), .B(KEYINPUT5), .Z(n1108) );
NAND2_X1 U802 ( .A1(n1038), .A2(n1110), .ZN(n1109) );
NAND2_X1 U803 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U804 ( .A1(n1040), .A2(n1113), .ZN(n1112) );
NOR3_X1 U805 ( .A1(n1114), .A2(n1111), .A3(n1115), .ZN(n1107) );
NOR2_X1 U806 ( .A1(n1106), .A2(n1116), .ZN(G63) );
XNOR2_X1 U807 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND3_X1 U808 ( .A1(G478), .A2(n1113), .A3(n1119), .ZN(n1117) );
XOR2_X1 U809 ( .A(n1120), .B(KEYINPUT53), .Z(n1119) );
NOR2_X1 U810 ( .A1(n1106), .A2(n1121), .ZN(G60) );
NOR3_X1 U811 ( .A1(n1055), .A2(n1122), .A3(n1123), .ZN(n1121) );
AND3_X1 U812 ( .A1(n1124), .A2(G475), .A3(n1125), .ZN(n1123) );
NOR2_X1 U813 ( .A1(n1126), .A2(n1124), .ZN(n1122) );
NOR2_X1 U814 ( .A1(n1127), .A2(n1053), .ZN(n1126) );
INV_X1 U815 ( .A(G475), .ZN(n1053) );
XOR2_X1 U816 ( .A(G104), .B(n1128), .Z(G6) );
NOR2_X1 U817 ( .A1(KEYINPUT29), .A2(n1129), .ZN(n1128) );
NOR3_X1 U818 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G57) );
NOR3_X1 U819 ( .A1(n1133), .A2(G953), .A3(G952), .ZN(n1132) );
AND2_X1 U820 ( .A1(n1133), .A2(n1106), .ZN(n1131) );
INV_X1 U821 ( .A(KEYINPUT39), .ZN(n1133) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(n1130) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1134) );
AND2_X1 U824 ( .A1(G472), .A2(n1125), .ZN(n1137) );
NAND2_X1 U825 ( .A1(n1138), .A2(KEYINPUT50), .ZN(n1136) );
XOR2_X1 U826 ( .A(n1139), .B(n1140), .Z(n1138) );
AND3_X1 U827 ( .A1(n1141), .A2(n1142), .A3(G210), .ZN(n1140) );
INV_X1 U828 ( .A(KEYINPUT32), .ZN(n1142) );
NOR2_X1 U829 ( .A1(n1106), .A2(n1143), .ZN(G54) );
XOR2_X1 U830 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U831 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1144) );
XNOR2_X1 U833 ( .A(n1150), .B(n1151), .ZN(n1148) );
NAND3_X1 U834 ( .A1(n1125), .A2(G469), .A3(KEYINPUT20), .ZN(n1151) );
INV_X1 U835 ( .A(n1114), .ZN(n1125) );
NAND2_X1 U836 ( .A1(KEYINPUT54), .A2(n1152), .ZN(n1150) );
XOR2_X1 U837 ( .A(KEYINPUT22), .B(G110), .Z(n1152) );
NOR2_X1 U838 ( .A1(n1106), .A2(n1153), .ZN(G51) );
XOR2_X1 U839 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U840 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
XOR2_X1 U841 ( .A(KEYINPUT43), .B(G210), .Z(n1158) );
NAND2_X1 U842 ( .A1(KEYINPUT17), .A2(n1114), .ZN(n1157) );
NAND2_X1 U843 ( .A1(G902), .A2(n1113), .ZN(n1114) );
INV_X1 U844 ( .A(n1127), .ZN(n1113) );
NAND2_X1 U845 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
INV_X1 U846 ( .A(KEYINPUT17), .ZN(n1160) );
NAND2_X1 U847 ( .A1(n1127), .A2(G902), .ZN(n1159) );
NOR2_X1 U848 ( .A1(n1087), .A2(n1030), .ZN(n1127) );
NAND4_X1 U849 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1030) );
NOR4_X1 U850 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
AND2_X1 U851 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
NAND3_X1 U852 ( .A1(n1013), .A2(n1027), .A3(n1171), .ZN(n1161) );
NAND2_X1 U853 ( .A1(n1172), .A2(n1173), .ZN(n1087) );
NOR4_X1 U854 ( .A1(n1174), .A2(n992), .A3(n1175), .A4(n1176), .ZN(n1173) );
AND3_X1 U855 ( .A1(n1026), .A2(n1177), .A3(n1178), .ZN(n992) );
AND4_X1 U856 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1129), .ZN(n1172) );
NAND3_X1 U857 ( .A1(n1178), .A2(n1177), .A3(n1027), .ZN(n1129) );
NOR2_X1 U858 ( .A1(n1061), .A2(G952), .ZN(n1106) );
XOR2_X1 U859 ( .A(G146), .B(n1182), .Z(G48) );
NOR3_X1 U860 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
XNOR2_X1 U861 ( .A(n1186), .B(KEYINPUT23), .ZN(n1184) );
XNOR2_X1 U862 ( .A(G143), .B(n1162), .ZN(G45) );
NAND4_X1 U863 ( .A1(n1013), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1162) );
XNOR2_X1 U864 ( .A(n1167), .B(n1190), .ZN(G42) );
XOR2_X1 U865 ( .A(n1078), .B(KEYINPUT63), .Z(n1190) );
AND4_X1 U866 ( .A1(n1191), .A2(n1027), .A3(n1192), .A4(n1018), .ZN(n1167) );
NOR2_X1 U867 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U868 ( .A(G137), .B(n1166), .Z(G39) );
NOR3_X1 U869 ( .A1(n1017), .A2(n1003), .A3(n1183), .ZN(n1166) );
INV_X1 U870 ( .A(n1191), .ZN(n1017) );
XOR2_X1 U871 ( .A(n1074), .B(n1170), .Z(G36) );
NAND3_X1 U872 ( .A1(n1191), .A2(n1026), .A3(n1187), .ZN(n1170) );
XOR2_X1 U873 ( .A(n1169), .B(n1195), .Z(G33) );
NOR2_X1 U874 ( .A1(G131), .A2(KEYINPUT30), .ZN(n1195) );
NAND3_X1 U875 ( .A1(n1191), .A2(n1027), .A3(n1187), .ZN(n1169) );
AND3_X1 U876 ( .A1(n1022), .A2(n1196), .A3(n1019), .ZN(n1187) );
NOR2_X1 U877 ( .A1(n1014), .A2(n1045), .ZN(n1191) );
INV_X1 U878 ( .A(n1015), .ZN(n1045) );
XOR2_X1 U879 ( .A(n1165), .B(n1197), .Z(G30) );
XOR2_X1 U880 ( .A(KEYINPUT45), .B(G128), .Z(n1197) );
AND3_X1 U881 ( .A1(n1013), .A2(n1026), .A3(n1171), .ZN(n1165) );
INV_X1 U882 ( .A(n1183), .ZN(n1171) );
NAND4_X1 U883 ( .A1(n1022), .A2(n1198), .A3(n1037), .A4(n1196), .ZN(n1183) );
INV_X1 U884 ( .A(n1194), .ZN(n1022) );
NAND2_X1 U885 ( .A1(n1199), .A2(n1200), .ZN(G3) );
NAND2_X1 U886 ( .A1(n1174), .A2(n1139), .ZN(n1200) );
XOR2_X1 U887 ( .A(KEYINPUT38), .B(n1201), .Z(n1199) );
NOR2_X1 U888 ( .A1(n1174), .A2(n1139), .ZN(n1201) );
AND3_X1 U889 ( .A1(n1019), .A2(n1178), .A3(n1202), .ZN(n1174) );
XOR2_X1 U890 ( .A(G125), .B(n1168), .Z(G27) );
AND4_X1 U891 ( .A1(n1013), .A2(n1027), .A3(n1203), .A4(n1018), .ZN(n1168) );
NOR2_X1 U892 ( .A1(n1193), .A2(n1007), .ZN(n1203) );
INV_X1 U893 ( .A(n1196), .ZN(n1193) );
NAND2_X1 U894 ( .A1(n1204), .A2(n1205), .ZN(n1196) );
NAND2_X1 U895 ( .A1(n1206), .A2(n1063), .ZN(n1205) );
INV_X1 U896 ( .A(G900), .ZN(n1063) );
XOR2_X1 U897 ( .A(n1181), .B(n1207), .Z(G24) );
XOR2_X1 U898 ( .A(KEYINPUT42), .B(G122), .Z(n1207) );
NAND4_X1 U899 ( .A1(n1208), .A2(n1177), .A3(n1188), .A4(n1189), .ZN(n1181) );
INV_X1 U900 ( .A(n1011), .ZN(n1177) );
NAND2_X1 U901 ( .A1(n1209), .A2(n1210), .ZN(n1011) );
XNOR2_X1 U902 ( .A(G119), .B(n1180), .ZN(G21) );
NAND4_X1 U903 ( .A1(n1208), .A2(n1202), .A3(n1198), .A4(n1037), .ZN(n1180) );
XOR2_X1 U904 ( .A(n1211), .B(n1179), .Z(G18) );
NAND3_X1 U905 ( .A1(n1019), .A2(n1026), .A3(n1208), .ZN(n1179) );
NOR3_X1 U906 ( .A1(n1007), .A2(n1212), .A3(n1186), .ZN(n1208) );
INV_X1 U907 ( .A(n1013), .ZN(n1186) );
XOR2_X1 U908 ( .A(n1213), .B(KEYINPUT44), .Z(n1013) );
AND2_X1 U909 ( .A1(n1214), .A2(n1189), .ZN(n1026) );
XNOR2_X1 U910 ( .A(n1176), .B(n1215), .ZN(G15) );
XNOR2_X1 U911 ( .A(G113), .B(KEYINPUT28), .ZN(n1215) );
AND3_X1 U912 ( .A1(n1027), .A2(n1019), .A3(n1216), .ZN(n1176) );
NOR3_X1 U913 ( .A1(n1007), .A2(n1212), .A3(n1213), .ZN(n1216) );
NAND2_X1 U914 ( .A1(n1217), .A2(n1024), .ZN(n1007) );
INV_X1 U915 ( .A(n1023), .ZN(n1217) );
AND2_X1 U916 ( .A1(n1037), .A2(n1210), .ZN(n1019) );
XNOR2_X1 U917 ( .A(n1218), .B(KEYINPUT26), .ZN(n1210) );
INV_X1 U918 ( .A(n1209), .ZN(n1037) );
INV_X1 U919 ( .A(n1185), .ZN(n1027) );
NAND2_X1 U920 ( .A1(n1219), .A2(n1188), .ZN(n1185) );
XOR2_X1 U921 ( .A(G110), .B(n1175), .Z(G12) );
AND3_X1 U922 ( .A1(n1202), .A2(n1178), .A3(n1018), .ZN(n1175) );
AND2_X1 U923 ( .A1(n1209), .A2(n1198), .ZN(n1018) );
XNOR2_X1 U924 ( .A(n1218), .B(KEYINPUT34), .ZN(n1198) );
XOR2_X1 U925 ( .A(n1220), .B(n1040), .Z(n1218) );
INV_X1 U926 ( .A(n1115), .ZN(n1040) );
NAND2_X1 U927 ( .A1(G217), .A2(n1221), .ZN(n1115) );
XOR2_X1 U928 ( .A(n1038), .B(KEYINPUT55), .Z(n1220) );
NAND2_X1 U929 ( .A1(n1111), .A2(n1120), .ZN(n1038) );
XOR2_X1 U930 ( .A(n1222), .B(n1223), .Z(n1111) );
XOR2_X1 U931 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U932 ( .A(n1226), .B(n1227), .Z(n1225) );
INV_X1 U933 ( .A(n1149), .ZN(n1224) );
XOR2_X1 U934 ( .A(n1228), .B(n1229), .Z(n1222) );
XOR2_X1 U935 ( .A(KEYINPUT12), .B(G137), .Z(n1229) );
XOR2_X1 U936 ( .A(n1230), .B(G128), .Z(n1228) );
NAND3_X1 U937 ( .A1(G221), .A2(n1061), .A3(n1231), .ZN(n1230) );
XOR2_X1 U938 ( .A(n1232), .B(KEYINPUT21), .Z(n1231) );
XOR2_X1 U939 ( .A(n1233), .B(G472), .Z(n1209) );
NAND3_X1 U940 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
XOR2_X1 U941 ( .A(n1120), .B(KEYINPUT19), .Z(n1236) );
NAND2_X1 U942 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
NAND2_X1 U943 ( .A1(n1141), .A2(G210), .ZN(n1238) );
XNOR2_X1 U944 ( .A(n1239), .B(n1135), .ZN(n1237) );
NAND2_X1 U945 ( .A1(KEYINPUT57), .A2(G101), .ZN(n1239) );
NAND3_X1 U946 ( .A1(G210), .A2(n1240), .A3(n1141), .ZN(n1234) );
XNOR2_X1 U947 ( .A(n1241), .B(n1135), .ZN(n1240) );
XNOR2_X1 U948 ( .A(n1242), .B(n1243), .ZN(n1135) );
XOR2_X1 U949 ( .A(G113), .B(n1244), .Z(n1243) );
XOR2_X1 U950 ( .A(KEYINPUT58), .B(G116), .Z(n1244) );
XOR2_X1 U951 ( .A(n1245), .B(n1246), .Z(n1242) );
INV_X1 U952 ( .A(n1247), .ZN(n1246) );
XOR2_X1 U953 ( .A(n1248), .B(n1249), .Z(n1245) );
INV_X1 U954 ( .A(n1226), .ZN(n1249) );
NAND2_X1 U955 ( .A1(n1250), .A2(KEYINPUT57), .ZN(n1241) );
XOR2_X1 U956 ( .A(n1139), .B(KEYINPUT52), .Z(n1250) );
INV_X1 U957 ( .A(G101), .ZN(n1139) );
NOR3_X1 U958 ( .A1(n1213), .A2(n1212), .A3(n1194), .ZN(n1178) );
NAND2_X1 U959 ( .A1(n1023), .A2(n1024), .ZN(n1194) );
NAND2_X1 U960 ( .A1(G221), .A2(n1221), .ZN(n1024) );
NAND2_X1 U961 ( .A1(G234), .A2(n1120), .ZN(n1221) );
XNOR2_X1 U962 ( .A(n1251), .B(G469), .ZN(n1023) );
NAND2_X1 U963 ( .A1(n1252), .A2(n1120), .ZN(n1251) );
XOR2_X1 U964 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U965 ( .A(n1146), .B(n1255), .Z(n1254) );
NOR2_X1 U966 ( .A1(KEYINPUT31), .A2(n1096), .ZN(n1255) );
INV_X1 U967 ( .A(G110), .ZN(n1096) );
XOR2_X1 U968 ( .A(n1256), .B(n1257), .Z(n1146) );
XOR2_X1 U969 ( .A(n1258), .B(n1247), .Z(n1257) );
XOR2_X1 U970 ( .A(n1259), .B(n1260), .Z(n1247) );
XOR2_X1 U971 ( .A(G137), .B(G134), .Z(n1260) );
NAND2_X1 U972 ( .A1(KEYINPUT2), .A2(G131), .ZN(n1259) );
NAND2_X1 U973 ( .A1(KEYINPUT49), .A2(n1261), .ZN(n1258) );
XOR2_X1 U974 ( .A(n1262), .B(n1263), .Z(n1256) );
NOR2_X1 U975 ( .A1(G101), .A2(KEYINPUT27), .ZN(n1263) );
XNOR2_X1 U976 ( .A(G107), .B(n1264), .ZN(n1262) );
NOR2_X1 U977 ( .A1(G953), .A2(n1062), .ZN(n1264) );
INV_X1 U978 ( .A(G227), .ZN(n1062) );
XOR2_X1 U979 ( .A(n1078), .B(n1265), .Z(n1253) );
NOR2_X1 U980 ( .A1(KEYINPUT40), .A2(n1072), .ZN(n1265) );
XOR2_X1 U981 ( .A(n1266), .B(n1147), .Z(n1072) );
AND2_X1 U982 ( .A1(n1204), .A2(n1267), .ZN(n1212) );
NAND2_X1 U983 ( .A1(n1206), .A2(n1101), .ZN(n1267) );
INV_X1 U984 ( .A(G898), .ZN(n1101) );
NOR3_X1 U985 ( .A1(n1120), .A2(n998), .A3(n1061), .ZN(n1206) );
NAND3_X1 U986 ( .A1(G952), .A2(n1061), .A3(n1268), .ZN(n1204) );
XNOR2_X1 U987 ( .A(n998), .B(KEYINPUT0), .ZN(n1268) );
NOR2_X1 U988 ( .A1(n1269), .A2(n1232), .ZN(n998) );
NAND2_X1 U989 ( .A1(n1014), .A2(n1015), .ZN(n1213) );
NAND2_X1 U990 ( .A1(n1270), .A2(n1271), .ZN(n1015) );
XNOR2_X1 U991 ( .A(G214), .B(KEYINPUT46), .ZN(n1270) );
OR2_X1 U992 ( .A1(n1047), .A2(n1272), .ZN(n1014) );
AND2_X1 U993 ( .A1(n1043), .A2(n1044), .ZN(n1272) );
NOR2_X1 U994 ( .A1(n1044), .A2(n1043), .ZN(n1047) );
AND2_X1 U995 ( .A1(G210), .A2(n1271), .ZN(n1043) );
NAND2_X1 U996 ( .A1(n1269), .A2(n1120), .ZN(n1271) );
INV_X1 U997 ( .A(G237), .ZN(n1269) );
NAND2_X1 U998 ( .A1(n1155), .A2(n1120), .ZN(n1044) );
INV_X1 U999 ( .A(G902), .ZN(n1120) );
XOR2_X1 U1000 ( .A(n1273), .B(n1274), .Z(n1155) );
XOR2_X1 U1001 ( .A(n1227), .B(n1275), .Z(n1274) );
XOR2_X1 U1002 ( .A(G122), .B(n1276), .Z(n1275) );
AND2_X1 U1003 ( .A1(n1061), .A2(G224), .ZN(n1276) );
INV_X1 U1004 ( .A(G953), .ZN(n1061) );
XOR2_X1 U1005 ( .A(G125), .B(G110), .Z(n1227) );
XOR2_X1 U1006 ( .A(n1277), .B(n1095), .Z(n1273) );
INV_X1 U1007 ( .A(n1099), .ZN(n1095) );
XOR2_X1 U1008 ( .A(n1226), .B(n1278), .Z(n1099) );
XNOR2_X1 U1009 ( .A(n1279), .B(n1280), .ZN(n1278) );
NOR2_X1 U1010 ( .A1(G113), .A2(KEYINPUT59), .ZN(n1280) );
NAND2_X1 U1011 ( .A1(KEYINPUT61), .A2(n1211), .ZN(n1279) );
INV_X1 U1012 ( .A(G116), .ZN(n1211) );
XNOR2_X1 U1013 ( .A(G119), .B(KEYINPUT7), .ZN(n1226) );
XNOR2_X1 U1014 ( .A(n1248), .B(n1100), .ZN(n1277) );
XNOR2_X1 U1015 ( .A(G101), .B(n1281), .ZN(n1100) );
XOR2_X1 U1016 ( .A(G107), .B(G104), .Z(n1281) );
XOR2_X1 U1017 ( .A(n1282), .B(G128), .Z(n1248) );
NAND2_X1 U1018 ( .A1(n1283), .A2(KEYINPUT14), .ZN(n1282) );
XOR2_X1 U1019 ( .A(G143), .B(n1266), .Z(n1283) );
INV_X1 U1020 ( .A(G146), .ZN(n1266) );
INV_X1 U1021 ( .A(n1003), .ZN(n1202) );
NAND2_X1 U1022 ( .A1(n1219), .A2(n1214), .ZN(n1003) );
XOR2_X1 U1023 ( .A(KEYINPUT36), .B(n1188), .Z(n1214) );
XOR2_X1 U1024 ( .A(n1055), .B(G475), .Z(n1188) );
NOR2_X1 U1025 ( .A1(n1124), .A2(G902), .ZN(n1055) );
XNOR2_X1 U1026 ( .A(n1284), .B(n1285), .ZN(n1124) );
XOR2_X1 U1027 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U1028 ( .A(n1288), .B(n1149), .Z(n1287) );
XNOR2_X1 U1029 ( .A(n1078), .B(G146), .ZN(n1149) );
INV_X1 U1030 ( .A(G140), .ZN(n1078) );
NAND2_X1 U1031 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1288) );
XOR2_X1 U1032 ( .A(n1289), .B(n1290), .Z(n1286) );
NOR2_X1 U1033 ( .A1(KEYINPUT4), .A2(G125), .ZN(n1290) );
NAND2_X1 U1034 ( .A1(n1141), .A2(G214), .ZN(n1289) );
NOR2_X1 U1035 ( .A1(G953), .A2(G237), .ZN(n1141) );
XOR2_X1 U1036 ( .A(n1291), .B(n1292), .Z(n1284) );
XOR2_X1 U1037 ( .A(G131), .B(G122), .Z(n1292) );
XOR2_X1 U1038 ( .A(n1261), .B(G113), .Z(n1291) );
INV_X1 U1039 ( .A(G104), .ZN(n1261) );
INV_X1 U1040 ( .A(n1189), .ZN(n1219) );
NAND2_X1 U1041 ( .A1(n1293), .A2(n1032), .ZN(n1189) );
NAND2_X1 U1042 ( .A1(G478), .A2(n1294), .ZN(n1032) );
OR2_X1 U1043 ( .A1(n1118), .A2(G902), .ZN(n1294) );
XOR2_X1 U1044 ( .A(KEYINPUT18), .B(n1046), .Z(n1293) );
NOR3_X1 U1045 ( .A1(G478), .A2(G902), .A3(n1118), .ZN(n1046) );
XOR2_X1 U1046 ( .A(n1295), .B(n1296), .Z(n1118) );
XOR2_X1 U1047 ( .A(G107), .B(n1297), .Z(n1296) );
XOR2_X1 U1048 ( .A(G122), .B(G116), .Z(n1297) );
XOR2_X1 U1049 ( .A(n1298), .B(n1299), .Z(n1295) );
NOR3_X1 U1050 ( .A1(n1300), .A2(n1232), .A3(n1301), .ZN(n1299) );
INV_X1 U1051 ( .A(G217), .ZN(n1301) );
INV_X1 U1052 ( .A(G234), .ZN(n1232) );
XOR2_X1 U1053 ( .A(KEYINPUT6), .B(G953), .Z(n1300) );
NAND2_X1 U1054 ( .A1(n1302), .A2(n1303), .ZN(n1298) );
OR2_X1 U1055 ( .A1(n1304), .A2(n1074), .ZN(n1303) );
XOR2_X1 U1056 ( .A(n1305), .B(KEYINPUT33), .Z(n1302) );
NAND2_X1 U1057 ( .A1(n1304), .A2(n1074), .ZN(n1305) );
INV_X1 U1058 ( .A(G134), .ZN(n1074) );
XOR2_X1 U1059 ( .A(n1147), .B(KEYINPUT47), .Z(n1304) );
XOR2_X1 U1060 ( .A(G128), .B(G143), .Z(n1147) );
endmodule


