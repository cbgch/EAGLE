//Key = 1101101100011111000010000111011100000010010000101010010011110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U745 ( .A(n1035), .B(G107), .Z(G9) );
NAND2_X1 U746 ( .A1(KEYINPUT3), .A2(n1036), .ZN(n1035) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
XOR2_X1 U760 ( .A(KEYINPUT44), .B(n1064), .Z(n1063) );
NOR3_X1 U761 ( .A1(n1059), .A2(n1065), .A3(n1055), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U763 ( .A1(KEYINPUT28), .A2(n1068), .ZN(n1066) );
NOR4_X1 U764 ( .A1(n1069), .A2(n1055), .A3(n1059), .A4(n1051), .ZN(n1044) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
AND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1039) );
NAND3_X1 U768 ( .A1(n1077), .A2(n1078), .A3(KEYINPUT28), .ZN(n1076) );
OR4_X1 U769 ( .A1(n1043), .A2(n1059), .A3(n1068), .A4(n1055), .ZN(n1078) );
INV_X1 U770 ( .A(n1079), .ZN(n1055) );
NOR3_X1 U771 ( .A1(n1080), .A2(G953), .A3(G952), .ZN(n1037) );
INV_X1 U772 ( .A(n1074), .ZN(n1080) );
NAND4_X1 U773 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1074) );
NOR4_X1 U774 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
XOR2_X1 U775 ( .A(KEYINPUT62), .B(n1064), .Z(n1088) );
XOR2_X1 U776 ( .A(n1089), .B(n1090), .Z(n1086) );
NAND2_X1 U777 ( .A1(KEYINPUT63), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U778 ( .A(n1092), .B(n1093), .ZN(n1085) );
NOR2_X1 U779 ( .A1(G478), .A2(KEYINPUT60), .ZN(n1093) );
NOR3_X1 U780 ( .A1(n1073), .A2(n1094), .A3(n1095), .ZN(n1083) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1082) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(G72) );
XOR2_X1 U783 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U784 ( .A1(G953), .A2(n1102), .ZN(n1101) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U787 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U788 ( .A(n1106), .B(n1107), .Z(n1103) );
XOR2_X1 U789 ( .A(G125), .B(n1108), .Z(n1107) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
NOR2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U792 ( .A(KEYINPUT41), .B(n1113), .Z(n1112) );
NOR2_X1 U793 ( .A1(G134), .A2(n1113), .ZN(n1109) );
NOR2_X1 U794 ( .A1(n1114), .A2(G953), .ZN(n1098) );
NAND2_X1 U795 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND3_X1 U796 ( .A1(G953), .A2(n1117), .A3(n1118), .ZN(n1116) );
XOR2_X1 U797 ( .A(n1119), .B(KEYINPUT23), .Z(n1115) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U799 ( .A1(G953), .A2(n1117), .ZN(n1121) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1117) );
XOR2_X1 U801 ( .A(n1118), .B(n1122), .Z(n1120) );
AND2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1118) );
OR3_X1 U803 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
INV_X1 U804 ( .A(KEYINPUT12), .ZN(n1127) );
OR2_X1 U805 ( .A1(n1128), .A2(KEYINPUT6), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1126), .A2(n1125), .ZN(n1128) );
XNOR2_X1 U807 ( .A(n1129), .B(n1130), .ZN(n1125) );
XOR2_X1 U808 ( .A(KEYINPUT2), .B(n1131), .Z(n1130) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR3_X1 U811 ( .A1(n1136), .A2(KEYINPUT16), .A3(n1137), .ZN(n1135) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1138), .ZN(G63) );
NOR3_X1 U813 ( .A1(n1092), .A2(n1139), .A3(n1140), .ZN(n1138) );
NOR3_X1 U814 ( .A1(n1141), .A2(n1142), .A3(n1136), .ZN(n1140) );
INV_X1 U815 ( .A(n1143), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1144), .A2(n1143), .ZN(n1139) );
AND2_X1 U817 ( .A1(n1041), .A2(G478), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1132), .A2(n1145), .ZN(G60) );
XNOR2_X1 U819 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U820 ( .A(KEYINPUT55), .B(n1148), .Z(n1147) );
NOR2_X1 U821 ( .A1(n1149), .A2(n1136), .ZN(n1148) );
INV_X1 U822 ( .A(G475), .ZN(n1149) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(G6) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(G57) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U828 ( .A(KEYINPUT17), .B(n1160), .Z(n1159) );
AND2_X1 U829 ( .A1(n1158), .A2(n1160), .ZN(n1156) );
NOR2_X1 U830 ( .A1(n1136), .A2(n1091), .ZN(n1160) );
XNOR2_X1 U831 ( .A(n1161), .B(n1162), .ZN(n1158) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1161) );
NOR2_X1 U833 ( .A1(KEYINPUT10), .A2(n1165), .ZN(n1164) );
NOR2_X1 U834 ( .A1(G952), .A2(n1166), .ZN(n1152) );
XOR2_X1 U835 ( .A(n1075), .B(KEYINPUT36), .Z(n1166) );
NOR2_X1 U836 ( .A1(n1132), .A2(n1167), .ZN(G54) );
XOR2_X1 U837 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U838 ( .A(n1170), .B(n1108), .Z(n1169) );
XOR2_X1 U839 ( .A(n1171), .B(n1165), .Z(n1108) );
XOR2_X1 U840 ( .A(n1172), .B(n1162), .Z(n1170) );
NAND3_X1 U841 ( .A1(G469), .A2(n1041), .A3(n1173), .ZN(n1172) );
XOR2_X1 U842 ( .A(n1174), .B(KEYINPUT4), .Z(n1173) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1168) );
NOR2_X1 U844 ( .A1(KEYINPUT37), .A2(n1177), .ZN(n1176) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1175) );
NOR2_X1 U846 ( .A1(n1132), .A2(n1180), .ZN(G51) );
XNOR2_X1 U847 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1136), .ZN(n1181) );
NAND2_X1 U849 ( .A1(G902), .A2(n1041), .ZN(n1136) );
NAND2_X1 U850 ( .A1(n1114), .A2(n1122), .ZN(n1041) );
AND4_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1122) );
NOR4_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
AND2_X1 U853 ( .A1(n1071), .A2(n1192), .ZN(n1191) );
NOR4_X1 U854 ( .A1(n1068), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1190) );
XOR2_X1 U855 ( .A(KEYINPUT33), .B(n1196), .Z(n1195) );
INV_X1 U856 ( .A(n1151), .ZN(n1189) );
NAND3_X1 U857 ( .A1(n1197), .A2(n1198), .A3(n1067), .ZN(n1151) );
AND2_X1 U858 ( .A1(n1036), .A2(n1199), .ZN(n1186) );
NAND3_X1 U859 ( .A1(n1198), .A2(n1200), .A3(n1197), .ZN(n1036) );
INV_X1 U860 ( .A(n1059), .ZN(n1198) );
AND4_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1114) );
NOR4_X1 U862 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NOR3_X1 U863 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1203) );
AND2_X1 U864 ( .A1(KEYINPUT59), .A2(n1212), .ZN(n1211) );
NOR3_X1 U865 ( .A1(KEYINPUT59), .A2(n1057), .A3(n1213), .ZN(n1210) );
NOR3_X1 U866 ( .A1(n1051), .A2(n1214), .A3(n1047), .ZN(n1209) );
OR3_X1 U867 ( .A1(n1196), .A2(n1215), .A3(n1216), .ZN(n1201) );
NOR2_X1 U868 ( .A1(n1075), .A2(G952), .ZN(n1132) );
XNOR2_X1 U869 ( .A(G146), .B(n1202), .ZN(G48) );
OR3_X1 U870 ( .A1(n1196), .A2(n1214), .A3(n1217), .ZN(n1202) );
XOR2_X1 U871 ( .A(n1218), .B(n1219), .Z(G45) );
NOR3_X1 U872 ( .A1(n1220), .A2(n1215), .A3(n1216), .ZN(n1219) );
XOR2_X1 U873 ( .A(KEYINPUT51), .B(n1196), .Z(n1220) );
NAND2_X1 U874 ( .A1(KEYINPUT58), .A2(n1221), .ZN(n1218) );
XOR2_X1 U875 ( .A(n1208), .B(n1222), .Z(G42) );
NOR2_X1 U876 ( .A1(KEYINPUT21), .A2(n1223), .ZN(n1222) );
AND4_X1 U877 ( .A1(n1061), .A2(n1224), .A3(n1077), .A4(n1225), .ZN(n1208) );
NOR2_X1 U878 ( .A1(n1217), .A2(n1226), .ZN(n1225) );
XOR2_X1 U879 ( .A(n1227), .B(n1228), .Z(G39) );
NOR2_X1 U880 ( .A1(KEYINPUT5), .A2(n1229), .ZN(n1228) );
NOR3_X1 U881 ( .A1(n1230), .A2(n1214), .A3(n1051), .ZN(n1227) );
INV_X1 U882 ( .A(n1231), .ZN(n1051) );
XOR2_X1 U883 ( .A(KEYINPUT14), .B(n1077), .Z(n1230) );
INV_X1 U884 ( .A(n1047), .ZN(n1077) );
XOR2_X1 U885 ( .A(n1207), .B(n1232), .Z(G36) );
NOR2_X1 U886 ( .A1(KEYINPUT24), .A2(n1111), .ZN(n1232) );
NOR3_X1 U887 ( .A1(n1215), .A2(n1068), .A3(n1047), .ZN(n1207) );
XOR2_X1 U888 ( .A(n1206), .B(n1233), .Z(G33) );
NOR2_X1 U889 ( .A1(KEYINPUT40), .A2(n1234), .ZN(n1233) );
NOR3_X1 U890 ( .A1(n1047), .A2(n1215), .A3(n1217), .ZN(n1206) );
INV_X1 U891 ( .A(n1067), .ZN(n1217) );
NAND3_X1 U892 ( .A1(n1061), .A2(n1224), .A3(n1056), .ZN(n1215) );
NAND2_X1 U893 ( .A1(n1072), .A2(n1235), .ZN(n1047) );
XOR2_X1 U894 ( .A(G128), .B(n1205), .Z(G30) );
NOR3_X1 U895 ( .A1(n1196), .A2(n1068), .A3(n1214), .ZN(n1205) );
NAND4_X1 U896 ( .A1(n1061), .A2(n1236), .A3(n1087), .A4(n1224), .ZN(n1214) );
XOR2_X1 U897 ( .A(G101), .B(n1188), .Z(G3) );
AND3_X1 U898 ( .A1(n1056), .A2(n1197), .A3(n1231), .ZN(n1188) );
XOR2_X1 U899 ( .A(G125), .B(n1212), .Z(G27) );
NOR2_X1 U900 ( .A1(n1213), .A2(n1226), .ZN(n1212) );
NAND4_X1 U901 ( .A1(n1071), .A2(n1067), .A3(n1079), .A4(n1224), .ZN(n1213) );
NAND2_X1 U902 ( .A1(n1043), .A2(n1237), .ZN(n1224) );
NAND4_X1 U903 ( .A1(n1238), .A2(G902), .A3(n1239), .A4(n1105), .ZN(n1237) );
INV_X1 U904 ( .A(G900), .ZN(n1105) );
XOR2_X1 U905 ( .A(n1075), .B(KEYINPUT7), .Z(n1238) );
XOR2_X1 U906 ( .A(n1240), .B(n1241), .Z(G24) );
NAND2_X1 U907 ( .A1(KEYINPUT0), .A2(G122), .ZN(n1241) );
NAND2_X1 U908 ( .A1(n1071), .A2(n1242), .ZN(n1240) );
XOR2_X1 U909 ( .A(KEYINPUT32), .B(n1192), .Z(n1242) );
NOR3_X1 U910 ( .A1(n1216), .A2(n1059), .A3(n1194), .ZN(n1192) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1244), .ZN(n1059) );
NAND2_X1 U912 ( .A1(n1245), .A2(n1246), .ZN(n1216) );
XNOR2_X1 U913 ( .A(G119), .B(n1184), .ZN(G21) );
NAND3_X1 U914 ( .A1(n1247), .A2(n1231), .A3(n1248), .ZN(n1184) );
NOR3_X1 U915 ( .A1(n1196), .A2(n1243), .A3(n1249), .ZN(n1248) );
INV_X1 U916 ( .A(n1071), .ZN(n1196) );
XOR2_X1 U917 ( .A(n1250), .B(n1251), .Z(G18) );
NAND4_X1 U918 ( .A1(n1071), .A2(n1247), .A3(n1200), .A4(n1252), .ZN(n1251) );
XOR2_X1 U919 ( .A(KEYINPUT45), .B(n1056), .Z(n1252) );
INV_X1 U920 ( .A(n1068), .ZN(n1200) );
NAND2_X1 U921 ( .A1(n1246), .A2(n1081), .ZN(n1068) );
XNOR2_X1 U922 ( .A(n1253), .B(KEYINPUT1), .ZN(n1071) );
XOR2_X1 U923 ( .A(n1254), .B(n1185), .Z(G15) );
NAND4_X1 U924 ( .A1(n1247), .A2(n1067), .A3(n1056), .A4(n1253), .ZN(n1185) );
INV_X1 U925 ( .A(n1193), .ZN(n1056) );
NAND2_X1 U926 ( .A1(n1243), .A2(n1236), .ZN(n1193) );
INV_X1 U927 ( .A(n1249), .ZN(n1236) );
XOR2_X1 U928 ( .A(n1255), .B(KEYINPUT31), .Z(n1249) );
NOR2_X1 U929 ( .A1(n1081), .A2(n1246), .ZN(n1067) );
INV_X1 U930 ( .A(n1245), .ZN(n1081) );
INV_X1 U931 ( .A(n1194), .ZN(n1247) );
NAND2_X1 U932 ( .A1(n1079), .A2(n1256), .ZN(n1194) );
NAND2_X1 U933 ( .A1(n1257), .A2(n1258), .ZN(n1079) );
OR3_X1 U934 ( .A1(n1064), .A2(n1095), .A3(KEYINPUT44), .ZN(n1258) );
INV_X1 U935 ( .A(n1062), .ZN(n1095) );
NAND2_X1 U936 ( .A1(KEYINPUT44), .A2(n1061), .ZN(n1257) );
XOR2_X1 U937 ( .A(n1178), .B(n1199), .Z(G12) );
NAND3_X1 U938 ( .A1(n1057), .A2(n1197), .A3(n1231), .ZN(n1199) );
NOR2_X1 U939 ( .A1(n1245), .A2(n1246), .ZN(n1231) );
XNOR2_X1 U940 ( .A(n1092), .B(n1259), .ZN(n1246) );
NOR2_X1 U941 ( .A1(KEYINPUT39), .A2(n1260), .ZN(n1259) );
XOR2_X1 U942 ( .A(n1142), .B(KEYINPUT26), .Z(n1260) );
INV_X1 U943 ( .A(G478), .ZN(n1142) );
NOR2_X1 U944 ( .A1(n1143), .A2(G902), .ZN(n1092) );
XOR2_X1 U945 ( .A(n1261), .B(n1262), .Z(n1143) );
XOR2_X1 U946 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U947 ( .A(n1265), .B(n1266), .Z(n1264) );
NOR2_X1 U948 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U949 ( .A(n1269), .B(KEYINPUT30), .Z(n1268) );
NAND2_X1 U950 ( .A1(G122), .A2(n1250), .ZN(n1269) );
NOR2_X1 U951 ( .A1(G122), .A2(n1250), .ZN(n1267) );
INV_X1 U952 ( .A(G116), .ZN(n1250) );
NAND2_X1 U953 ( .A1(KEYINPUT15), .A2(n1221), .ZN(n1265) );
INV_X1 U954 ( .A(G143), .ZN(n1221) );
NAND2_X1 U955 ( .A1(n1270), .A2(G217), .ZN(n1263) );
XOR2_X1 U956 ( .A(n1271), .B(n1272), .Z(n1261) );
XOR2_X1 U957 ( .A(KEYINPUT22), .B(G134), .Z(n1272) );
XOR2_X1 U958 ( .A(n1273), .B(G128), .Z(n1271) );
XOR2_X1 U959 ( .A(n1274), .B(n1275), .Z(n1245) );
XOR2_X1 U960 ( .A(KEYINPUT25), .B(G475), .Z(n1275) );
NAND2_X1 U961 ( .A1(n1146), .A2(n1174), .ZN(n1274) );
XNOR2_X1 U962 ( .A(n1276), .B(n1277), .ZN(n1146) );
XOR2_X1 U963 ( .A(n1171), .B(n1278), .Z(n1277) );
INV_X1 U964 ( .A(n1279), .ZN(n1171) );
XOR2_X1 U965 ( .A(n1280), .B(n1281), .Z(n1276) );
XOR2_X1 U966 ( .A(G146), .B(G113), .Z(n1281) );
NAND3_X1 U967 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1280) );
OR2_X1 U968 ( .A1(n1285), .A2(n1234), .ZN(n1284) );
NAND2_X1 U969 ( .A1(KEYINPUT18), .A2(n1286), .ZN(n1283) );
NAND2_X1 U970 ( .A1(n1287), .A2(n1234), .ZN(n1286) );
XNOR2_X1 U971 ( .A(n1285), .B(KEYINPUT57), .ZN(n1287) );
NAND2_X1 U972 ( .A1(n1288), .A2(n1289), .ZN(n1282) );
INV_X1 U973 ( .A(KEYINPUT18), .ZN(n1289) );
NAND2_X1 U974 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
OR2_X1 U975 ( .A1(n1285), .A2(KEYINPUT57), .ZN(n1291) );
NAND3_X1 U976 ( .A1(n1285), .A2(n1234), .A3(KEYINPUT57), .ZN(n1290) );
INV_X1 U977 ( .A(G131), .ZN(n1234) );
XNOR2_X1 U978 ( .A(n1292), .B(G143), .ZN(n1285) );
NAND2_X1 U979 ( .A1(n1293), .A2(G214), .ZN(n1292) );
AND3_X1 U980 ( .A1(n1253), .A2(n1256), .A3(n1061), .ZN(n1197) );
AND2_X1 U981 ( .A1(n1064), .A2(n1062), .ZN(n1061) );
NAND2_X1 U982 ( .A1(G221), .A2(n1294), .ZN(n1062) );
XNOR2_X1 U983 ( .A(n1295), .B(G469), .ZN(n1064) );
NAND2_X1 U984 ( .A1(n1296), .A2(n1174), .ZN(n1295) );
XOR2_X1 U985 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U986 ( .A(n1179), .B(n1299), .Z(n1298) );
NOR3_X1 U987 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1299) );
AND2_X1 U988 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NOR3_X1 U989 ( .A1(n1304), .A2(n1305), .A3(n1303), .ZN(n1301) );
NOR2_X1 U990 ( .A1(n1306), .A2(n1162), .ZN(n1300) );
NOR2_X1 U991 ( .A1(n1307), .A2(n1303), .ZN(n1306) );
INV_X1 U992 ( .A(KEYINPUT27), .ZN(n1303) );
XOR2_X1 U993 ( .A(n1304), .B(KEYINPUT8), .Z(n1307) );
NAND3_X1 U994 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1304) );
OR2_X1 U995 ( .A1(n1165), .A2(n1311), .ZN(n1310) );
NAND2_X1 U996 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
INV_X1 U997 ( .A(KEYINPUT46), .ZN(n1313) );
NAND2_X1 U998 ( .A1(n1314), .A2(n1311), .ZN(n1312) );
XOR2_X1 U999 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U1000 ( .A1(KEYINPUT46), .A2(n1317), .ZN(n1308) );
NAND2_X1 U1001 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND3_X1 U1002 ( .A1(n1311), .A2(n1165), .A3(n1315), .ZN(n1319) );
INV_X1 U1003 ( .A(KEYINPUT43), .ZN(n1315) );
XNOR2_X1 U1004 ( .A(n1177), .B(KEYINPUT42), .ZN(n1311) );
XOR2_X1 U1005 ( .A(n1320), .B(n1321), .Z(n1177) );
XOR2_X1 U1006 ( .A(n1322), .B(n1323), .Z(n1321) );
NOR2_X1 U1007 ( .A1(KEYINPUT54), .A2(n1150), .ZN(n1322) );
INV_X1 U1008 ( .A(G104), .ZN(n1150) );
XOR2_X1 U1009 ( .A(n1273), .B(KEYINPUT13), .Z(n1320) );
INV_X1 U1010 ( .A(G107), .ZN(n1273) );
NAND2_X1 U1011 ( .A1(KEYINPUT43), .A2(n1316), .ZN(n1318) );
AND2_X1 U1012 ( .A1(G227), .A2(n1075), .ZN(n1179) );
NAND2_X1 U1013 ( .A1(KEYINPUT56), .A2(n1324), .ZN(n1297) );
XOR2_X1 U1014 ( .A(n1325), .B(n1279), .Z(n1324) );
NAND2_X1 U1015 ( .A1(KEYINPUT20), .A2(G110), .ZN(n1325) );
NAND2_X1 U1016 ( .A1(n1043), .A2(n1326), .ZN(n1256) );
NAND3_X1 U1017 ( .A1(n1126), .A2(n1239), .A3(G902), .ZN(n1326) );
NOR2_X1 U1018 ( .A1(n1075), .A2(G898), .ZN(n1126) );
NAND3_X1 U1019 ( .A1(n1239), .A2(n1075), .A3(G952), .ZN(n1043) );
NAND2_X1 U1020 ( .A1(G237), .A2(G234), .ZN(n1239) );
NOR2_X1 U1021 ( .A1(n1072), .A2(n1073), .ZN(n1253) );
INV_X1 U1022 ( .A(n1235), .ZN(n1073) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1327), .ZN(n1235) );
NOR2_X1 U1024 ( .A1(n1328), .A2(n1094), .ZN(n1072) );
AND3_X1 U1025 ( .A1(n1183), .A2(n1174), .A3(n1182), .ZN(n1094) );
AND2_X1 U1026 ( .A1(n1329), .A2(n1097), .ZN(n1328) );
NAND2_X1 U1027 ( .A1(n1182), .A2(n1174), .ZN(n1097) );
XOR2_X1 U1028 ( .A(n1330), .B(n1331), .Z(n1182) );
XOR2_X1 U1029 ( .A(n1278), .B(n1332), .Z(n1331) );
XOR2_X1 U1030 ( .A(KEYINPUT53), .B(n1333), .Z(n1332) );
AND2_X1 U1031 ( .A1(n1075), .A2(G224), .ZN(n1333) );
XOR2_X1 U1032 ( .A(G125), .B(n1131), .Z(n1278) );
XOR2_X1 U1033 ( .A(G104), .B(G122), .Z(n1131) );
XOR2_X1 U1034 ( .A(n1129), .B(n1165), .Z(n1330) );
INV_X1 U1035 ( .A(n1316), .ZN(n1165) );
XOR2_X1 U1036 ( .A(n1334), .B(n1335), .Z(n1129) );
XOR2_X1 U1037 ( .A(G107), .B(n1336), .Z(n1335) );
XOR2_X1 U1038 ( .A(KEYINPUT49), .B(G110), .Z(n1336) );
XOR2_X1 U1039 ( .A(n1337), .B(n1338), .Z(n1334) );
NOR2_X1 U1040 ( .A1(KEYINPUT9), .A2(n1323), .ZN(n1338) );
XOR2_X1 U1041 ( .A(KEYINPUT47), .B(n1096), .Z(n1329) );
INV_X1 U1042 ( .A(n1183), .ZN(n1096) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1327), .ZN(n1183) );
NAND2_X1 U1044 ( .A1(n1339), .A2(n1174), .ZN(n1327) );
INV_X1 U1045 ( .A(G237), .ZN(n1339) );
INV_X1 U1046 ( .A(n1226), .ZN(n1057) );
NAND2_X1 U1047 ( .A1(n1244), .A2(n1087), .ZN(n1226) );
INV_X1 U1048 ( .A(n1243), .ZN(n1087) );
XNOR2_X1 U1049 ( .A(n1340), .B(n1137), .ZN(n1243) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1294), .ZN(n1137) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1174), .ZN(n1294) );
NAND2_X1 U1052 ( .A1(n1134), .A2(n1174), .ZN(n1340) );
XNOR2_X1 U1053 ( .A(n1341), .B(n1342), .ZN(n1134) );
XOR2_X1 U1054 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1055 ( .A(n1345), .B(n1346), .Z(n1344) );
NAND2_X1 U1056 ( .A1(KEYINPUT38), .A2(G146), .ZN(n1346) );
NAND2_X1 U1057 ( .A1(n1270), .A2(G221), .ZN(n1345) );
AND2_X1 U1058 ( .A1(G234), .A2(n1075), .ZN(n1270) );
INV_X1 U1059 ( .A(G953), .ZN(n1075) );
NOR2_X1 U1060 ( .A1(KEYINPUT19), .A2(n1279), .ZN(n1343) );
XOR2_X1 U1061 ( .A(n1223), .B(KEYINPUT29), .Z(n1279) );
INV_X1 U1062 ( .A(G140), .ZN(n1223) );
XOR2_X1 U1063 ( .A(n1347), .B(n1348), .Z(n1341) );
XNOR2_X1 U1064 ( .A(G125), .B(n1349), .ZN(n1348) );
NAND2_X1 U1065 ( .A1(n1350), .A2(KEYINPUT50), .ZN(n1349) );
XOR2_X1 U1066 ( .A(n1178), .B(n1351), .Z(n1350) );
XOR2_X1 U1067 ( .A(G128), .B(G119), .Z(n1351) );
XOR2_X1 U1068 ( .A(n1229), .B(KEYINPUT35), .Z(n1347) );
INV_X1 U1069 ( .A(G137), .ZN(n1229) );
INV_X1 U1070 ( .A(n1255), .ZN(n1244) );
XOR2_X1 U1071 ( .A(n1091), .B(n1352), .Z(n1255) );
NOR2_X1 U1072 ( .A1(n1090), .A2(KEYINPUT34), .ZN(n1352) );
AND2_X1 U1073 ( .A1(n1353), .A2(n1174), .ZN(n1090) );
INV_X1 U1074 ( .A(G902), .ZN(n1174) );
XOR2_X1 U1075 ( .A(n1354), .B(n1355), .Z(n1353) );
XOR2_X1 U1076 ( .A(n1162), .B(n1155), .Z(n1355) );
XNOR2_X1 U1077 ( .A(n1356), .B(n1323), .ZN(n1155) );
XOR2_X1 U1078 ( .A(G101), .B(KEYINPUT48), .Z(n1323) );
NAND2_X1 U1079 ( .A1(n1293), .A2(G210), .ZN(n1356) );
NOR2_X1 U1080 ( .A1(G953), .A2(G237), .ZN(n1293) );
INV_X1 U1081 ( .A(n1305), .ZN(n1162) );
XOR2_X1 U1082 ( .A(n1111), .B(n1113), .Z(n1305) );
XOR2_X1 U1083 ( .A(G137), .B(G131), .Z(n1113) );
INV_X1 U1084 ( .A(G134), .ZN(n1111) );
XOR2_X1 U1085 ( .A(n1163), .B(n1357), .Z(n1354) );
XNOR2_X1 U1086 ( .A(n1358), .B(KEYINPUT52), .ZN(n1357) );
NAND2_X1 U1087 ( .A1(KEYINPUT61), .A2(n1316), .ZN(n1358) );
XOR2_X1 U1088 ( .A(n1359), .B(n1360), .Z(n1316) );
XOR2_X1 U1089 ( .A(G146), .B(G143), .Z(n1360) );
INV_X1 U1090 ( .A(G128), .ZN(n1359) );
XOR2_X1 U1091 ( .A(n1337), .B(KEYINPUT11), .Z(n1163) );
XOR2_X1 U1092 ( .A(n1254), .B(n1361), .Z(n1337) );
XOR2_X1 U1093 ( .A(G119), .B(G116), .Z(n1361) );
INV_X1 U1094 ( .A(G113), .ZN(n1254) );
INV_X1 U1095 ( .A(G472), .ZN(n1091) );
INV_X1 U1096 ( .A(G110), .ZN(n1178) );
endmodule


