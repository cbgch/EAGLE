//Key = 1101111010100011011101101110100100111100101000111110101110010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;

XNOR2_X1 U782 ( .A(n1083), .B(n1084), .ZN(G9) );
NOR2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(G75) );
NOR4_X1 U784 ( .A1(n1087), .A2(n1088), .A3(G953), .A4(n1089), .ZN(n1086) );
NOR3_X1 U785 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
NOR2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR3_X1 U787 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1093) );
NAND3_X1 U788 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1087) );
XNOR2_X1 U789 ( .A(n1101), .B(KEYINPUT19), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U792 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U794 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND3_X1 U801 ( .A1(n1119), .A2(n1115), .A3(n1125), .ZN(n1108) );
XOR2_X1 U802 ( .A(n1126), .B(KEYINPUT44), .Z(n1104) );
OR2_X1 U803 ( .A1(n1090), .A2(n1112), .ZN(n1126) );
NAND4_X1 U804 ( .A1(n1106), .A2(n1119), .A3(n1115), .A4(n1110), .ZN(n1090) );
INV_X1 U805 ( .A(n1127), .ZN(n1106) );
NOR3_X1 U806 ( .A1(n1089), .A2(G953), .A3(G952), .ZN(n1085) );
AND4_X1 U807 ( .A1(n1128), .A2(n1115), .A3(n1129), .A4(n1130), .ZN(n1089) );
NOR4_X1 U808 ( .A1(n1131), .A2(n1132), .A3(n1092), .A4(n1133), .ZN(n1130) );
XOR2_X1 U809 ( .A(n1134), .B(KEYINPUT43), .Z(n1132) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U811 ( .A(KEYINPUT25), .B(n1137), .ZN(n1135) );
XOR2_X1 U812 ( .A(n1138), .B(G478), .Z(n1129) );
NAND2_X1 U813 ( .A1(KEYINPUT59), .A2(n1139), .ZN(n1138) );
XNOR2_X1 U814 ( .A(n1140), .B(n1141), .ZN(n1128) );
NAND2_X1 U815 ( .A1(KEYINPUT1), .A2(n1142), .ZN(n1140) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(G72) );
XOR2_X1 U817 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND3_X1 U818 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
OR2_X1 U819 ( .A1(n1150), .A2(KEYINPUT45), .ZN(n1148) );
NAND2_X1 U820 ( .A1(n1151), .A2(KEYINPUT45), .ZN(n1147) );
NAND2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1145) );
NAND2_X1 U822 ( .A1(G953), .A2(n1154), .ZN(n1153) );
XOR2_X1 U823 ( .A(n1155), .B(n1156), .Z(n1152) );
XNOR2_X1 U824 ( .A(G140), .B(n1157), .ZN(n1156) );
NOR2_X1 U825 ( .A1(KEYINPUT51), .A2(n1158), .ZN(n1155) );
XNOR2_X1 U826 ( .A(n1159), .B(n1160), .ZN(n1158) );
XNOR2_X1 U827 ( .A(n1161), .B(n1162), .ZN(n1160) );
NAND2_X1 U828 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
NAND2_X1 U829 ( .A1(G137), .A2(n1165), .ZN(n1164) );
XOR2_X1 U830 ( .A(n1166), .B(KEYINPUT16), .Z(n1163) );
NAND2_X1 U831 ( .A1(G134), .A2(n1167), .ZN(n1166) );
NOR3_X1 U832 ( .A1(n1149), .A2(KEYINPUT32), .A3(n1168), .ZN(n1143) );
AND2_X1 U833 ( .A1(G227), .A2(G900), .ZN(n1168) );
XOR2_X1 U834 ( .A(n1169), .B(n1170), .Z(G69) );
XOR2_X1 U835 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U836 ( .A1(n1098), .A2(G953), .ZN(n1172) );
NAND3_X1 U837 ( .A1(KEYINPUT62), .A2(n1173), .A3(n1174), .ZN(n1171) );
NOR3_X1 U838 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
NAND2_X1 U839 ( .A1(n1178), .A2(n1179), .ZN(n1173) );
XOR2_X1 U840 ( .A(KEYINPUT42), .B(n1180), .Z(n1179) );
NAND2_X1 U841 ( .A1(G953), .A2(n1181), .ZN(n1169) );
NAND2_X1 U842 ( .A1(G898), .A2(G224), .ZN(n1181) );
NOR2_X1 U843 ( .A1(n1182), .A2(n1183), .ZN(G66) );
NOR2_X1 U844 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U845 ( .A(KEYINPUT58), .B(n1186), .Z(n1185) );
AND2_X1 U846 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U847 ( .A1(n1188), .A2(n1187), .ZN(n1184) );
NOR2_X1 U848 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR2_X1 U849 ( .A1(n1182), .A2(n1191), .ZN(G63) );
XOR2_X1 U850 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U851 ( .A1(KEYINPUT11), .A2(n1194), .ZN(n1193) );
NAND2_X1 U852 ( .A1(n1195), .A2(G478), .ZN(n1192) );
NOR2_X1 U853 ( .A1(n1182), .A2(n1196), .ZN(G60) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1196) );
AND2_X1 U855 ( .A1(G475), .A2(n1195), .ZN(n1198) );
NAND2_X1 U856 ( .A1(KEYINPUT46), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U857 ( .A(n1200), .B(n1201), .ZN(G6) );
NOR3_X1 U858 ( .A1(n1117), .A2(n1202), .A3(n1203), .ZN(n1201) );
XNOR2_X1 U859 ( .A(n1204), .B(KEYINPUT27), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1182), .A2(n1205), .ZN(G57) );
XOR2_X1 U861 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U862 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U863 ( .A(n1210), .B(n1211), .Z(n1206) );
XOR2_X1 U864 ( .A(KEYINPUT6), .B(n1212), .Z(n1211) );
NOR2_X1 U865 ( .A1(n1141), .A2(n1189), .ZN(n1212) );
INV_X1 U866 ( .A(G472), .ZN(n1141) );
NAND2_X1 U867 ( .A1(KEYINPUT48), .A2(n1213), .ZN(n1210) );
NOR3_X1 U868 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(G54) );
AND2_X1 U869 ( .A1(KEYINPUT55), .A2(n1182), .ZN(n1216) );
NOR3_X1 U870 ( .A1(KEYINPUT55), .A2(G952), .A3(n1217), .ZN(n1215) );
INV_X1 U871 ( .A(n1218), .ZN(n1217) );
XOR2_X1 U872 ( .A(n1219), .B(n1220), .Z(n1214) );
XNOR2_X1 U873 ( .A(n1221), .B(n1222), .ZN(n1220) );
NAND2_X1 U874 ( .A1(KEYINPUT3), .A2(n1223), .ZN(n1221) );
NAND2_X1 U875 ( .A1(n1195), .A2(G469), .ZN(n1223) );
INV_X1 U876 ( .A(n1189), .ZN(n1195) );
XOR2_X1 U877 ( .A(n1224), .B(n1225), .Z(n1219) );
NAND2_X1 U878 ( .A1(n1226), .A2(KEYINPUT54), .ZN(n1224) );
XOR2_X1 U879 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND2_X1 U880 ( .A1(KEYINPUT31), .A2(n1229), .ZN(n1227) );
NOR2_X1 U881 ( .A1(n1182), .A2(n1230), .ZN(G51) );
XOR2_X1 U882 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U883 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U884 ( .A1(n1235), .A2(n1189), .ZN(n1234) );
NAND2_X1 U885 ( .A1(G902), .A2(n1236), .ZN(n1189) );
NAND2_X1 U886 ( .A1(n1098), .A2(n1101), .ZN(n1236) );
INV_X1 U887 ( .A(n1150), .ZN(n1101) );
NAND2_X1 U888 ( .A1(n1237), .A2(n1238), .ZN(n1150) );
NOR4_X1 U889 ( .A1(n1151), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1238) );
NOR4_X1 U890 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1237) );
NOR2_X1 U891 ( .A1(n1118), .A2(n1246), .ZN(n1245) );
NOR2_X1 U892 ( .A1(n1117), .A2(n1246), .ZN(n1244) );
NOR3_X1 U893 ( .A1(n1247), .A2(n1248), .A3(n1110), .ZN(n1243) );
NAND3_X1 U894 ( .A1(n1249), .A2(n1092), .A3(n1250), .ZN(n1247) );
XNOR2_X1 U895 ( .A(KEYINPUT41), .B(n1121), .ZN(n1250) );
AND4_X1 U896 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1098) );
AND4_X1 U897 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
INV_X1 U898 ( .A(n1259), .ZN(n1257) );
NOR2_X1 U899 ( .A1(n1260), .A2(n1084), .ZN(n1253) );
NOR3_X1 U900 ( .A1(n1118), .A2(n1203), .A3(n1121), .ZN(n1084) );
NOR4_X1 U901 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1117), .ZN(n1260) );
XNOR2_X1 U902 ( .A(n1115), .B(KEYINPUT60), .ZN(n1261) );
NAND2_X1 U903 ( .A1(n1264), .A2(n1265), .ZN(n1252) );
XNOR2_X1 U904 ( .A(n1266), .B(KEYINPUT18), .ZN(n1264) );
OR3_X1 U905 ( .A1(n1121), .A2(n1203), .A3(n1117), .ZN(n1251) );
INV_X1 U906 ( .A(n1204), .ZN(n1121) );
NOR3_X1 U907 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1233) );
NOR2_X1 U908 ( .A1(n1270), .A2(n1157), .ZN(n1269) );
XNOR2_X1 U909 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR3_X1 U910 ( .A1(G125), .A2(n1273), .A3(n1274), .ZN(n1268) );
NOR2_X1 U911 ( .A1(n1271), .A2(n1275), .ZN(n1267) );
XNOR2_X1 U912 ( .A(n1276), .B(KEYINPUT7), .ZN(n1231) );
NOR2_X1 U913 ( .A1(n1218), .A2(G952), .ZN(n1182) );
XOR2_X1 U914 ( .A(n1149), .B(KEYINPUT57), .Z(n1218) );
XOR2_X1 U915 ( .A(G146), .B(n1242), .Z(G48) );
AND3_X1 U916 ( .A1(n1277), .A2(n1094), .A3(n1278), .ZN(n1242) );
XOR2_X1 U917 ( .A(G143), .B(n1241), .Z(G45) );
AND4_X1 U918 ( .A1(n1279), .A2(n1094), .A3(n1280), .A4(n1133), .ZN(n1241) );
XOR2_X1 U919 ( .A(G140), .B(n1240), .Z(G42) );
AND3_X1 U920 ( .A1(n1102), .A2(n1204), .A3(n1281), .ZN(n1240) );
XNOR2_X1 U921 ( .A(G137), .B(n1282), .ZN(G39) );
NAND2_X1 U922 ( .A1(n1283), .A2(n1278), .ZN(n1282) );
INV_X1 U923 ( .A(n1248), .ZN(n1283) );
NAND2_X1 U924 ( .A1(n1102), .A2(n1119), .ZN(n1248) );
XNOR2_X1 U925 ( .A(n1165), .B(n1284), .ZN(G36) );
NOR3_X1 U926 ( .A1(n1285), .A2(n1118), .A3(n1286), .ZN(n1284) );
XOR2_X1 U927 ( .A(KEYINPUT21), .B(n1102), .Z(n1285) );
NAND2_X1 U928 ( .A1(n1287), .A2(n1288), .ZN(G33) );
NAND2_X1 U929 ( .A1(n1162), .A2(n1289), .ZN(n1288) );
XOR2_X1 U930 ( .A(n1290), .B(n1291), .Z(n1287) );
NOR2_X1 U931 ( .A1(n1162), .A2(n1289), .ZN(n1291) );
INV_X1 U932 ( .A(KEYINPUT36), .ZN(n1289) );
NAND2_X1 U933 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
INV_X1 U934 ( .A(n1246), .ZN(n1293) );
NAND2_X1 U935 ( .A1(n1279), .A2(n1102), .ZN(n1246) );
NOR3_X1 U936 ( .A1(n1096), .A2(n1131), .A3(n1097), .ZN(n1102) );
INV_X1 U937 ( .A(n1136), .ZN(n1097) );
INV_X1 U938 ( .A(n1095), .ZN(n1131) );
INV_X1 U939 ( .A(n1137), .ZN(n1096) );
INV_X1 U940 ( .A(n1286), .ZN(n1279) );
NAND3_X1 U941 ( .A1(n1204), .A2(n1249), .A3(n1125), .ZN(n1286) );
XNOR2_X1 U942 ( .A(n1277), .B(KEYINPUT4), .ZN(n1292) );
XOR2_X1 U943 ( .A(G128), .B(n1239), .Z(G30) );
AND3_X1 U944 ( .A1(n1266), .A2(n1094), .A3(n1278), .ZN(n1239) );
AND4_X1 U945 ( .A1(n1294), .A2(n1204), .A3(n1249), .A4(n1092), .ZN(n1278) );
XNOR2_X1 U946 ( .A(G101), .B(n1258), .ZN(G3) );
NAND4_X1 U947 ( .A1(n1125), .A2(n1119), .A3(n1204), .A4(n1295), .ZN(n1258) );
XNOR2_X1 U948 ( .A(n1151), .B(n1296), .ZN(G27) );
NOR2_X1 U949 ( .A1(G125), .A2(KEYINPUT61), .ZN(n1296) );
AND3_X1 U950 ( .A1(n1115), .A2(n1094), .A3(n1281), .ZN(n1151) );
AND4_X1 U951 ( .A1(n1277), .A2(n1110), .A3(n1249), .A4(n1092), .ZN(n1281) );
NAND2_X1 U952 ( .A1(n1127), .A2(n1297), .ZN(n1249) );
NAND4_X1 U953 ( .A1(G902), .A2(G953), .A3(n1298), .A4(n1154), .ZN(n1297) );
INV_X1 U954 ( .A(G900), .ZN(n1154) );
NAND2_X1 U955 ( .A1(n1299), .A2(n1300), .ZN(G24) );
NAND2_X1 U956 ( .A1(n1259), .A2(n1301), .ZN(n1300) );
XOR2_X1 U957 ( .A(KEYINPUT26), .B(n1302), .Z(n1299) );
NOR2_X1 U958 ( .A1(n1259), .A2(n1301), .ZN(n1302) );
NOR4_X1 U959 ( .A1(n1303), .A2(n1203), .A3(n1304), .A4(n1305), .ZN(n1259) );
NAND3_X1 U960 ( .A1(n1295), .A2(n1110), .A3(n1112), .ZN(n1203) );
INV_X1 U961 ( .A(n1092), .ZN(n1112) );
XNOR2_X1 U962 ( .A(G119), .B(n1256), .ZN(G21) );
NAND3_X1 U963 ( .A1(n1306), .A2(n1115), .A3(n1294), .ZN(n1256) );
INV_X1 U964 ( .A(n1110), .ZN(n1294) );
INV_X1 U965 ( .A(n1303), .ZN(n1115) );
NAND2_X1 U966 ( .A1(n1307), .A2(n1308), .ZN(G18) );
NAND2_X1 U967 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U968 ( .A(KEYINPUT29), .B(n1311), .Z(n1309) );
NAND2_X1 U969 ( .A1(n1312), .A2(G116), .ZN(n1307) );
XOR2_X1 U970 ( .A(KEYINPUT22), .B(n1311), .Z(n1312) );
NOR2_X1 U971 ( .A1(n1313), .A2(n1118), .ZN(n1311) );
INV_X1 U972 ( .A(n1266), .ZN(n1118) );
NOR2_X1 U973 ( .A1(n1133), .A2(n1304), .ZN(n1266) );
XNOR2_X1 U974 ( .A(n1314), .B(n1315), .ZN(G15) );
NOR2_X1 U975 ( .A1(n1117), .A2(n1313), .ZN(n1315) );
INV_X1 U976 ( .A(n1265), .ZN(n1313) );
NOR3_X1 U977 ( .A1(n1303), .A2(n1262), .A3(n1263), .ZN(n1265) );
INV_X1 U978 ( .A(n1125), .ZN(n1263) );
NOR2_X1 U979 ( .A1(n1110), .A2(n1092), .ZN(n1125) );
NAND2_X1 U980 ( .A1(n1124), .A2(n1316), .ZN(n1303) );
INV_X1 U981 ( .A(n1277), .ZN(n1117) );
NOR2_X1 U982 ( .A1(n1280), .A2(n1305), .ZN(n1277) );
INV_X1 U983 ( .A(n1133), .ZN(n1305) );
XNOR2_X1 U984 ( .A(G110), .B(n1255), .ZN(G12) );
NAND3_X1 U985 ( .A1(n1204), .A2(n1110), .A3(n1306), .ZN(n1255) );
AND3_X1 U986 ( .A1(n1295), .A2(n1092), .A3(n1119), .ZN(n1306) );
NOR2_X1 U987 ( .A1(n1133), .A2(n1280), .ZN(n1119) );
INV_X1 U988 ( .A(n1304), .ZN(n1280) );
XOR2_X1 U989 ( .A(n1139), .B(n1317), .Z(n1304) );
XOR2_X1 U990 ( .A(KEYINPUT24), .B(G478), .Z(n1317) );
NOR2_X1 U991 ( .A1(n1194), .A2(G902), .ZN(n1139) );
XOR2_X1 U992 ( .A(n1318), .B(n1319), .Z(n1194) );
AND3_X1 U993 ( .A1(G217), .A2(n1320), .A3(G234), .ZN(n1319) );
NAND2_X1 U994 ( .A1(n1321), .A2(KEYINPUT50), .ZN(n1318) );
XOR2_X1 U995 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U996 ( .A(G128), .B(n1324), .Z(n1323) );
NOR2_X1 U997 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U998 ( .A(n1327), .B(KEYINPUT40), .Z(n1326) );
NAND2_X1 U999 ( .A1(n1328), .A2(n1083), .ZN(n1327) );
XOR2_X1 U1000 ( .A(KEYINPUT39), .B(n1329), .Z(n1328) );
NOR2_X1 U1001 ( .A1(n1083), .A2(n1329), .ZN(n1325) );
XNOR2_X1 U1002 ( .A(n1310), .B(n1330), .ZN(n1329) );
XNOR2_X1 U1003 ( .A(G134), .B(n1331), .ZN(n1322) );
XOR2_X1 U1004 ( .A(KEYINPUT28), .B(G143), .Z(n1331) );
XNOR2_X1 U1005 ( .A(n1332), .B(G475), .ZN(n1133) );
NAND2_X1 U1006 ( .A1(n1199), .A2(n1333), .ZN(n1332) );
XNOR2_X1 U1007 ( .A(n1334), .B(n1335), .ZN(n1199) );
XOR2_X1 U1008 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1009 ( .A(n1200), .B(n1338), .ZN(n1337) );
NOR2_X1 U1010 ( .A1(KEYINPUT38), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U1011 ( .A(n1340), .B(n1314), .ZN(n1339) );
INV_X1 U1012 ( .A(G113), .ZN(n1314) );
NAND2_X1 U1013 ( .A1(KEYINPUT17), .A2(n1330), .ZN(n1340) );
XNOR2_X1 U1014 ( .A(G140), .B(n1162), .ZN(n1336) );
INV_X1 U1015 ( .A(G131), .ZN(n1162) );
XOR2_X1 U1016 ( .A(n1341), .B(n1342), .Z(n1334) );
XOR2_X1 U1017 ( .A(n1343), .B(n1344), .Z(n1342) );
NOR2_X1 U1018 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
INV_X1 U1019 ( .A(G214), .ZN(n1346) );
NOR2_X1 U1020 ( .A1(KEYINPUT13), .A2(n1347), .ZN(n1343) );
XNOR2_X1 U1021 ( .A(G125), .B(KEYINPUT9), .ZN(n1347) );
XOR2_X1 U1022 ( .A(n1348), .B(n1349), .Z(n1341) );
NOR2_X1 U1023 ( .A1(G143), .A2(KEYINPUT63), .ZN(n1349) );
NAND2_X1 U1024 ( .A1(KEYINPUT56), .A2(G146), .ZN(n1348) );
NAND3_X1 U1025 ( .A1(n1350), .A2(n1351), .A3(n1352), .ZN(n1092) );
NAND2_X1 U1026 ( .A1(G902), .A2(G217), .ZN(n1352) );
OR3_X1 U1027 ( .A1(n1187), .A2(G902), .A3(n1353), .ZN(n1351) );
NAND2_X1 U1028 ( .A1(n1353), .A2(n1187), .ZN(n1350) );
XNOR2_X1 U1029 ( .A(n1354), .B(n1355), .ZN(n1187) );
XOR2_X1 U1030 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1031 ( .A(n1358), .B(n1359), .Z(n1357) );
NAND2_X1 U1032 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1033 ( .A1(n1362), .A2(n1167), .ZN(n1361) );
XOR2_X1 U1034 ( .A(KEYINPUT10), .B(n1363), .Z(n1360) );
NOR2_X1 U1035 ( .A1(n1167), .A2(n1362), .ZN(n1363) );
NAND3_X1 U1036 ( .A1(G234), .A2(n1320), .A3(G221), .ZN(n1362) );
NAND2_X1 U1037 ( .A1(n1364), .A2(KEYINPUT14), .ZN(n1358) );
XNOR2_X1 U1038 ( .A(G110), .B(n1365), .ZN(n1364) );
XOR2_X1 U1039 ( .A(G128), .B(G119), .Z(n1365) );
NOR2_X1 U1040 ( .A1(G140), .A2(KEYINPUT30), .ZN(n1356) );
XNOR2_X1 U1041 ( .A(G125), .B(n1366), .ZN(n1354) );
XOR2_X1 U1042 ( .A(KEYINPUT34), .B(G146), .Z(n1366) );
NOR2_X1 U1043 ( .A1(n1190), .A2(G234), .ZN(n1353) );
INV_X1 U1044 ( .A(G217), .ZN(n1190) );
INV_X1 U1045 ( .A(n1262), .ZN(n1295) );
NAND2_X1 U1046 ( .A1(n1094), .A2(n1367), .ZN(n1262) );
NAND2_X1 U1047 ( .A1(n1368), .A2(n1127), .ZN(n1367) );
NAND3_X1 U1048 ( .A1(n1298), .A2(n1149), .A3(G952), .ZN(n1127) );
NAND3_X1 U1049 ( .A1(G902), .A2(n1298), .A3(n1175), .ZN(n1368) );
NOR2_X1 U1050 ( .A1(n1149), .A2(G898), .ZN(n1175) );
INV_X1 U1051 ( .A(G953), .ZN(n1149) );
NAND2_X1 U1052 ( .A1(G237), .A2(G234), .ZN(n1298) );
AND2_X1 U1053 ( .A1(n1369), .A2(n1095), .ZN(n1094) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1370), .ZN(n1095) );
NAND2_X1 U1055 ( .A1(n1333), .A2(n1371), .ZN(n1370) );
NAND2_X1 U1056 ( .A1(n1137), .A2(n1136), .ZN(n1369) );
NAND2_X1 U1057 ( .A1(G210), .A2(n1372), .ZN(n1136) );
NAND2_X1 U1058 ( .A1(n1373), .A2(n1333), .ZN(n1372) );
NAND2_X1 U1059 ( .A1(n1374), .A2(G237), .ZN(n1373) );
XNOR2_X1 U1060 ( .A(n1276), .B(n1375), .ZN(n1374) );
NAND3_X1 U1061 ( .A1(n1376), .A2(n1333), .A3(n1377), .ZN(n1137) );
XOR2_X1 U1062 ( .A(n1375), .B(n1276), .Z(n1377) );
NOR3_X1 U1063 ( .A1(n1177), .A2(n1176), .A3(n1378), .ZN(n1276) );
NOR2_X1 U1064 ( .A1(n1379), .A2(n1180), .ZN(n1378) );
XNOR2_X1 U1065 ( .A(n1380), .B(n1381), .ZN(n1180) );
AND3_X1 U1066 ( .A1(n1380), .A2(n1379), .A3(n1381), .ZN(n1176) );
NOR3_X1 U1067 ( .A1(n1381), .A2(n1178), .A3(n1380), .ZN(n1177) );
XOR2_X1 U1068 ( .A(n1382), .B(n1383), .Z(n1380) );
NOR2_X1 U1069 ( .A1(G119), .A2(KEYINPUT20), .ZN(n1383) );
INV_X1 U1070 ( .A(n1379), .ZN(n1178) );
NAND3_X1 U1071 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n1379) );
NAND2_X1 U1072 ( .A1(n1387), .A2(n1083), .ZN(n1385) );
XNOR2_X1 U1073 ( .A(G104), .B(G101), .ZN(n1387) );
NAND3_X1 U1074 ( .A1(G104), .A2(n1388), .A3(G107), .ZN(n1384) );
XOR2_X1 U1075 ( .A(n1389), .B(G110), .Z(n1381) );
NAND2_X1 U1076 ( .A1(KEYINPUT8), .A2(n1330), .ZN(n1389) );
XNOR2_X1 U1077 ( .A(n1301), .B(KEYINPUT0), .ZN(n1330) );
INV_X1 U1078 ( .A(G122), .ZN(n1301) );
AND2_X1 U1079 ( .A1(n1390), .A2(n1391), .ZN(n1375) );
NAND2_X1 U1080 ( .A1(n1274), .A2(n1392), .ZN(n1391) );
NAND2_X1 U1081 ( .A1(n1275), .A2(n1393), .ZN(n1392) );
XOR2_X1 U1082 ( .A(KEYINPUT35), .B(n1394), .Z(n1390) );
AND3_X1 U1083 ( .A1(n1271), .A2(n1393), .A3(n1275), .ZN(n1394) );
NAND2_X1 U1084 ( .A1(n1273), .A2(n1157), .ZN(n1275) );
INV_X1 U1085 ( .A(G125), .ZN(n1157) );
NAND2_X1 U1086 ( .A1(n1395), .A2(n1272), .ZN(n1393) );
XNOR2_X1 U1087 ( .A(G125), .B(KEYINPUT15), .ZN(n1395) );
INV_X1 U1088 ( .A(n1274), .ZN(n1271) );
NAND2_X1 U1089 ( .A1(G224), .A2(n1320), .ZN(n1274) );
NAND2_X1 U1090 ( .A1(G210), .A2(G237), .ZN(n1376) );
XOR2_X1 U1091 ( .A(G472), .B(n1396), .Z(n1110) );
NOR2_X1 U1092 ( .A1(KEYINPUT23), .A2(n1142), .ZN(n1396) );
AND2_X1 U1093 ( .A1(n1397), .A2(n1333), .ZN(n1142) );
XOR2_X1 U1094 ( .A(n1398), .B(n1208), .Z(n1397) );
XNOR2_X1 U1095 ( .A(n1272), .B(n1228), .ZN(n1208) );
INV_X1 U1096 ( .A(n1273), .ZN(n1272) );
XNOR2_X1 U1097 ( .A(n1399), .B(n1400), .ZN(n1273) );
NAND2_X1 U1098 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1399) );
XNOR2_X1 U1099 ( .A(n1401), .B(n1402), .ZN(n1398) );
NOR2_X1 U1100 ( .A1(KEYINPUT53), .A2(n1209), .ZN(n1402) );
XNOR2_X1 U1101 ( .A(n1388), .B(n1403), .ZN(n1209) );
NOR2_X1 U1102 ( .A1(n1345), .A2(n1235), .ZN(n1403) );
INV_X1 U1103 ( .A(G210), .ZN(n1235) );
NAND2_X1 U1104 ( .A1(n1320), .A2(n1371), .ZN(n1345) );
INV_X1 U1105 ( .A(G237), .ZN(n1371) );
NOR2_X1 U1106 ( .A1(KEYINPUT33), .A2(n1213), .ZN(n1401) );
XOR2_X1 U1107 ( .A(G119), .B(n1382), .Z(n1213) );
XNOR2_X1 U1108 ( .A(G113), .B(n1310), .ZN(n1382) );
INV_X1 U1109 ( .A(G116), .ZN(n1310) );
NOR2_X1 U1110 ( .A1(n1124), .A2(n1123), .ZN(n1204) );
INV_X1 U1111 ( .A(n1316), .ZN(n1123) );
NAND2_X1 U1112 ( .A1(G221), .A2(n1404), .ZN(n1316) );
NAND2_X1 U1113 ( .A1(G234), .A2(n1333), .ZN(n1404) );
XOR2_X1 U1114 ( .A(n1405), .B(G469), .Z(n1124) );
NAND2_X1 U1115 ( .A1(n1406), .A2(n1333), .ZN(n1405) );
INV_X1 U1116 ( .A(G902), .ZN(n1333) );
XOR2_X1 U1117 ( .A(n1407), .B(n1408), .Z(n1406) );
XNOR2_X1 U1118 ( .A(n1229), .B(n1228), .ZN(n1408) );
XNOR2_X1 U1119 ( .A(n1409), .B(n1410), .ZN(n1228) );
XNOR2_X1 U1120 ( .A(n1167), .B(G131), .ZN(n1410) );
INV_X1 U1121 ( .A(G137), .ZN(n1167) );
NAND2_X1 U1122 ( .A1(KEYINPUT49), .A2(n1165), .ZN(n1409) );
INV_X1 U1123 ( .A(G134), .ZN(n1165) );
XOR2_X1 U1124 ( .A(n1411), .B(n1412), .Z(n1229) );
INV_X1 U1125 ( .A(n1159), .ZN(n1412) );
XNOR2_X1 U1126 ( .A(n1413), .B(n1400), .ZN(n1159) );
XOR2_X1 U1127 ( .A(G143), .B(G146), .Z(n1400) );
XNOR2_X1 U1128 ( .A(G128), .B(KEYINPUT5), .ZN(n1413) );
NAND3_X1 U1129 ( .A1(n1414), .A2(n1415), .A3(n1386), .ZN(n1411) );
NAND3_X1 U1130 ( .A1(G101), .A2(n1200), .A3(G107), .ZN(n1386) );
NAND2_X1 U1131 ( .A1(n1416), .A2(n1083), .ZN(n1415) );
INV_X1 U1132 ( .A(G107), .ZN(n1083) );
XNOR2_X1 U1133 ( .A(n1417), .B(G101), .ZN(n1416) );
NAND2_X1 U1134 ( .A1(n1418), .A2(G107), .ZN(n1414) );
NAND2_X1 U1135 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
NAND2_X1 U1136 ( .A1(n1417), .A2(n1388), .ZN(n1420) );
INV_X1 U1137 ( .A(G101), .ZN(n1388) );
NOR2_X1 U1138 ( .A1(n1200), .A2(KEYINPUT2), .ZN(n1417) );
INV_X1 U1139 ( .A(G104), .ZN(n1200) );
NAND2_X1 U1140 ( .A1(KEYINPUT2), .A2(G101), .ZN(n1419) );
XOR2_X1 U1141 ( .A(n1421), .B(n1225), .Z(n1407) );
AND2_X1 U1142 ( .A1(G227), .A2(n1320), .ZN(n1225) );
XOR2_X1 U1143 ( .A(G953), .B(KEYINPUT37), .Z(n1320) );
NAND2_X1 U1144 ( .A1(KEYINPUT47), .A2(n1222), .ZN(n1421) );
XOR2_X1 U1145 ( .A(G110), .B(n1422), .Z(n1222) );
XOR2_X1 U1146 ( .A(KEYINPUT12), .B(G140), .Z(n1422) );
endmodule


