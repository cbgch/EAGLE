//Key = 1000100011110001011100010101000011011111000000010100101100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359;

XNOR2_X1 U740 ( .A(G107), .B(n1025), .ZN(G9) );
NAND2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U743 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
INV_X1 U744 ( .A(n1033), .ZN(n1032) );
NOR2_X1 U745 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U748 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U753 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1053), .A2(n1052), .ZN(n1040) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U756 ( .A1(n1056), .A2(n1047), .A3(n1057), .ZN(n1054) );
NOR4_X1 U757 ( .A1(n1058), .A2(n1052), .A3(n1047), .A4(n1043), .ZN(n1036) );
INV_X1 U758 ( .A(n1059), .ZN(n1047) );
NOR3_X1 U759 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U760 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1030) );
NOR4_X1 U761 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XOR2_X1 U762 ( .A(n1068), .B(n1069), .Z(n1067) );
XNOR2_X1 U763 ( .A(KEYINPUT39), .B(n1070), .ZN(n1069) );
NOR4_X1 U764 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1062) );
AND3_X1 U765 ( .A1(KEYINPUT19), .A2(n1075), .A3(n1076), .ZN(n1074) );
NOR2_X1 U766 ( .A1(KEYINPUT19), .A2(n1076), .ZN(n1073) );
NOR2_X1 U767 ( .A1(KEYINPUT40), .A2(n1077), .ZN(n1072) );
NOR2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U769 ( .A1(KEYINPUT44), .A2(n1080), .ZN(n1079) );
AND2_X1 U770 ( .A1(n1081), .A2(KEYINPUT44), .ZN(n1078) );
NOR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1071) );
INV_X1 U772 ( .A(KEYINPUT40), .ZN(n1083) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
XNOR2_X1 U774 ( .A(KEYINPUT44), .B(n1086), .ZN(n1084) );
XNOR2_X1 U775 ( .A(n1087), .B(G475), .ZN(n1060) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND2_X1 U779 ( .A1(G227), .A2(G900), .ZN(n1092) );
NOR3_X1 U780 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1090) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U782 ( .A(n1099), .B(KEYINPUT52), .Z(n1094) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1099) );
NAND3_X1 U784 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
NAND2_X1 U785 ( .A1(KEYINPUT2), .A2(n1103), .ZN(n1102) );
NAND3_X1 U786 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1101) );
INV_X1 U787 ( .A(KEYINPUT2), .ZN(n1105) );
OR2_X1 U788 ( .A1(n1106), .A2(n1104), .ZN(n1100) );
NOR2_X1 U789 ( .A1(KEYINPUT28), .A2(n1103), .ZN(n1104) );
AND2_X1 U790 ( .A1(n1107), .A2(n1093), .ZN(n1088) );
XOR2_X1 U791 ( .A(n1108), .B(n1109), .Z(G69) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U793 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XNOR2_X1 U794 ( .A(KEYINPUT41), .B(n1093), .ZN(n1113) );
NOR2_X1 U795 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1116), .B(KEYINPUT30), .Z(n1114) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1110) );
XOR2_X1 U798 ( .A(n1119), .B(n1120), .Z(n1118) );
XNOR2_X1 U799 ( .A(n1121), .B(n1122), .ZN(n1120) );
XOR2_X1 U800 ( .A(n1123), .B(n1124), .Z(n1119) );
NAND2_X1 U801 ( .A1(KEYINPUT33), .A2(n1125), .ZN(n1123) );
NOR2_X1 U802 ( .A1(n1126), .A2(n1093), .ZN(n1108) );
AND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1126) );
NOR2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U806 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
XOR2_X1 U807 ( .A(KEYINPUT31), .B(G217), .Z(n1132) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1133), .ZN(G63) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U810 ( .A1(n1131), .A2(G478), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1136), .ZN(G60) );
NOR3_X1 U812 ( .A1(n1087), .A2(n1137), .A3(n1138), .ZN(n1136) );
NOR3_X1 U813 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NOR2_X1 U814 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1033), .A2(n1140), .ZN(n1142) );
XNOR2_X1 U816 ( .A(G104), .B(n1144), .ZN(G6) );
NAND2_X1 U817 ( .A1(n1145), .A2(n1027), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1127), .A2(n1146), .ZN(G57) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U820 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U821 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
XOR2_X1 U822 ( .A(n1153), .B(KEYINPUT4), .Z(n1152) );
NAND2_X1 U823 ( .A1(G101), .A2(n1154), .ZN(n1153) );
NOR2_X1 U824 ( .A1(G101), .A2(n1154), .ZN(n1151) );
XOR2_X1 U825 ( .A(KEYINPUT43), .B(n1155), .Z(n1154) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(n1147) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U828 ( .A(KEYINPUT50), .B(n1160), .Z(n1159) );
AND2_X1 U829 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1162), .A2(n1161), .ZN(n1158) );
NAND2_X1 U831 ( .A1(n1131), .A2(G472), .ZN(n1156) );
NOR2_X1 U832 ( .A1(n1127), .A2(n1163), .ZN(G54) );
XOR2_X1 U833 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U835 ( .A1(KEYINPUT13), .A2(n1168), .ZN(n1167) );
NAND3_X1 U836 ( .A1(n1169), .A2(n1170), .A3(G469), .ZN(n1166) );
NAND2_X1 U837 ( .A1(KEYINPUT61), .A2(n1141), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
INV_X1 U839 ( .A(KEYINPUT61), .ZN(n1172) );
NAND2_X1 U840 ( .A1(n1033), .A2(G902), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1173), .A2(n1174), .ZN(n1164) );
NAND2_X1 U842 ( .A1(G110), .A2(n1175), .ZN(n1174) );
NAND2_X1 U843 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
XNOR2_X1 U844 ( .A(KEYINPUT6), .B(n1175), .ZN(n1176) );
XNOR2_X1 U845 ( .A(n1178), .B(n1179), .ZN(n1175) );
NOR2_X1 U846 ( .A1(n1127), .A2(n1180), .ZN(G51) );
XOR2_X1 U847 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U848 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U849 ( .A1(KEYINPUT10), .A2(n1162), .ZN(n1184) );
OR2_X1 U850 ( .A1(n1141), .A2(n1075), .ZN(n1183) );
INV_X1 U851 ( .A(n1131), .ZN(n1141) );
NOR2_X1 U852 ( .A1(n1185), .A2(n1033), .ZN(n1131) );
NOR3_X1 U853 ( .A1(n1107), .A2(n1115), .A3(n1116), .ZN(n1033) );
NAND3_X1 U854 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1116) );
NAND3_X1 U855 ( .A1(n1189), .A2(n1190), .A3(n1027), .ZN(n1188) );
AND2_X1 U856 ( .A1(n1080), .A2(n1191), .ZN(n1027) );
NAND2_X1 U857 ( .A1(n1026), .A2(n1192), .ZN(n1190) );
INV_X1 U858 ( .A(KEYINPUT15), .ZN(n1192) );
NAND2_X1 U859 ( .A1(n1058), .A2(KEYINPUT15), .ZN(n1189) );
NOR2_X1 U860 ( .A1(n1145), .A2(n1026), .ZN(n1058) );
NAND3_X1 U861 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1115) );
OR2_X1 U862 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND4_X1 U863 ( .A1(n1198), .A2(n1145), .A3(n1199), .A4(n1048), .ZN(n1194) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1193) );
NAND3_X1 U865 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1201) );
NAND4_X1 U866 ( .A1(n1052), .A2(n1196), .A3(n1205), .A4(n1206), .ZN(n1204) );
INV_X1 U867 ( .A(KEYINPUT25), .ZN(n1196) );
INV_X1 U868 ( .A(n1080), .ZN(n1052) );
NAND4_X1 U869 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1107) );
AND4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1209) );
NOR2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND4_X1 U873 ( .A1(n1059), .A2(n1048), .A3(n1219), .A4(n1220), .ZN(n1208) );
INV_X1 U874 ( .A(n1221), .ZN(n1220) );
AND3_X1 U875 ( .A1(n1026), .A2(n1218), .A3(n1222), .ZN(n1219) );
INV_X1 U876 ( .A(KEYINPUT36), .ZN(n1218) );
NAND4_X1 U877 ( .A1(n1049), .A2(n1055), .A3(n1145), .A4(n1221), .ZN(n1207) );
NAND2_X1 U878 ( .A1(n1223), .A2(n1224), .ZN(n1055) );
NAND2_X1 U879 ( .A1(n1059), .A2(n1222), .ZN(n1224) );
NAND2_X1 U880 ( .A1(n1225), .A2(n1200), .ZN(n1223) );
XOR2_X1 U881 ( .A(n1226), .B(n1227), .Z(n1181) );
NAND2_X1 U882 ( .A1(KEYINPUT9), .A2(n1228), .ZN(n1226) );
NOR2_X1 U883 ( .A1(n1093), .A2(G952), .ZN(n1127) );
XOR2_X1 U884 ( .A(G146), .B(n1215), .Z(G48) );
AND3_X1 U885 ( .A1(n1229), .A2(n1200), .A3(n1145), .ZN(n1215) );
XNOR2_X1 U886 ( .A(G143), .B(n1214), .ZN(G45) );
NAND4_X1 U887 ( .A1(n1230), .A2(n1231), .A3(n1200), .A4(n1205), .ZN(n1214) );
XNOR2_X1 U888 ( .A(G140), .B(n1232), .ZN(G42) );
NAND3_X1 U889 ( .A1(n1145), .A2(n1059), .A3(n1233), .ZN(n1232) );
NOR3_X1 U890 ( .A1(n1234), .A2(KEYINPUT16), .A3(n1081), .ZN(n1233) );
INV_X1 U891 ( .A(n1049), .ZN(n1081) );
XNOR2_X1 U892 ( .A(G137), .B(n1213), .ZN(G39) );
NAND3_X1 U893 ( .A1(n1229), .A2(n1235), .A3(n1059), .ZN(n1213) );
XNOR2_X1 U894 ( .A(G134), .B(n1217), .ZN(G36) );
NAND3_X1 U895 ( .A1(n1231), .A2(n1026), .A3(n1059), .ZN(n1217) );
XNOR2_X1 U896 ( .A(G131), .B(n1212), .ZN(G33) );
NAND3_X1 U897 ( .A1(n1059), .A2(n1231), .A3(n1145), .ZN(n1212) );
AND2_X1 U898 ( .A1(n1236), .A2(n1048), .ZN(n1231) );
NOR2_X1 U899 ( .A1(n1050), .A2(n1066), .ZN(n1059) );
INV_X1 U900 ( .A(n1051), .ZN(n1066) );
XNOR2_X1 U901 ( .A(n1211), .B(n1237), .ZN(G30) );
NOR2_X1 U902 ( .A1(KEYINPUT45), .A2(n1238), .ZN(n1237) );
NAND3_X1 U903 ( .A1(n1026), .A2(n1200), .A3(n1229), .ZN(n1211) );
AND3_X1 U904 ( .A1(n1239), .A2(n1085), .A3(n1236), .ZN(n1229) );
INV_X1 U905 ( .A(n1234), .ZN(n1236) );
NAND2_X1 U906 ( .A1(n1222), .A2(n1221), .ZN(n1234) );
XNOR2_X1 U907 ( .A(n1240), .B(n1186), .ZN(G3) );
NAND3_X1 U908 ( .A1(n1235), .A2(n1191), .A3(n1048), .ZN(n1186) );
XNOR2_X1 U909 ( .A(G101), .B(KEYINPUT62), .ZN(n1240) );
XNOR2_X1 U910 ( .A(G125), .B(n1241), .ZN(G27) );
NAND4_X1 U911 ( .A1(n1200), .A2(n1221), .A3(n1049), .A4(n1242), .ZN(n1241) );
NOR2_X1 U912 ( .A1(n1043), .A2(n1243), .ZN(n1242) );
XOR2_X1 U913 ( .A(KEYINPUT37), .B(n1145), .Z(n1243) );
NAND2_X1 U914 ( .A1(n1035), .A2(n1244), .ZN(n1221) );
NAND3_X1 U915 ( .A1(G902), .A2(n1245), .A3(n1095), .ZN(n1244) );
AND2_X1 U916 ( .A1(n1246), .A2(G953), .ZN(n1095) );
XNOR2_X1 U917 ( .A(G900), .B(KEYINPUT22), .ZN(n1246) );
XNOR2_X1 U918 ( .A(G122), .B(n1197), .ZN(G24) );
NAND4_X1 U919 ( .A1(n1200), .A2(n1205), .A3(n1080), .A4(n1206), .ZN(n1197) );
NOR2_X1 U920 ( .A1(n1247), .A2(n1248), .ZN(n1206) );
NOR2_X1 U921 ( .A1(n1085), .A2(n1239), .ZN(n1080) );
XNOR2_X1 U922 ( .A(n1249), .B(n1250), .ZN(G21) );
NOR2_X1 U923 ( .A1(n1251), .A2(n1203), .ZN(n1250) );
NAND4_X1 U924 ( .A1(n1198), .A2(n1235), .A3(n1239), .A4(n1085), .ZN(n1203) );
XNOR2_X1 U925 ( .A(n1200), .B(KEYINPUT60), .ZN(n1251) );
XOR2_X1 U926 ( .A(n1252), .B(n1253), .Z(G18) );
NAND2_X1 U927 ( .A1(KEYINPUT23), .A2(G116), .ZN(n1253) );
NAND2_X1 U928 ( .A1(n1200), .A2(n1254), .ZN(n1252) );
XNOR2_X1 U929 ( .A(KEYINPUT26), .B(n1202), .ZN(n1254) );
NAND3_X1 U930 ( .A1(n1048), .A2(n1026), .A3(n1198), .ZN(n1202) );
NOR2_X1 U931 ( .A1(n1230), .A2(n1061), .ZN(n1026) );
INV_X1 U932 ( .A(n1248), .ZN(n1230) );
XNOR2_X1 U933 ( .A(G113), .B(n1255), .ZN(G15) );
NAND4_X1 U934 ( .A1(n1256), .A2(n1145), .A3(n1199), .A4(n1048), .ZN(n1255) );
AND2_X1 U935 ( .A1(n1257), .A2(n1085), .ZN(n1048) );
NOR2_X1 U936 ( .A1(n1248), .A2(n1205), .ZN(n1145) );
NOR2_X1 U937 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
NOR2_X1 U938 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U939 ( .A(KEYINPUT5), .ZN(n1261) );
AND2_X1 U940 ( .A1(n1043), .A2(n1262), .ZN(n1260) );
NOR2_X1 U941 ( .A1(KEYINPUT5), .A2(n1198), .ZN(n1258) );
INV_X1 U942 ( .A(n1247), .ZN(n1198) );
NAND2_X1 U943 ( .A1(n1225), .A2(n1262), .ZN(n1247) );
INV_X1 U944 ( .A(n1043), .ZN(n1225) );
NAND2_X1 U945 ( .A1(n1263), .A2(n1264), .ZN(n1043) );
XNOR2_X1 U946 ( .A(n1064), .B(KEYINPUT1), .ZN(n1263) );
XNOR2_X1 U947 ( .A(G110), .B(n1187), .ZN(G12) );
NAND3_X1 U948 ( .A1(n1235), .A2(n1191), .A3(n1049), .ZN(n1187) );
NOR2_X1 U949 ( .A1(n1085), .A2(n1257), .ZN(n1049) );
INV_X1 U950 ( .A(n1239), .ZN(n1257) );
XNOR2_X1 U951 ( .A(n1265), .B(n1086), .ZN(n1239) );
AND2_X1 U952 ( .A1(G217), .A2(n1266), .ZN(n1086) );
NAND2_X1 U953 ( .A1(n1130), .A2(n1185), .ZN(n1265) );
XOR2_X1 U954 ( .A(n1267), .B(n1268), .Z(n1130) );
XOR2_X1 U955 ( .A(n1122), .B(n1269), .Z(n1268) );
XOR2_X1 U956 ( .A(n1097), .B(n1270), .Z(n1269) );
NOR2_X1 U957 ( .A1(KEYINPUT48), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U958 ( .A(G125), .B(G140), .ZN(n1097) );
XNOR2_X1 U959 ( .A(G119), .B(G110), .ZN(n1122) );
XOR2_X1 U960 ( .A(n1272), .B(n1273), .Z(n1267) );
XNOR2_X1 U961 ( .A(G137), .B(n1238), .ZN(n1273) );
NAND2_X1 U962 ( .A1(G221), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U963 ( .A(n1275), .B(G472), .ZN(n1085) );
NAND2_X1 U964 ( .A1(n1276), .A2(n1185), .ZN(n1275) );
XOR2_X1 U965 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U966 ( .A(n1161), .B(n1279), .ZN(n1278) );
NOR2_X1 U967 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR2_X1 U968 ( .A1(KEYINPUT42), .A2(n1162), .ZN(n1281) );
AND2_X1 U969 ( .A1(KEYINPUT14), .A2(n1162), .ZN(n1280) );
XOR2_X1 U970 ( .A(n1282), .B(n1283), .Z(n1277) );
XNOR2_X1 U971 ( .A(G101), .B(n1150), .ZN(n1283) );
NAND3_X1 U972 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1150) );
OR2_X1 U973 ( .A1(G113), .A2(KEYINPUT55), .ZN(n1286) );
NAND3_X1 U974 ( .A1(KEYINPUT55), .A2(G113), .A3(n1287), .ZN(n1285) );
INV_X1 U975 ( .A(n1288), .ZN(n1287) );
NAND2_X1 U976 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
NAND2_X1 U977 ( .A1(KEYINPUT55), .A2(n1290), .ZN(n1289) );
XOR2_X1 U978 ( .A(KEYINPUT3), .B(G113), .Z(n1290) );
XOR2_X1 U979 ( .A(G116), .B(n1249), .Z(n1288) );
INV_X1 U980 ( .A(G119), .ZN(n1249) );
NAND2_X1 U981 ( .A1(KEYINPUT47), .A2(n1155), .ZN(n1282) );
AND3_X1 U982 ( .A1(n1291), .A2(n1093), .A3(G210), .ZN(n1155) );
AND3_X1 U983 ( .A1(n1199), .A2(n1262), .A3(n1222), .ZN(n1191) );
NOR2_X1 U984 ( .A1(n1264), .A2(n1064), .ZN(n1222) );
INV_X1 U985 ( .A(n1057), .ZN(n1064) );
NAND2_X1 U986 ( .A1(G221), .A2(n1266), .ZN(n1057) );
NAND2_X1 U987 ( .A1(G234), .A2(n1185), .ZN(n1266) );
INV_X1 U988 ( .A(n1056), .ZN(n1264) );
NAND3_X1 U989 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1056) );
NAND2_X1 U990 ( .A1(G469), .A2(n1068), .ZN(n1294) );
NAND2_X1 U991 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
INV_X1 U992 ( .A(KEYINPUT32), .ZN(n1296) );
NAND2_X1 U993 ( .A1(n1297), .A2(n1070), .ZN(n1295) );
INV_X1 U994 ( .A(G469), .ZN(n1070) );
XNOR2_X1 U995 ( .A(n1068), .B(n1298), .ZN(n1297) );
NAND2_X1 U996 ( .A1(KEYINPUT32), .A2(n1299), .ZN(n1292) );
NAND2_X1 U997 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U998 ( .A1(n1068), .A2(n1298), .ZN(n1301) );
OR3_X1 U999 ( .A1(n1068), .A2(G469), .A3(n1298), .ZN(n1300) );
INV_X1 U1000 ( .A(KEYINPUT18), .ZN(n1298) );
NAND2_X1 U1001 ( .A1(n1302), .A2(n1185), .ZN(n1068) );
XOR2_X1 U1002 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1003 ( .A(n1178), .B(n1305), .Z(n1304) );
XNOR2_X1 U1004 ( .A(KEYINPUT20), .B(n1177), .ZN(n1305) );
INV_X1 U1005 ( .A(G110), .ZN(n1177) );
AND2_X1 U1006 ( .A1(G227), .A2(n1093), .ZN(n1178) );
XNOR2_X1 U1007 ( .A(n1168), .B(n1179), .ZN(n1303) );
XOR2_X1 U1008 ( .A(G140), .B(KEYINPUT21), .Z(n1179) );
XNOR2_X1 U1009 ( .A(n1306), .B(n1307), .ZN(n1168) );
XNOR2_X1 U1010 ( .A(n1308), .B(n1309), .ZN(n1307) );
XNOR2_X1 U1011 ( .A(n1106), .B(n1103), .ZN(n1306) );
XNOR2_X1 U1012 ( .A(G128), .B(n1310), .ZN(n1103) );
INV_X1 U1013 ( .A(n1161), .ZN(n1106) );
XOR2_X1 U1014 ( .A(G131), .B(n1311), .Z(n1161) );
XOR2_X1 U1015 ( .A(G137), .B(G134), .Z(n1311) );
NAND2_X1 U1016 ( .A1(n1035), .A2(n1312), .ZN(n1262) );
NAND3_X1 U1017 ( .A1(n1117), .A2(n1245), .A3(G902), .ZN(n1312) );
AND2_X1 U1018 ( .A1(n1313), .A2(G953), .ZN(n1117) );
XNOR2_X1 U1019 ( .A(G898), .B(KEYINPUT56), .ZN(n1313) );
NAND3_X1 U1020 ( .A1(n1245), .A2(n1093), .A3(G952), .ZN(n1035) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1245) );
XNOR2_X1 U1022 ( .A(n1200), .B(KEYINPUT54), .ZN(n1199) );
AND2_X1 U1023 ( .A1(n1314), .A2(n1050), .ZN(n1200) );
OR2_X1 U1024 ( .A1(n1065), .A2(n1315), .ZN(n1050) );
AND2_X1 U1025 ( .A1(n1076), .A2(n1075), .ZN(n1315) );
NOR2_X1 U1026 ( .A1(n1075), .A2(n1076), .ZN(n1065) );
AND2_X1 U1027 ( .A1(n1316), .A2(n1185), .ZN(n1076) );
XNOR2_X1 U1028 ( .A(n1162), .B(n1317), .ZN(n1316) );
XNOR2_X1 U1029 ( .A(n1227), .B(n1228), .ZN(n1317) );
AND2_X1 U1030 ( .A1(G224), .A2(n1093), .ZN(n1228) );
XNOR2_X1 U1031 ( .A(n1318), .B(n1319), .ZN(n1227) );
XNOR2_X1 U1032 ( .A(n1320), .B(G110), .ZN(n1319) );
XOR2_X1 U1033 ( .A(n1321), .B(n1124), .Z(n1318) );
XNOR2_X1 U1034 ( .A(n1322), .B(KEYINPUT0), .ZN(n1124) );
NAND2_X1 U1035 ( .A1(KEYINPUT35), .A2(n1323), .ZN(n1321) );
XNOR2_X1 U1036 ( .A(n1324), .B(n1125), .ZN(n1323) );
XOR2_X1 U1037 ( .A(n1308), .B(n1325), .Z(n1125) );
NOR2_X1 U1038 ( .A1(KEYINPUT12), .A2(n1309), .ZN(n1325) );
XOR2_X1 U1039 ( .A(G104), .B(n1326), .Z(n1309) );
XNOR2_X1 U1040 ( .A(KEYINPUT27), .B(n1327), .ZN(n1326) );
INV_X1 U1041 ( .A(G101), .ZN(n1308) );
NOR2_X1 U1042 ( .A1(KEYINPUT24), .A2(n1328), .ZN(n1324) );
XNOR2_X1 U1043 ( .A(G119), .B(n1121), .ZN(n1328) );
XOR2_X1 U1044 ( .A(G113), .B(n1329), .Z(n1121) );
NOR2_X1 U1045 ( .A1(G116), .A2(KEYINPUT34), .ZN(n1329) );
XOR2_X1 U1046 ( .A(n1310), .B(n1330), .Z(n1162) );
XNOR2_X1 U1047 ( .A(n1331), .B(KEYINPUT57), .ZN(n1330) );
NAND2_X1 U1048 ( .A1(KEYINPUT38), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1049 ( .A(KEYINPUT46), .B(n1238), .ZN(n1332) );
XNOR2_X1 U1050 ( .A(G146), .B(n1333), .ZN(n1310) );
INV_X1 U1051 ( .A(G143), .ZN(n1333) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1334), .ZN(n1075) );
XNOR2_X1 U1053 ( .A(KEYINPUT58), .B(n1051), .ZN(n1314) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1334), .ZN(n1051) );
NAND2_X1 U1055 ( .A1(n1335), .A2(n1185), .ZN(n1334) );
XNOR2_X1 U1056 ( .A(G237), .B(KEYINPUT29), .ZN(n1335) );
INV_X1 U1057 ( .A(n1039), .ZN(n1235) );
NAND2_X1 U1058 ( .A1(n1336), .A2(n1248), .ZN(n1039) );
XOR2_X1 U1059 ( .A(n1337), .B(n1140), .Z(n1248) );
INV_X1 U1060 ( .A(G475), .ZN(n1140) );
NAND2_X1 U1061 ( .A1(KEYINPUT49), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1062 ( .A(KEYINPUT17), .B(n1339), .ZN(n1338) );
INV_X1 U1063 ( .A(n1087), .ZN(n1339) );
NOR2_X1 U1064 ( .A1(n1143), .A2(G902), .ZN(n1087) );
INV_X1 U1065 ( .A(n1139), .ZN(n1143) );
XNOR2_X1 U1066 ( .A(n1340), .B(n1341), .ZN(n1139) );
XOR2_X1 U1067 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1068 ( .A(G104), .B(n1344), .Z(n1343) );
NOR2_X1 U1069 ( .A1(KEYINPUT51), .A2(n1345), .ZN(n1344) );
XNOR2_X1 U1070 ( .A(G122), .B(G113), .ZN(n1345) );
XNOR2_X1 U1071 ( .A(G131), .B(n1320), .ZN(n1342) );
INV_X1 U1072 ( .A(G125), .ZN(n1320) );
XNOR2_X1 U1073 ( .A(n1271), .B(n1346), .ZN(n1340) );
XNOR2_X1 U1074 ( .A(n1347), .B(n1348), .ZN(n1346) );
NOR2_X1 U1075 ( .A1(G140), .A2(KEYINPUT7), .ZN(n1348) );
NAND2_X1 U1076 ( .A1(n1349), .A2(KEYINPUT59), .ZN(n1347) );
XNOR2_X1 U1077 ( .A(G143), .B(n1350), .ZN(n1349) );
AND3_X1 U1078 ( .A1(G214), .A2(n1093), .A3(n1291), .ZN(n1350) );
INV_X1 U1079 ( .A(G237), .ZN(n1291) );
XOR2_X1 U1080 ( .A(G146), .B(KEYINPUT53), .Z(n1271) );
XNOR2_X1 U1081 ( .A(KEYINPUT8), .B(n1061), .ZN(n1336) );
INV_X1 U1082 ( .A(n1205), .ZN(n1061) );
XNOR2_X1 U1083 ( .A(n1351), .B(G478), .ZN(n1205) );
NAND2_X1 U1084 ( .A1(n1135), .A2(n1185), .ZN(n1351) );
INV_X1 U1085 ( .A(G902), .ZN(n1185) );
XNOR2_X1 U1086 ( .A(n1352), .B(n1353), .ZN(n1135) );
XOR2_X1 U1087 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1088 ( .A(n1356), .B(n1357), .ZN(n1355) );
NAND2_X1 U1089 ( .A1(KEYINPUT63), .A2(n1327), .ZN(n1357) );
INV_X1 U1090 ( .A(G107), .ZN(n1327) );
NAND2_X1 U1091 ( .A1(KEYINPUT11), .A2(n1322), .ZN(n1356) );
INV_X1 U1092 ( .A(G122), .ZN(n1322) );
NAND2_X1 U1093 ( .A1(G217), .A2(n1274), .ZN(n1354) );
AND2_X1 U1094 ( .A1(G234), .A2(n1093), .ZN(n1274) );
INV_X1 U1095 ( .A(G953), .ZN(n1093) );
XOR2_X1 U1096 ( .A(n1358), .B(n1359), .Z(n1352) );
XNOR2_X1 U1097 ( .A(n1238), .B(G116), .ZN(n1359) );
INV_X1 U1098 ( .A(G128), .ZN(n1238) );
XNOR2_X1 U1099 ( .A(G134), .B(G143), .ZN(n1358) );
endmodule


