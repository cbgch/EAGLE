//Key = 0011111111101001000101010110110010010101101001011001101010101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329;

XOR2_X1 U734 ( .A(G107), .B(n1016), .Z(G9) );
NOR2_X1 U735 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U736 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NOR2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
XOR2_X1 U738 ( .A(n1025), .B(KEYINPUT43), .Z(n1023) );
NAND3_X1 U739 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1019) );
OR3_X1 U740 ( .A1(n1029), .A2(n1025), .A3(n1030), .ZN(n1028) );
NAND4_X1 U741 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1025) );
NAND3_X1 U742 ( .A1(n1035), .A2(n1036), .A3(n1031), .ZN(n1026) );
INV_X1 U743 ( .A(n1037), .ZN(n1031) );
NAND2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND3_X1 U745 ( .A1(n1034), .A2(n1040), .A3(n1032), .ZN(n1039) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U747 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U748 ( .A1(n1033), .A2(n1045), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U750 ( .A1(n1032), .A2(n1048), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U753 ( .A1(n1034), .A2(n1053), .ZN(n1046) );
NAND2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U755 ( .A(n1056), .B(KEYINPUT27), .Z(n1054) );
NOR3_X1 U756 ( .A1(n1022), .A2(G952), .A3(n1057), .ZN(n1017) );
INV_X1 U757 ( .A(n1027), .ZN(n1057) );
NAND4_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1027) );
NOR4_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NOR2_X1 U760 ( .A1(KEYINPUT61), .A2(G475), .ZN(n1063) );
AND2_X1 U761 ( .A1(n1066), .A2(KEYINPUT61), .ZN(n1062) );
XNOR2_X1 U762 ( .A(n1067), .B(n1068), .ZN(n1058) );
NOR2_X1 U763 ( .A1(G478), .A2(KEYINPUT38), .ZN(n1068) );
XOR2_X1 U764 ( .A(n1069), .B(n1070), .Z(G72) );
XOR2_X1 U765 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U766 ( .A1(G953), .A2(n1073), .ZN(n1072) );
NAND2_X1 U767 ( .A1(G900), .A2(G227), .ZN(n1073) );
NAND2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
NAND2_X1 U769 ( .A1(G953), .A2(n1076), .ZN(n1075) );
XOR2_X1 U770 ( .A(n1077), .B(n1078), .Z(n1074) );
XOR2_X1 U771 ( .A(n1079), .B(n1080), .Z(n1078) );
XOR2_X1 U772 ( .A(n1081), .B(n1082), .Z(n1077) );
NAND2_X1 U773 ( .A1(KEYINPUT28), .A2(n1083), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1084), .A2(G953), .ZN(n1069) );
XOR2_X1 U775 ( .A(n1085), .B(n1086), .Z(G69) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(n1086) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U778 ( .A1(G898), .A2(n1091), .ZN(n1089) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1091), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U781 ( .A(KEYINPUT40), .B(n1095), .ZN(n1094) );
NAND2_X1 U782 ( .A1(G953), .A2(n1096), .ZN(n1085) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1097), .A2(n1098), .ZN(G66) );
XNOR2_X1 U785 ( .A(n1099), .B(n1100), .ZN(n1098) );
NOR3_X1 U786 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
INV_X1 U787 ( .A(G217), .ZN(n1103) );
XOR2_X1 U788 ( .A(n1104), .B(KEYINPUT15), .Z(n1102) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1105), .ZN(G63) );
XOR2_X1 U790 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U791 ( .A1(KEYINPUT1), .A2(n1108), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U793 ( .A(n1111), .ZN(n1110) );
NOR2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1114), .A2(G478), .ZN(n1106) );
NOR2_X1 U796 ( .A1(n1097), .A2(n1115), .ZN(G60) );
XOR2_X1 U797 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U798 ( .A1(KEYINPUT17), .A2(n1118), .ZN(n1117) );
NAND2_X1 U799 ( .A1(n1114), .A2(G475), .ZN(n1116) );
XNOR2_X1 U800 ( .A(G104), .B(n1119), .ZN(G6) );
NOR2_X1 U801 ( .A1(n1097), .A2(n1120), .ZN(G57) );
XOR2_X1 U802 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1122) );
AND2_X1 U804 ( .A1(G472), .A2(n1114), .ZN(n1123) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1121) );
NOR2_X1 U806 ( .A1(KEYINPUT30), .A2(n1127), .ZN(n1126) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1125) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
XOR2_X1 U810 ( .A(n1134), .B(KEYINPUT7), .Z(n1132) );
NOR2_X1 U811 ( .A1(n1097), .A2(n1135), .ZN(G54) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U813 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U814 ( .A(n1140), .B(G110), .Z(n1139) );
XNOR2_X1 U815 ( .A(KEYINPUT5), .B(KEYINPUT13), .ZN(n1138) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1136) );
XNOR2_X1 U817 ( .A(n1143), .B(n1080), .ZN(n1142) );
XOR2_X1 U818 ( .A(G140), .B(n1144), .Z(n1080) );
NAND2_X1 U819 ( .A1(n1145), .A2(KEYINPUT37), .ZN(n1143) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U821 ( .A(n1148), .B(n1149), .ZN(n1141) );
NOR3_X1 U822 ( .A1(n1101), .A2(KEYINPUT57), .A3(n1150), .ZN(n1149) );
INV_X1 U823 ( .A(G469), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1097), .A2(n1151), .ZN(G51) );
NOR2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U826 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
XNOR2_X1 U828 ( .A(KEYINPUT11), .B(n1155), .ZN(n1157) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1155) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U831 ( .A1(KEYINPUT60), .A2(n1081), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1090), .B(n1079), .Z(n1158) );
XNOR2_X1 U833 ( .A(n1154), .B(KEYINPUT33), .ZN(n1156) );
AND2_X1 U834 ( .A1(n1114), .A2(n1162), .ZN(n1154) );
INV_X1 U835 ( .A(n1101), .ZN(n1114) );
NAND2_X1 U836 ( .A1(G902), .A2(n1020), .ZN(n1101) );
NAND3_X1 U837 ( .A1(n1093), .A2(n1095), .A3(n1084), .ZN(n1020) );
AND4_X1 U838 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1084) );
NOR4_X1 U839 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
NOR3_X1 U841 ( .A1(n1173), .A2(n1056), .A3(n1174), .ZN(n1172) );
XOR2_X1 U842 ( .A(KEYINPUT56), .B(n1035), .Z(n1173) );
AND4_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1119), .A4(n1177), .ZN(n1093) );
NOR4_X1 U844 ( .A1(n1016), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1177) );
AND3_X1 U845 ( .A1(n1034), .A2(n1181), .A3(n1182), .ZN(n1016) );
NAND3_X1 U846 ( .A1(n1034), .A2(n1181), .A3(n1183), .ZN(n1119) );
NOR2_X1 U847 ( .A1(n1091), .A2(G952), .ZN(n1097) );
XOR2_X1 U848 ( .A(G146), .B(n1171), .Z(G48) );
AND3_X1 U849 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1171) );
XOR2_X1 U850 ( .A(n1187), .B(n1163), .Z(G45) );
NAND4_X1 U851 ( .A1(n1188), .A2(n1184), .A3(n1189), .A4(n1066), .ZN(n1163) );
XNOR2_X1 U852 ( .A(G140), .B(n1164), .ZN(G42) );
NAND3_X1 U853 ( .A1(n1051), .A2(n1035), .A3(n1186), .ZN(n1164) );
NOR4_X1 U854 ( .A1(n1055), .A2(n1041), .A3(n1190), .A4(n1191), .ZN(n1186) );
XOR2_X1 U855 ( .A(G137), .B(n1168), .Z(G39) );
AND4_X1 U856 ( .A1(n1032), .A2(n1192), .A3(n1035), .A4(n1193), .ZN(n1168) );
INV_X1 U857 ( .A(n1041), .ZN(n1193) );
XOR2_X1 U858 ( .A(G134), .B(n1194), .Z(G36) );
NOR3_X1 U859 ( .A1(n1174), .A2(n1056), .A3(n1065), .ZN(n1194) );
XOR2_X1 U860 ( .A(G131), .B(n1170), .Z(G33) );
NOR3_X1 U861 ( .A1(n1055), .A2(n1065), .A3(n1174), .ZN(n1170) );
INV_X1 U862 ( .A(n1188), .ZN(n1174) );
NOR3_X1 U863 ( .A1(n1041), .A2(n1191), .A3(n1049), .ZN(n1188) );
INV_X1 U864 ( .A(n1035), .ZN(n1065) );
NOR2_X1 U865 ( .A1(n1029), .A2(n1195), .ZN(n1035) );
INV_X1 U866 ( .A(n1030), .ZN(n1195) );
INV_X1 U867 ( .A(n1183), .ZN(n1055) );
XOR2_X1 U868 ( .A(n1196), .B(n1197), .Z(G30) );
NOR2_X1 U869 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
AND2_X1 U870 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1199) );
AND4_X1 U871 ( .A1(n1192), .A2(n1182), .A3(n1200), .A4(n1184), .ZN(n1169) );
NOR2_X1 U872 ( .A1(KEYINPUT29), .A2(n1201), .ZN(n1198) );
NAND4_X1 U873 ( .A1(n1192), .A2(n1182), .A3(n1200), .A4(n1024), .ZN(n1201) );
NOR3_X1 U874 ( .A1(n1190), .A2(n1191), .A3(n1051), .ZN(n1192) );
XNOR2_X1 U875 ( .A(G101), .B(n1175), .ZN(G3) );
NAND3_X1 U876 ( .A1(n1032), .A2(n1181), .A3(n1202), .ZN(n1175) );
XOR2_X1 U877 ( .A(n1203), .B(n1204), .Z(G27) );
XOR2_X1 U878 ( .A(KEYINPUT58), .B(G125), .Z(n1204) );
NOR2_X1 U879 ( .A1(n1167), .A2(KEYINPUT59), .ZN(n1203) );
AND4_X1 U880 ( .A1(n1033), .A2(n1184), .A3(n1183), .A4(n1205), .ZN(n1167) );
NOR3_X1 U881 ( .A1(n1185), .A2(n1191), .A3(n1190), .ZN(n1205) );
AND2_X1 U882 ( .A1(n1037), .A2(n1206), .ZN(n1191) );
NAND4_X1 U883 ( .A1(G953), .A2(G902), .A3(n1207), .A4(n1076), .ZN(n1206) );
INV_X1 U884 ( .A(G900), .ZN(n1076) );
XNOR2_X1 U885 ( .A(G122), .B(n1176), .ZN(G24) );
NAND4_X1 U886 ( .A1(n1208), .A2(n1034), .A3(n1189), .A4(n1066), .ZN(n1176) );
INV_X1 U887 ( .A(n1064), .ZN(n1034) );
NAND2_X1 U888 ( .A1(n1190), .A2(n1051), .ZN(n1064) );
XOR2_X1 U889 ( .A(n1180), .B(n1209), .Z(G21) );
NOR2_X1 U890 ( .A1(KEYINPUT36), .A2(n1210), .ZN(n1209) );
AND4_X1 U891 ( .A1(n1208), .A2(n1032), .A3(n1185), .A4(n1052), .ZN(n1180) );
XNOR2_X1 U892 ( .A(G116), .B(n1095), .ZN(G18) );
NAND3_X1 U893 ( .A1(n1202), .A2(n1182), .A3(n1208), .ZN(n1095) );
INV_X1 U894 ( .A(n1056), .ZN(n1182) );
NAND2_X1 U895 ( .A1(n1211), .A2(n1189), .ZN(n1056) );
XOR2_X1 U896 ( .A(G113), .B(n1179), .Z(G15) );
AND3_X1 U897 ( .A1(n1202), .A2(n1183), .A3(n1208), .ZN(n1179) );
AND2_X1 U898 ( .A1(n1033), .A2(n1212), .ZN(n1208) );
NOR2_X1 U899 ( .A1(n1213), .A2(n1043), .ZN(n1033) );
INV_X1 U900 ( .A(n1059), .ZN(n1043) );
NOR2_X1 U901 ( .A1(n1189), .A2(n1211), .ZN(n1183) );
INV_X1 U902 ( .A(n1049), .ZN(n1202) );
NAND2_X1 U903 ( .A1(n1190), .A2(n1185), .ZN(n1049) );
INV_X1 U904 ( .A(n1051), .ZN(n1185) );
XOR2_X1 U905 ( .A(n1214), .B(n1215), .Z(G12) );
NAND2_X1 U906 ( .A1(KEYINPUT21), .A2(n1178), .ZN(n1215) );
AND4_X1 U907 ( .A1(n1032), .A2(n1181), .A3(n1051), .A4(n1052), .ZN(n1178) );
INV_X1 U908 ( .A(n1190), .ZN(n1052) );
XOR2_X1 U909 ( .A(n1216), .B(n1217), .Z(n1190) );
AND2_X1 U910 ( .A1(n1104), .A2(G217), .ZN(n1217) );
NAND2_X1 U911 ( .A1(n1218), .A2(n1099), .ZN(n1216) );
NAND2_X1 U912 ( .A1(n1219), .A2(n1220), .ZN(n1099) );
NAND2_X1 U913 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XNOR2_X1 U914 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U915 ( .A(n1225), .B(KEYINPUT48), .Z(n1221) );
NAND2_X1 U916 ( .A1(n1226), .A2(n1227), .ZN(n1219) );
XOR2_X1 U917 ( .A(n1223), .B(n1224), .Z(n1227) );
NAND2_X1 U918 ( .A1(KEYINPUT42), .A2(n1228), .ZN(n1224) );
INV_X1 U919 ( .A(G137), .ZN(n1228) );
NAND3_X1 U920 ( .A1(G234), .A2(n1091), .A3(G221), .ZN(n1223) );
XOR2_X1 U921 ( .A(n1225), .B(KEYINPUT16), .Z(n1226) );
XOR2_X1 U922 ( .A(n1229), .B(n1230), .Z(n1225) );
XNOR2_X1 U923 ( .A(n1231), .B(n1232), .ZN(n1230) );
NAND2_X1 U924 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
OR2_X1 U925 ( .A1(n1081), .A2(G140), .ZN(n1234) );
XOR2_X1 U926 ( .A(n1235), .B(KEYINPUT18), .Z(n1233) );
NAND2_X1 U927 ( .A1(G140), .A2(n1081), .ZN(n1235) );
XOR2_X1 U928 ( .A(n1214), .B(n1236), .Z(n1229) );
NOR2_X1 U929 ( .A1(KEYINPUT55), .A2(n1210), .ZN(n1236) );
XOR2_X1 U930 ( .A(n1237), .B(G472), .Z(n1051) );
NAND2_X1 U931 ( .A1(n1238), .A2(n1218), .ZN(n1237) );
XOR2_X1 U932 ( .A(n1127), .B(n1239), .Z(n1238) );
XOR2_X1 U933 ( .A(n1240), .B(G101), .Z(n1239) );
NAND2_X1 U934 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U935 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U936 ( .A(KEYINPUT6), .B(n1245), .Z(n1241) );
NOR2_X1 U937 ( .A1(n1243), .A2(n1244), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1246), .A2(n1131), .ZN(n1244) );
NAND2_X1 U939 ( .A1(n1134), .A2(n1247), .ZN(n1131) );
NAND2_X1 U940 ( .A1(n1248), .A2(n1133), .ZN(n1246) );
INV_X1 U941 ( .A(n1247), .ZN(n1133) );
XOR2_X1 U942 ( .A(n1134), .B(KEYINPUT63), .Z(n1248) );
XNOR2_X1 U943 ( .A(n1249), .B(n1129), .ZN(n1243) );
NOR2_X1 U944 ( .A1(KEYINPUT41), .A2(n1250), .ZN(n1129) );
XOR2_X1 U945 ( .A(n1210), .B(n1251), .Z(n1250) );
XOR2_X1 U946 ( .A(n1252), .B(KEYINPUT62), .Z(n1249) );
NAND3_X1 U947 ( .A1(n1253), .A2(n1091), .A3(G210), .ZN(n1127) );
AND2_X1 U948 ( .A1(n1212), .A2(n1200), .ZN(n1181) );
XOR2_X1 U949 ( .A(n1041), .B(KEYINPUT8), .Z(n1200) );
NAND2_X1 U950 ( .A1(n1213), .A2(n1059), .ZN(n1041) );
NAND2_X1 U951 ( .A1(G221), .A2(n1104), .ZN(n1059) );
NAND2_X1 U952 ( .A1(n1254), .A2(G234), .ZN(n1104) );
XOR2_X1 U953 ( .A(n1218), .B(KEYINPUT53), .Z(n1254) );
INV_X1 U954 ( .A(n1044), .ZN(n1213) );
XOR2_X1 U955 ( .A(n1060), .B(KEYINPUT31), .Z(n1044) );
XOR2_X1 U956 ( .A(n1255), .B(G469), .Z(n1060) );
NAND2_X1 U957 ( .A1(n1256), .A2(n1218), .ZN(n1255) );
XOR2_X1 U958 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U959 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U960 ( .A(n1214), .B(n1261), .Z(n1260) );
NOR2_X1 U961 ( .A1(G140), .A2(KEYINPUT50), .ZN(n1261) );
NAND2_X1 U962 ( .A1(KEYINPUT51), .A2(n1146), .ZN(n1259) );
XOR2_X1 U963 ( .A(n1134), .B(KEYINPUT47), .Z(n1146) );
XOR2_X1 U964 ( .A(n1262), .B(n1147), .Z(n1257) );
XNOR2_X1 U965 ( .A(n1263), .B(G101), .ZN(n1147) );
NAND2_X1 U966 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U967 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U968 ( .A(KEYINPUT10), .B(n1268), .Z(n1264) );
NOR2_X1 U969 ( .A1(n1266), .A2(n1267), .ZN(n1268) );
INV_X1 U970 ( .A(G107), .ZN(n1267) );
XNOR2_X1 U971 ( .A(n1269), .B(n1270), .ZN(n1262) );
NAND2_X1 U972 ( .A1(KEYINPUT25), .A2(n1247), .ZN(n1270) );
XOR2_X1 U973 ( .A(n1140), .B(n1144), .Z(n1247) );
XOR2_X1 U974 ( .A(G134), .B(G137), .Z(n1144) );
NAND2_X1 U975 ( .A1(KEYINPUT4), .A2(G131), .ZN(n1140) );
NAND2_X1 U976 ( .A1(KEYINPUT3), .A2(n1148), .ZN(n1269) );
AND2_X1 U977 ( .A1(G227), .A2(n1091), .ZN(n1148) );
AND2_X1 U978 ( .A1(n1184), .A2(n1271), .ZN(n1212) );
NAND2_X1 U979 ( .A1(n1272), .A2(n1037), .ZN(n1271) );
NAND3_X1 U980 ( .A1(n1273), .A2(n1207), .A3(G952), .ZN(n1037) );
INV_X1 U981 ( .A(n1022), .ZN(n1273) );
XOR2_X1 U982 ( .A(n1091), .B(KEYINPUT26), .Z(n1022) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1207), .A4(n1274), .ZN(n1272) );
INV_X1 U984 ( .A(G898), .ZN(n1274) );
NAND2_X1 U985 ( .A1(G234), .A2(G237), .ZN(n1207) );
INV_X1 U986 ( .A(n1024), .ZN(n1184) );
NAND2_X1 U987 ( .A1(n1029), .A2(n1030), .ZN(n1024) );
NAND2_X1 U988 ( .A1(G214), .A2(n1275), .ZN(n1030) );
XNOR2_X1 U989 ( .A(n1276), .B(n1162), .ZN(n1029) );
AND2_X1 U990 ( .A1(G210), .A2(n1275), .ZN(n1162) );
NAND2_X1 U991 ( .A1(n1253), .A2(n1218), .ZN(n1275) );
INV_X1 U992 ( .A(G237), .ZN(n1253) );
NAND2_X1 U993 ( .A1(n1277), .A2(n1218), .ZN(n1276) );
XOR2_X1 U994 ( .A(n1278), .B(n1279), .Z(n1277) );
INV_X1 U995 ( .A(n1090), .ZN(n1279) );
XOR2_X1 U996 ( .A(n1280), .B(n1281), .Z(n1090) );
XNOR2_X1 U997 ( .A(n1124), .B(n1282), .ZN(n1281) );
XOR2_X1 U998 ( .A(n1283), .B(n1251), .Z(n1282) );
NAND2_X1 U999 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
OR2_X1 U1000 ( .A1(n1214), .A2(G122), .ZN(n1285) );
XOR2_X1 U1001 ( .A(n1286), .B(KEYINPUT20), .Z(n1284) );
NAND2_X1 U1002 ( .A1(G122), .A2(n1214), .ZN(n1286) );
XOR2_X1 U1003 ( .A(G101), .B(G113), .Z(n1124) );
XOR2_X1 U1004 ( .A(n1287), .B(n1288), .Z(n1280) );
XOR2_X1 U1005 ( .A(G107), .B(n1289), .Z(n1288) );
NOR2_X1 U1006 ( .A1(KEYINPUT24), .A2(n1266), .ZN(n1289) );
NAND2_X1 U1007 ( .A1(KEYINPUT35), .A2(n1210), .ZN(n1287) );
INV_X1 U1008 ( .A(G119), .ZN(n1210) );
XNOR2_X1 U1009 ( .A(KEYINPUT45), .B(n1290), .ZN(n1278) );
NOR3_X1 U1010 ( .A1(KEYINPUT46), .A2(n1291), .A3(n1292), .ZN(n1290) );
NOR2_X1 U1011 ( .A1(n1081), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1012 ( .A(n1294), .B(KEYINPUT23), .Z(n1293) );
INV_X1 U1013 ( .A(G125), .ZN(n1081) );
NOR2_X1 U1014 ( .A1(G125), .A2(n1295), .ZN(n1291) );
XOR2_X1 U1015 ( .A(KEYINPUT39), .B(n1296), .Z(n1295) );
INV_X1 U1016 ( .A(n1294), .ZN(n1296) );
XOR2_X1 U1017 ( .A(n1160), .B(n1079), .Z(n1294) );
INV_X1 U1018 ( .A(n1134), .ZN(n1079) );
XOR2_X1 U1019 ( .A(n1187), .B(n1232), .Z(n1134) );
XNOR2_X1 U1020 ( .A(n1196), .B(G146), .ZN(n1232) );
INV_X1 U1021 ( .A(G128), .ZN(n1196) );
NAND2_X1 U1022 ( .A1(G224), .A2(n1091), .ZN(n1160) );
NOR2_X1 U1023 ( .A1(n1066), .A2(n1189), .ZN(n1032) );
XOR2_X1 U1024 ( .A(n1067), .B(n1297), .Z(n1189) );
XOR2_X1 U1025 ( .A(KEYINPUT32), .B(G478), .Z(n1297) );
NAND2_X1 U1026 ( .A1(n1218), .A2(n1298), .ZN(n1067) );
NAND2_X1 U1027 ( .A1(n1299), .A2(n1111), .ZN(n1298) );
NAND2_X1 U1028 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
OR2_X1 U1029 ( .A1(n1113), .A2(n1112), .ZN(n1299) );
XOR2_X1 U1030 ( .A(n1300), .B(n1301), .Z(n1112) );
XOR2_X1 U1031 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1032 ( .A(G128), .B(G122), .Z(n1303) );
XOR2_X1 U1033 ( .A(KEYINPUT34), .B(G143), .Z(n1302) );
XOR2_X1 U1034 ( .A(n1304), .B(n1251), .Z(n1300) );
XOR2_X1 U1035 ( .A(G116), .B(KEYINPUT14), .Z(n1251) );
XOR2_X1 U1036 ( .A(n1305), .B(G107), .Z(n1304) );
NAND2_X1 U1037 ( .A1(KEYINPUT12), .A2(n1306), .ZN(n1305) );
INV_X1 U1038 ( .A(G134), .ZN(n1306) );
NAND3_X1 U1039 ( .A1(G217), .A2(n1091), .A3(G234), .ZN(n1113) );
INV_X1 U1040 ( .A(G902), .ZN(n1218) );
INV_X1 U1041 ( .A(n1211), .ZN(n1066) );
XOR2_X1 U1042 ( .A(n1307), .B(G475), .Z(n1211) );
OR2_X1 U1043 ( .A1(n1118), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1044 ( .A(n1308), .B(n1309), .ZN(n1118) );
XOR2_X1 U1045 ( .A(n1310), .B(n1311), .Z(n1309) );
NAND2_X1 U1046 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1047 ( .A1(KEYINPUT0), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1048 ( .A1(KEYINPUT9), .A2(n1315), .ZN(n1312) );
INV_X1 U1049 ( .A(n1314), .ZN(n1315) );
XOR2_X1 U1050 ( .A(n1316), .B(G146), .Z(n1314) );
NAND2_X1 U1051 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
OR2_X1 U1052 ( .A1(n1319), .A2(G125), .ZN(n1318) );
XOR2_X1 U1053 ( .A(n1320), .B(KEYINPUT44), .Z(n1317) );
NAND2_X1 U1054 ( .A1(G125), .A2(n1319), .ZN(n1320) );
XOR2_X1 U1055 ( .A(G140), .B(KEYINPUT19), .Z(n1319) );
NAND2_X1 U1056 ( .A1(n1321), .A2(n1322), .ZN(n1310) );
NAND2_X1 U1057 ( .A1(n1323), .A2(n1083), .ZN(n1322) );
INV_X1 U1058 ( .A(G131), .ZN(n1083) );
XOR2_X1 U1059 ( .A(n1324), .B(KEYINPUT22), .Z(n1323) );
NAND2_X1 U1060 ( .A1(n1325), .A2(G131), .ZN(n1321) );
XOR2_X1 U1061 ( .A(n1324), .B(KEYINPUT54), .Z(n1325) );
XOR2_X1 U1062 ( .A(n1326), .B(n1327), .Z(n1324) );
NOR2_X1 U1063 ( .A1(KEYINPUT49), .A2(n1187), .ZN(n1327) );
INV_X1 U1064 ( .A(G143), .ZN(n1187) );
NAND3_X1 U1065 ( .A1(n1328), .A2(n1091), .A3(G214), .ZN(n1326) );
INV_X1 U1066 ( .A(G953), .ZN(n1091) );
XOR2_X1 U1067 ( .A(KEYINPUT52), .B(G237), .Z(n1328) );
XNOR2_X1 U1068 ( .A(n1329), .B(n1266), .ZN(n1308) );
XNOR2_X1 U1069 ( .A(G104), .B(KEYINPUT2), .ZN(n1266) );
XOR2_X1 U1070 ( .A(n1252), .B(G122), .Z(n1329) );
INV_X1 U1071 ( .A(G113), .ZN(n1252) );
INV_X1 U1072 ( .A(G110), .ZN(n1214) );
endmodule


