//Key = 0110011100101001001000100101110010100101100011111110111010011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;

XNOR2_X1 U731 ( .A(G107), .B(n1002), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
NAND2_X1 U734 ( .A1(G952), .A2(n1009), .ZN(n1006) );
NAND2_X1 U735 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U736 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U737 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U738 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND3_X1 U739 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1018) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1021) );
NAND2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U745 ( .A1(n1023), .A2(n1031), .A3(n1027), .ZN(n1016) );
XOR2_X1 U746 ( .A(KEYINPUT40), .B(n1032), .Z(n1012) );
NOR3_X1 U747 ( .A1(n1019), .A2(n1033), .A3(n1034), .ZN(n1032) );
XNOR2_X1 U748 ( .A(n1027), .B(KEYINPUT30), .ZN(n1033) );
NAND4_X1 U749 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1005) );
NAND3_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1036) );
XNOR2_X1 U751 ( .A(KEYINPUT59), .B(n1042), .ZN(n1041) );
NAND2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1035) );
XNOR2_X1 U753 ( .A(n1039), .B(KEYINPUT53), .ZN(n1043) );
NOR3_X1 U754 ( .A1(n1045), .A2(n1046), .A3(n1034), .ZN(n1039) );
NAND3_X1 U755 ( .A1(n1020), .A2(n1023), .A3(n1014), .ZN(n1034) );
INV_X1 U756 ( .A(n1047), .ZN(n1014) );
NOR3_X1 U757 ( .A1(n1048), .A2(G953), .A3(n1049), .ZN(n1003) );
INV_X1 U758 ( .A(n1037), .ZN(n1049) );
NAND4_X1 U759 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1037) );
NOR4_X1 U760 ( .A1(n1054), .A2(n1040), .A3(n1046), .A4(n1055), .ZN(n1053) );
NAND3_X1 U761 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1054) );
NAND2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR3_X1 U763 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1052) );
AND2_X1 U764 ( .A1(G469), .A2(KEYINPUT31), .ZN(n1063) );
NOR2_X1 U765 ( .A1(KEYINPUT31), .A2(n1064), .ZN(n1062) );
XNOR2_X1 U766 ( .A(n1065), .B(n1066), .ZN(n1061) );
XOR2_X1 U767 ( .A(n1067), .B(KEYINPUT23), .Z(n1051) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1050) );
XNOR2_X1 U769 ( .A(KEYINPUT20), .B(n1070), .ZN(n1048) );
XOR2_X1 U770 ( .A(n1071), .B(n1072), .Z(G72) );
XOR2_X1 U771 ( .A(n1073), .B(n1074), .Z(n1072) );
NAND2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
INV_X1 U773 ( .A(n1077), .ZN(n1076) );
XOR2_X1 U774 ( .A(n1078), .B(n1079), .Z(n1075) );
XNOR2_X1 U775 ( .A(n1080), .B(n1081), .ZN(n1079) );
XOR2_X1 U776 ( .A(n1082), .B(n1083), .Z(n1078) );
XNOR2_X1 U777 ( .A(n1084), .B(n1085), .ZN(n1082) );
NAND2_X1 U778 ( .A1(KEYINPUT47), .A2(G125), .ZN(n1085) );
NAND3_X1 U779 ( .A1(n1086), .A2(n1087), .A3(KEYINPUT44), .ZN(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT52), .A2(n1088), .ZN(n1087) );
OR3_X1 U781 ( .A1(n1089), .A2(G134), .A3(KEYINPUT52), .ZN(n1086) );
INV_X1 U782 ( .A(G137), .ZN(n1089) );
NAND2_X1 U783 ( .A1(n1090), .A2(n1007), .ZN(n1073) );
XNOR2_X1 U784 ( .A(G953), .B(KEYINPUT4), .ZN(n1090) );
NOR2_X1 U785 ( .A1(n1091), .A2(n1038), .ZN(n1071) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1091) );
XOR2_X1 U787 ( .A(n1092), .B(n1093), .Z(G69) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U789 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U790 ( .A(KEYINPUT21), .B(n1098), .Z(n1097) );
NOR2_X1 U791 ( .A1(G898), .A2(n1038), .ZN(n1098) );
XOR2_X1 U792 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U793 ( .A(n1101), .B(KEYINPUT8), .ZN(n1100) );
NAND2_X1 U794 ( .A1(KEYINPUT49), .A2(n1102), .ZN(n1101) );
NAND3_X1 U795 ( .A1(n1008), .A2(n1038), .A3(KEYINPUT54), .ZN(n1094) );
NAND2_X1 U796 ( .A1(G953), .A2(n1103), .ZN(n1092) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1103) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U800 ( .A1(n1108), .A2(n1059), .ZN(n1106) );
NOR3_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G63) );
AND2_X1 U802 ( .A1(KEYINPUT1), .A2(n1104), .ZN(n1111) );
NOR3_X1 U803 ( .A1(KEYINPUT1), .A2(G953), .A3(G952), .ZN(n1110) );
NOR3_X1 U804 ( .A1(n1066), .A2(n1112), .A3(n1113), .ZN(n1109) );
AND3_X1 U805 ( .A1(n1114), .A2(G478), .A3(n1108), .ZN(n1113) );
NOR2_X1 U806 ( .A1(n1115), .A2(n1114), .ZN(n1112) );
NOR2_X1 U807 ( .A1(n1116), .A2(n1065), .ZN(n1115) );
NOR2_X1 U808 ( .A1(n1007), .A2(n1008), .ZN(n1116) );
NOR2_X1 U809 ( .A1(n1104), .A2(n1117), .ZN(G60) );
XOR2_X1 U810 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U811 ( .A1(n1108), .A2(G475), .ZN(n1118) );
XNOR2_X1 U812 ( .A(G104), .B(n1120), .ZN(G6) );
NOR2_X1 U813 ( .A1(n1104), .A2(n1121), .ZN(G57) );
XOR2_X1 U814 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U815 ( .A(n1124), .B(n1125), .ZN(n1123) );
NOR2_X1 U816 ( .A1(KEYINPUT0), .A2(n1126), .ZN(n1122) );
XOR2_X1 U817 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U818 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U819 ( .A1(KEYINPUT51), .A2(n1131), .ZN(n1130) );
XOR2_X1 U820 ( .A(G116), .B(n1132), .Z(n1131) );
NAND2_X1 U821 ( .A1(KEYINPUT28), .A2(n1133), .ZN(n1129) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(n1127) );
NAND2_X1 U823 ( .A1(n1108), .A2(G472), .ZN(n1134) );
NOR3_X1 U824 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(G54) );
AND2_X1 U825 ( .A1(n1104), .A2(KEYINPUT50), .ZN(n1138) );
NOR3_X1 U826 ( .A1(KEYINPUT50), .A2(n1038), .A3(n1070), .ZN(n1137) );
INV_X1 U827 ( .A(G952), .ZN(n1070) );
XOR2_X1 U828 ( .A(n1139), .B(n1140), .Z(n1136) );
XOR2_X1 U829 ( .A(n1080), .B(n1141), .Z(n1140) );
XOR2_X1 U830 ( .A(n1142), .B(n1133), .Z(n1141) );
NAND2_X1 U831 ( .A1(KEYINPUT37), .A2(n1143), .ZN(n1142) );
XOR2_X1 U832 ( .A(n1144), .B(n1145), .Z(n1139) );
XOR2_X1 U833 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U834 ( .A1(n1108), .A2(G469), .ZN(n1147) );
NAND2_X1 U835 ( .A1(KEYINPUT5), .A2(n1148), .ZN(n1144) );
NOR2_X1 U836 ( .A1(n1104), .A2(n1149), .ZN(G51) );
XOR2_X1 U837 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U838 ( .A(n1152), .B(n1153), .Z(n1150) );
NOR2_X1 U839 ( .A1(KEYINPUT57), .A2(n1154), .ZN(n1153) );
NAND2_X1 U840 ( .A1(n1108), .A2(n1155), .ZN(n1152) );
AND2_X1 U841 ( .A1(G902), .A2(n1156), .ZN(n1108) );
OR2_X1 U842 ( .A1(n1008), .A2(n1007), .ZN(n1156) );
NAND4_X1 U843 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1007) );
AND4_X1 U844 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NOR3_X1 U845 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1159) );
NOR2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
INV_X1 U847 ( .A(KEYINPUT7), .ZN(n1169) );
NOR4_X1 U848 ( .A1(KEYINPUT7), .A2(n1170), .A3(n1045), .A4(n1171), .ZN(n1166) );
NAND3_X1 U849 ( .A1(n1172), .A2(n1173), .A3(n1068), .ZN(n1170) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1175), .ZN(n1165) );
XNOR2_X1 U851 ( .A(n1176), .B(KEYINPUT41), .ZN(n1174) );
NAND4_X1 U852 ( .A1(n1120), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1008) );
AND4_X1 U853 ( .A1(n1002), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1179) );
NAND3_X1 U854 ( .A1(n1183), .A2(n1023), .A3(n1184), .ZN(n1002) );
NOR3_X1 U855 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1178) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U857 ( .A(n1190), .B(KEYINPUT63), .Z(n1189) );
NAND2_X1 U858 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR4_X1 U859 ( .A1(n1044), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1186) );
INV_X1 U860 ( .A(n1023), .ZN(n1194) );
NAND3_X1 U861 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
NOR2_X1 U862 ( .A1(n1199), .A2(n1197), .ZN(n1185) );
INV_X1 U863 ( .A(KEYINPUT46), .ZN(n1197) );
NAND3_X1 U864 ( .A1(n1184), .A2(n1023), .A3(n1191), .ZN(n1120) );
NOR2_X1 U865 ( .A1(n1038), .A2(G952), .ZN(n1104) );
XNOR2_X1 U866 ( .A(G146), .B(n1157), .ZN(G48) );
NAND3_X1 U867 ( .A1(n1191), .A2(n1200), .A3(n1201), .ZN(n1157) );
XNOR2_X1 U868 ( .A(G143), .B(n1158), .ZN(G45) );
NAND3_X1 U869 ( .A1(n1202), .A2(n1176), .A3(n1201), .ZN(n1158) );
INV_X1 U870 ( .A(n1171), .ZN(n1201) );
XNOR2_X1 U871 ( .A(G140), .B(n1164), .ZN(G42) );
OR2_X1 U872 ( .A1(n1175), .A2(n1030), .ZN(n1164) );
NAND2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(G39) );
OR2_X1 U874 ( .A1(n1205), .A2(n1168), .ZN(n1204) );
XOR2_X1 U875 ( .A(n1206), .B(KEYINPUT9), .Z(n1203) );
NAND2_X1 U876 ( .A1(n1205), .A2(n1168), .ZN(n1206) );
NAND4_X1 U877 ( .A1(n1207), .A2(n1027), .A3(n1068), .A4(n1173), .ZN(n1168) );
XOR2_X1 U878 ( .A(G137), .B(KEYINPUT19), .Z(n1205) );
XNOR2_X1 U879 ( .A(G134), .B(n1163), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1176), .A2(n1183), .A3(n1207), .ZN(n1163) );
NAND2_X1 U881 ( .A1(n1208), .A2(n1209), .ZN(G33) );
NAND4_X1 U882 ( .A1(n1210), .A2(n1176), .A3(n1211), .A4(n1212), .ZN(n1209) );
NAND2_X1 U883 ( .A1(G131), .A2(n1213), .ZN(n1212) );
OR2_X1 U884 ( .A1(G131), .A2(KEYINPUT56), .ZN(n1211) );
NAND3_X1 U885 ( .A1(n1214), .A2(n1213), .A3(G131), .ZN(n1208) );
INV_X1 U886 ( .A(KEYINPUT36), .ZN(n1213) );
NAND3_X1 U887 ( .A1(n1210), .A2(n1176), .A3(KEYINPUT56), .ZN(n1214) );
INV_X1 U888 ( .A(n1175), .ZN(n1210) );
NAND2_X1 U889 ( .A1(n1207), .A2(n1191), .ZN(n1175) );
INV_X1 U890 ( .A(n1025), .ZN(n1191) );
NOR2_X1 U891 ( .A1(n1171), .A2(n1172), .ZN(n1207) );
INV_X1 U892 ( .A(n1010), .ZN(n1172) );
NAND2_X1 U893 ( .A1(n1215), .A2(n1216), .ZN(n1010) );
OR2_X1 U894 ( .A1(n1188), .A2(KEYINPUT59), .ZN(n1216) );
INV_X1 U895 ( .A(n1044), .ZN(n1188) );
NAND3_X1 U896 ( .A1(n1042), .A2(n1217), .A3(KEYINPUT59), .ZN(n1215) );
NAND2_X1 U897 ( .A1(n1031), .A2(n1218), .ZN(n1171) );
XOR2_X1 U898 ( .A(n1219), .B(KEYINPUT14), .Z(n1031) );
XNOR2_X1 U899 ( .A(G128), .B(n1162), .ZN(G30) );
NAND4_X1 U900 ( .A1(n1200), .A2(n1183), .A3(n1219), .A4(n1218), .ZN(n1162) );
XOR2_X1 U901 ( .A(n1177), .B(n1220), .Z(G3) );
XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n1124), .ZN(n1220) );
NAND3_X1 U903 ( .A1(n1027), .A2(n1184), .A3(n1176), .ZN(n1177) );
INV_X1 U904 ( .A(n1221), .ZN(n1184) );
XNOR2_X1 U905 ( .A(G125), .B(n1161), .ZN(G27) );
NAND4_X1 U906 ( .A1(n1218), .A2(n1019), .A3(n1044), .A4(n1222), .ZN(n1161) );
NOR3_X1 U907 ( .A1(n1025), .A2(n1030), .A3(n1223), .ZN(n1222) );
NAND2_X1 U908 ( .A1(n1047), .A2(n1224), .ZN(n1218) );
NAND3_X1 U909 ( .A1(G902), .A2(n1225), .A3(n1077), .ZN(n1224) );
NOR2_X1 U910 ( .A1(n1038), .A2(G900), .ZN(n1077) );
XNOR2_X1 U911 ( .A(n1199), .B(n1226), .ZN(G24) );
NOR2_X1 U912 ( .A1(KEYINPUT38), .A2(n1227), .ZN(n1226) );
NAND3_X1 U913 ( .A1(n1228), .A2(n1023), .A3(n1202), .ZN(n1199) );
AND3_X1 U914 ( .A1(n1198), .A2(n1196), .A3(n1044), .ZN(n1202) );
NOR2_X1 U915 ( .A1(n1173), .A2(n1068), .ZN(n1023) );
XNOR2_X1 U916 ( .A(G119), .B(n1182), .ZN(G21) );
NAND3_X1 U917 ( .A1(n1228), .A2(n1027), .A3(n1200), .ZN(n1182) );
AND3_X1 U918 ( .A1(n1068), .A2(n1173), .A3(n1044), .ZN(n1200) );
INV_X1 U919 ( .A(n1195), .ZN(n1228) );
XNOR2_X1 U920 ( .A(G116), .B(n1181), .ZN(G18) );
NAND3_X1 U921 ( .A1(n1183), .A2(n1044), .A3(n1192), .ZN(n1181) );
INV_X1 U922 ( .A(n1026), .ZN(n1183) );
NAND2_X1 U923 ( .A1(n1229), .A2(n1198), .ZN(n1026) );
XOR2_X1 U924 ( .A(n1196), .B(KEYINPUT25), .Z(n1229) );
XNOR2_X1 U925 ( .A(G113), .B(n1230), .ZN(G15) );
NAND3_X1 U926 ( .A1(n1192), .A2(n1231), .A3(n1232), .ZN(n1230) );
XNOR2_X1 U927 ( .A(n1044), .B(KEYINPUT34), .ZN(n1232) );
XNOR2_X1 U928 ( .A(KEYINPUT11), .B(n1025), .ZN(n1231) );
NAND2_X1 U929 ( .A1(n1233), .A2(n1196), .ZN(n1025) );
INV_X1 U930 ( .A(n1198), .ZN(n1233) );
NOR2_X1 U931 ( .A1(n1029), .A2(n1195), .ZN(n1192) );
NAND3_X1 U932 ( .A1(n1234), .A2(n1019), .A3(n1020), .ZN(n1195) );
INV_X1 U933 ( .A(n1176), .ZN(n1029) );
NOR2_X1 U934 ( .A1(n1173), .A2(n1235), .ZN(n1176) );
XNOR2_X1 U935 ( .A(G110), .B(n1180), .ZN(G12) );
OR3_X1 U936 ( .A1(n1030), .A2(n1221), .A3(n1045), .ZN(n1180) );
INV_X1 U937 ( .A(n1027), .ZN(n1045) );
NOR2_X1 U938 ( .A1(n1198), .A2(n1196), .ZN(n1027) );
NAND2_X1 U939 ( .A1(n1056), .A2(n1067), .ZN(n1196) );
NAND3_X1 U940 ( .A1(n1236), .A2(n1237), .A3(n1119), .ZN(n1067) );
INV_X1 U941 ( .A(G475), .ZN(n1236) );
NAND2_X1 U942 ( .A1(G475), .A2(n1238), .ZN(n1056) );
NAND2_X1 U943 ( .A1(n1119), .A2(n1237), .ZN(n1238) );
XOR2_X1 U944 ( .A(n1239), .B(n1240), .Z(n1119) );
XOR2_X1 U945 ( .A(n1241), .B(n1242), .Z(n1240) );
NAND2_X1 U946 ( .A1(KEYINPUT15), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U947 ( .A(n1083), .B(n1244), .ZN(n1243) );
XOR2_X1 U948 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U949 ( .A1(KEYINPUT58), .A2(n1247), .ZN(n1246) );
NAND3_X1 U950 ( .A1(n1248), .A2(n1038), .A3(G214), .ZN(n1245) );
NAND2_X1 U951 ( .A1(n1249), .A2(n1250), .ZN(n1241) );
NAND2_X1 U952 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U953 ( .A(n1253), .ZN(n1251) );
XOR2_X1 U954 ( .A(n1254), .B(KEYINPUT42), .Z(n1249) );
NAND2_X1 U955 ( .A1(G146), .A2(n1253), .ZN(n1254) );
XNOR2_X1 U956 ( .A(G104), .B(n1255), .ZN(n1239) );
XNOR2_X1 U957 ( .A(n1227), .B(G113), .ZN(n1255) );
NAND2_X1 U958 ( .A1(n1256), .A2(n1257), .ZN(n1198) );
NAND2_X1 U959 ( .A1(n1258), .A2(n1065), .ZN(n1257) );
XOR2_X1 U960 ( .A(KEYINPUT18), .B(n1259), .Z(n1256) );
NOR2_X1 U961 ( .A1(n1065), .A2(n1258), .ZN(n1259) );
XOR2_X1 U962 ( .A(KEYINPUT55), .B(n1066), .Z(n1258) );
NOR2_X1 U963 ( .A1(n1114), .A2(G902), .ZN(n1066) );
XOR2_X1 U964 ( .A(n1260), .B(n1261), .Z(n1114) );
NOR2_X1 U965 ( .A1(KEYINPUT33), .A2(n1262), .ZN(n1261) );
XOR2_X1 U966 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U967 ( .A(G116), .B(n1265), .Z(n1264) );
XNOR2_X1 U968 ( .A(G134), .B(n1227), .ZN(n1265) );
XNOR2_X1 U969 ( .A(n1266), .B(n1267), .ZN(n1263) );
XNOR2_X1 U970 ( .A(G107), .B(n1247), .ZN(n1266) );
NAND2_X1 U971 ( .A1(G217), .A2(n1268), .ZN(n1260) );
INV_X1 U972 ( .A(G478), .ZN(n1065) );
NAND3_X1 U973 ( .A1(n1219), .A2(n1234), .A3(n1044), .ZN(n1221) );
NOR2_X1 U974 ( .A1(n1042), .A2(n1040), .ZN(n1044) );
INV_X1 U975 ( .A(n1217), .ZN(n1040) );
NAND2_X1 U976 ( .A1(G214), .A2(n1269), .ZN(n1217) );
XOR2_X1 U977 ( .A(n1069), .B(KEYINPUT27), .Z(n1042) );
XNOR2_X1 U978 ( .A(n1270), .B(n1155), .ZN(n1069) );
AND2_X1 U979 ( .A1(G210), .A2(n1269), .ZN(n1155) );
NAND2_X1 U980 ( .A1(n1248), .A2(n1237), .ZN(n1269) );
NAND2_X1 U981 ( .A1(n1271), .A2(n1237), .ZN(n1270) );
XOR2_X1 U982 ( .A(n1154), .B(n1272), .Z(n1271) );
XNOR2_X1 U983 ( .A(n1151), .B(KEYINPUT43), .ZN(n1272) );
XNOR2_X1 U984 ( .A(n1273), .B(n1099), .ZN(n1151) );
XNOR2_X1 U985 ( .A(G110), .B(n1227), .ZN(n1099) );
INV_X1 U986 ( .A(G122), .ZN(n1227) );
XOR2_X1 U987 ( .A(n1274), .B(n1275), .Z(n1273) );
AND2_X1 U988 ( .A1(n1038), .A2(G224), .ZN(n1275) );
NAND2_X1 U989 ( .A1(KEYINPUT2), .A2(n1102), .ZN(n1274) );
XOR2_X1 U990 ( .A(n1276), .B(n1277), .Z(n1102) );
XNOR2_X1 U991 ( .A(n1278), .B(n1279), .ZN(n1276) );
NOR2_X1 U992 ( .A1(G116), .A2(KEYINPUT26), .ZN(n1279) );
XNOR2_X1 U993 ( .A(n1135), .B(G125), .ZN(n1154) );
NAND2_X1 U994 ( .A1(n1047), .A2(n1280), .ZN(n1234) );
NAND4_X1 U995 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1281), .ZN(n1280) );
INV_X1 U996 ( .A(G898), .ZN(n1281) );
NAND3_X1 U997 ( .A1(n1225), .A2(n1038), .A3(G952), .ZN(n1047) );
NAND2_X1 U998 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U999 ( .A1(n1020), .A2(n1046), .ZN(n1219) );
INV_X1 U1000 ( .A(n1019), .ZN(n1046) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1282), .ZN(n1019) );
INV_X1 U1002 ( .A(n1223), .ZN(n1020) );
NAND2_X1 U1003 ( .A1(n1283), .A2(n1064), .ZN(n1223) );
NAND3_X1 U1004 ( .A1(n1284), .A2(n1237), .A3(n1285), .ZN(n1064) );
INV_X1 U1005 ( .A(G469), .ZN(n1284) );
XOR2_X1 U1006 ( .A(n1057), .B(KEYINPUT17), .Z(n1283) );
NAND2_X1 U1007 ( .A1(G469), .A2(n1286), .ZN(n1057) );
NAND2_X1 U1008 ( .A1(n1285), .A2(n1237), .ZN(n1286) );
XNOR2_X1 U1009 ( .A(n1287), .B(n1288), .ZN(n1285) );
XOR2_X1 U1010 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1011 ( .A(n1291), .B(n1146), .ZN(n1290) );
NAND2_X1 U1012 ( .A1(n1292), .A2(G227), .ZN(n1146) );
XNOR2_X1 U1013 ( .A(G953), .B(KEYINPUT16), .ZN(n1292) );
NAND2_X1 U1014 ( .A1(KEYINPUT48), .A2(n1293), .ZN(n1291) );
XOR2_X1 U1015 ( .A(KEYINPUT60), .B(n1143), .Z(n1293) );
XNOR2_X1 U1016 ( .A(n1294), .B(n1277), .ZN(n1143) );
XNOR2_X1 U1017 ( .A(n1295), .B(G107), .ZN(n1277) );
INV_X1 U1018 ( .A(G104), .ZN(n1295) );
NAND2_X1 U1019 ( .A1(KEYINPUT45), .A2(n1124), .ZN(n1294) );
INV_X1 U1020 ( .A(G101), .ZN(n1124) );
NAND2_X1 U1021 ( .A1(KEYINPUT12), .A2(n1133), .ZN(n1289) );
XNOR2_X1 U1022 ( .A(n1080), .B(n1148), .ZN(n1287) );
XOR2_X1 U1023 ( .A(G110), .B(n1081), .Z(n1148) );
XNOR2_X1 U1024 ( .A(n1296), .B(n1297), .ZN(n1080) );
NAND2_X1 U1025 ( .A1(KEYINPUT32), .A2(n1247), .ZN(n1296) );
NAND2_X1 U1026 ( .A1(n1235), .A2(n1173), .ZN(n1030) );
NAND3_X1 U1027 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1173) );
INV_X1 U1028 ( .A(n1055), .ZN(n1300) );
NOR2_X1 U1029 ( .A1(n1060), .A2(n1059), .ZN(n1055) );
NAND2_X1 U1030 ( .A1(KEYINPUT24), .A2(n1301), .ZN(n1299) );
NAND3_X1 U1031 ( .A1(n1060), .A2(n1302), .A3(n1059), .ZN(n1298) );
INV_X1 U1032 ( .A(n1301), .ZN(n1059) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1282), .ZN(n1301) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1237), .ZN(n1282) );
INV_X1 U1035 ( .A(KEYINPUT24), .ZN(n1302) );
NAND2_X1 U1036 ( .A1(n1107), .A2(n1237), .ZN(n1060) );
XOR2_X1 U1037 ( .A(n1303), .B(n1304), .Z(n1107) );
XNOR2_X1 U1038 ( .A(n1305), .B(n1306), .ZN(n1304) );
XOR2_X1 U1039 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U1040 ( .A1(KEYINPUT35), .A2(G110), .ZN(n1308) );
NAND2_X1 U1041 ( .A1(n1268), .A2(G221), .ZN(n1307) );
AND2_X1 U1042 ( .A1(G234), .A2(n1038), .ZN(n1268) );
XOR2_X1 U1043 ( .A(n1309), .B(n1310), .Z(n1303) );
NOR2_X1 U1044 ( .A1(KEYINPUT61), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1045 ( .A(n1253), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1046 ( .A(KEYINPUT22), .B(n1252), .ZN(n1312) );
INV_X1 U1047 ( .A(G146), .ZN(n1252) );
XOR2_X1 U1048 ( .A(G125), .B(n1081), .Z(n1253) );
XOR2_X1 U1049 ( .A(G140), .B(KEYINPUT13), .Z(n1081) );
XNOR2_X1 U1050 ( .A(G119), .B(G137), .ZN(n1309) );
INV_X1 U1051 ( .A(n1068), .ZN(n1235) );
XNOR2_X1 U1052 ( .A(n1313), .B(G472), .ZN(n1068) );
NAND2_X1 U1053 ( .A1(n1314), .A2(n1237), .ZN(n1313) );
INV_X1 U1054 ( .A(G902), .ZN(n1237) );
XOR2_X1 U1055 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1056 ( .A(n1317), .B(n1318), .ZN(n1316) );
INV_X1 U1057 ( .A(n1278), .ZN(n1318) );
XOR2_X1 U1058 ( .A(G101), .B(n1132), .Z(n1278) );
XOR2_X1 U1059 ( .A(G113), .B(G119), .Z(n1132) );
XOR2_X1 U1060 ( .A(n1135), .B(n1133), .Z(n1317) );
XOR2_X1 U1061 ( .A(n1083), .B(n1088), .Z(n1133) );
XNOR2_X1 U1062 ( .A(G134), .B(G137), .ZN(n1088) );
XOR2_X1 U1063 ( .A(G131), .B(KEYINPUT29), .Z(n1083) );
XOR2_X1 U1064 ( .A(n1297), .B(n1319), .Z(n1135) );
XOR2_X1 U1065 ( .A(KEYINPUT3), .B(n1247), .Z(n1319) );
XOR2_X1 U1066 ( .A(G143), .B(KEYINPUT62), .Z(n1247) );
XNOR2_X1 U1067 ( .A(G146), .B(n1267), .ZN(n1297) );
INV_X1 U1068 ( .A(n1305), .ZN(n1267) );
XOR2_X1 U1069 ( .A(G128), .B(KEYINPUT6), .Z(n1305) );
XNOR2_X1 U1070 ( .A(n1125), .B(n1320), .ZN(n1315) );
XOR2_X1 U1071 ( .A(KEYINPUT10), .B(G116), .Z(n1320) );
AND3_X1 U1072 ( .A1(n1248), .A2(n1038), .A3(G210), .ZN(n1125) );
INV_X1 U1073 ( .A(G953), .ZN(n1038) );
INV_X1 U1074 ( .A(G237), .ZN(n1248) );
endmodule


