//Key = 0010100101100101010011011011001110010011011111000001100110000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;

XOR2_X1 U716 ( .A(n975), .B(n976), .Z(G9) );
NAND2_X1 U717 ( .A1(KEYINPUT20), .A2(G107), .ZN(n976) );
NOR2_X1 U718 ( .A1(n977), .A2(n978), .ZN(G75) );
NOR4_X1 U719 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n978) );
XOR2_X1 U720 ( .A(n983), .B(KEYINPUT57), .Z(n981) );
NAND2_X1 U721 ( .A1(n984), .A2(n985), .ZN(n983) );
NAND3_X1 U722 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n985) );
NAND3_X1 U723 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n987) );
NAND4_X1 U724 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .ZN(n991) );
NAND3_X1 U725 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n990) );
NAND3_X1 U726 ( .A1(n999), .A2(n1000), .A3(n992), .ZN(n989) );
NAND2_X1 U727 ( .A1(n1001), .A2(n1002), .ZN(n984) );
NAND4_X1 U728 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n979) );
NAND3_X1 U729 ( .A1(n986), .A2(n1007), .A3(n988), .ZN(n1004) );
NAND2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U731 ( .A1(n992), .A2(n1010), .ZN(n1009) );
NAND2_X1 U732 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U733 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
XNOR2_X1 U734 ( .A(n1000), .B(KEYINPUT52), .ZN(n1013) );
NAND2_X1 U735 ( .A1(n993), .A2(n1015), .ZN(n1011) );
NAND2_X1 U736 ( .A1(n996), .A2(n1016), .ZN(n1008) );
NAND2_X1 U737 ( .A1(n1001), .A2(n1017), .ZN(n1003) );
AND3_X1 U738 ( .A1(n996), .A2(n992), .A3(n988), .ZN(n1001) );
INV_X1 U739 ( .A(n1018), .ZN(n988) );
AND2_X1 U740 ( .A1(n1000), .A2(n993), .ZN(n996) );
NOR3_X1 U741 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n977) );
INV_X1 U742 ( .A(n1005), .ZN(n1019) );
NAND4_X1 U743 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1005) );
NOR4_X1 U744 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
XOR2_X1 U745 ( .A(G475), .B(n1028), .Z(n1027) );
XOR2_X1 U746 ( .A(KEYINPUT12), .B(n1029), .Z(n1026) );
XOR2_X1 U747 ( .A(n1030), .B(KEYINPUT24), .Z(n1024) );
NOR3_X1 U748 ( .A1(n1031), .A2(n994), .A3(n998), .ZN(n1022) );
XOR2_X1 U749 ( .A(n1032), .B(n1033), .Z(n1021) );
XNOR2_X1 U750 ( .A(G469), .B(KEYINPUT56), .ZN(n1033) );
XOR2_X1 U751 ( .A(KEYINPUT30), .B(n1034), .Z(n1020) );
XOR2_X1 U752 ( .A(n1035), .B(n1036), .Z(G72) );
NOR2_X1 U753 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR3_X1 U754 ( .A1(n980), .A2(KEYINPUT14), .A3(n1039), .ZN(n1038) );
NOR2_X1 U755 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NOR2_X1 U756 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U757 ( .A1(G953), .A2(n1044), .ZN(n1043) );
AND2_X1 U758 ( .A1(n1044), .A2(KEYINPUT14), .ZN(n1042) );
INV_X1 U759 ( .A(n1039), .ZN(n1044) );
NAND2_X1 U760 ( .A1(n1045), .A2(n1046), .ZN(n1039) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XOR2_X1 U762 ( .A(n1049), .B(n1050), .Z(n1045) );
XOR2_X1 U763 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U764 ( .A(G125), .B(n1053), .Z(n1049) );
INV_X1 U765 ( .A(n980), .ZN(n1040) );
NAND2_X1 U766 ( .A1(G953), .A2(n1054), .ZN(n1035) );
NAND2_X1 U767 ( .A1(G900), .A2(G227), .ZN(n1054) );
XOR2_X1 U768 ( .A(n1055), .B(n1056), .Z(G69) );
XOR2_X1 U769 ( .A(n1057), .B(n1058), .Z(n1056) );
NAND2_X1 U770 ( .A1(n1006), .A2(n1059), .ZN(n1058) );
NAND3_X1 U771 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR3_X1 U772 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
INV_X1 U773 ( .A(n975), .ZN(n1064) );
XNOR2_X1 U774 ( .A(KEYINPUT44), .B(n1066), .ZN(n1061) );
NAND2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(n1057) );
NAND2_X1 U776 ( .A1(n1047), .A2(n1069), .ZN(n1068) );
XOR2_X1 U777 ( .A(KEYINPUT13), .B(n1070), .Z(n1067) );
NOR2_X1 U778 ( .A1(n1071), .A2(n1006), .ZN(n1055) );
AND2_X1 U779 ( .A1(G224), .A2(G898), .ZN(n1071) );
NOR2_X1 U780 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XOR2_X1 U781 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U782 ( .A1(n1076), .A2(G217), .ZN(n1074) );
NOR2_X1 U783 ( .A1(n1072), .A2(n1077), .ZN(G63) );
XOR2_X1 U784 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U785 ( .A1(n1076), .A2(G478), .ZN(n1078) );
NOR2_X1 U786 ( .A1(n1072), .A2(n1080), .ZN(G60) );
NOR3_X1 U787 ( .A1(n1028), .A2(n1081), .A3(n1082), .ZN(n1080) );
AND3_X1 U788 ( .A1(n1083), .A2(G475), .A3(n1076), .ZN(n1082) );
NOR2_X1 U789 ( .A1(n1084), .A2(n1083), .ZN(n1081) );
NOR2_X1 U790 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U791 ( .A(G475), .ZN(n1086) );
XOR2_X1 U792 ( .A(n1087), .B(n1066), .Z(G6) );
NOR2_X1 U793 ( .A1(n1072), .A2(n1088), .ZN(G57) );
NOR2_X1 U794 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U795 ( .A(KEYINPUT54), .B(n1091), .Z(n1090) );
NOR2_X1 U796 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U797 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U798 ( .A1(n1096), .A2(n1097), .ZN(n1089) );
XOR2_X1 U799 ( .A(n1095), .B(n1094), .Z(n1097) );
NAND2_X1 U800 ( .A1(KEYINPUT32), .A2(n1098), .ZN(n1094) );
NAND3_X1 U801 ( .A1(n1099), .A2(n1100), .A3(G472), .ZN(n1098) );
OR2_X1 U802 ( .A1(n1076), .A2(KEYINPUT37), .ZN(n1100) );
NAND2_X1 U803 ( .A1(KEYINPUT37), .A2(n1101), .ZN(n1099) );
OR2_X1 U804 ( .A1(n1085), .A2(G902), .ZN(n1101) );
NAND2_X1 U805 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
NAND2_X1 U806 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U807 ( .A(n1106), .B(KEYINPUT18), .Z(n1104) );
XOR2_X1 U808 ( .A(n1107), .B(KEYINPUT50), .Z(n1102) );
OR2_X1 U809 ( .A1(n1105), .A2(n1106), .ZN(n1107) );
NOR2_X1 U810 ( .A1(n1072), .A2(n1108), .ZN(G54) );
XOR2_X1 U811 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U812 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U813 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U814 ( .A(n1115), .B(n1116), .Z(n1111) );
NOR2_X1 U815 ( .A1(KEYINPUT28), .A2(n1117), .ZN(n1116) );
NAND2_X1 U816 ( .A1(n1076), .A2(G469), .ZN(n1115) );
XOR2_X1 U817 ( .A(n1118), .B(n1119), .Z(n1109) );
XOR2_X1 U818 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U819 ( .A(n1122), .B(G131), .Z(n1118) );
NAND2_X1 U820 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND4_X1 U821 ( .A1(KEYINPUT42), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1124) );
NAND2_X1 U822 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
NAND2_X1 U823 ( .A1(n1126), .A2(n1130), .ZN(n1129) );
OR2_X1 U824 ( .A1(n1127), .A2(n1125), .ZN(n1130) );
INV_X1 U825 ( .A(KEYINPUT19), .ZN(n1127) );
NAND2_X1 U826 ( .A1(KEYINPUT42), .A2(n1125), .ZN(n1128) );
XNOR2_X1 U827 ( .A(n1131), .B(n1132), .ZN(n1125) );
XOR2_X1 U828 ( .A(n1133), .B(KEYINPUT34), .Z(n1131) );
NOR2_X1 U829 ( .A1(n1134), .A2(n1135), .ZN(G51) );
XOR2_X1 U830 ( .A(KEYINPUT47), .B(n1072), .Z(n1135) );
NOR2_X1 U831 ( .A1(n1006), .A2(G952), .ZN(n1072) );
XNOR2_X1 U832 ( .A(n1136), .B(n1137), .ZN(n1134) );
XOR2_X1 U833 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U834 ( .A1(n1076), .A2(n1140), .ZN(n1138) );
NOR2_X1 U835 ( .A1(n1141), .A2(n1085), .ZN(n1076) );
NOR2_X1 U836 ( .A1(n982), .A2(n1142), .ZN(n1085) );
XOR2_X1 U837 ( .A(KEYINPUT11), .B(n980), .Z(n1142) );
NAND4_X1 U838 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n980) );
AND4_X1 U839 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NAND2_X1 U840 ( .A1(n1002), .A2(n1151), .ZN(n1145) );
NAND2_X1 U841 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U842 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XNOR2_X1 U843 ( .A(KEYINPUT26), .B(n1156), .ZN(n1154) );
NAND2_X1 U844 ( .A1(n1014), .A2(n1157), .ZN(n1152) );
NAND2_X1 U845 ( .A1(n1158), .A2(n1060), .ZN(n982) );
AND4_X1 U846 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1060) );
NOR2_X1 U847 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U848 ( .A1(KEYINPUT36), .A2(n1165), .ZN(n1164) );
NOR3_X1 U849 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1163) );
INV_X1 U850 ( .A(KEYINPUT27), .ZN(n1166) );
NAND4_X1 U851 ( .A1(n992), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1161) );
NAND2_X1 U852 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
NAND3_X1 U853 ( .A1(n986), .A2(n1156), .A3(KEYINPUT36), .ZN(n1173) );
OR2_X1 U854 ( .A1(n1168), .A2(KEYINPUT27), .ZN(n1172) );
XOR2_X1 U855 ( .A(n1174), .B(KEYINPUT41), .Z(n1158) );
NAND4_X1 U856 ( .A1(n1175), .A2(n1066), .A3(n1176), .A4(n975), .ZN(n1174) );
NAND3_X1 U857 ( .A1(n1002), .A2(n993), .A3(n1177), .ZN(n975) );
NAND3_X1 U858 ( .A1(n1177), .A2(n993), .A3(n1017), .ZN(n1066) );
XOR2_X1 U859 ( .A(KEYINPUT9), .B(n1063), .Z(n1175) );
XNOR2_X1 U860 ( .A(G146), .B(n1150), .ZN(G48) );
NAND3_X1 U861 ( .A1(n1017), .A2(n1156), .A3(n1155), .ZN(n1150) );
XNOR2_X1 U862 ( .A(G143), .B(n1143), .ZN(G45) );
NAND4_X1 U863 ( .A1(n1155), .A2(n1014), .A3(n1178), .A4(n1179), .ZN(n1143) );
XNOR2_X1 U864 ( .A(G140), .B(n1149), .ZN(G42) );
NAND3_X1 U865 ( .A1(n1017), .A2(n1157), .A3(n999), .ZN(n1149) );
XNOR2_X1 U866 ( .A(G137), .B(n1148), .ZN(G39) );
NAND3_X1 U867 ( .A1(n1157), .A2(n1156), .A3(n986), .ZN(n1148) );
XOR2_X1 U868 ( .A(n1180), .B(n1181), .Z(G36) );
NOR3_X1 U869 ( .A1(n1168), .A2(KEYINPUT0), .A3(n1182), .ZN(n1181) );
NAND2_X1 U870 ( .A1(n1014), .A2(n1002), .ZN(n1168) );
XNOR2_X1 U871 ( .A(G134), .B(KEYINPUT15), .ZN(n1180) );
XOR2_X1 U872 ( .A(n1183), .B(n1147), .Z(G33) );
NAND3_X1 U873 ( .A1(n1017), .A2(n1157), .A3(n1014), .ZN(n1147) );
INV_X1 U874 ( .A(n1182), .ZN(n1157) );
NAND3_X1 U875 ( .A1(n1016), .A2(n1184), .A3(n1000), .ZN(n1182) );
AND2_X1 U876 ( .A1(n995), .A2(n1185), .ZN(n1000) );
XNOR2_X1 U877 ( .A(n1186), .B(KEYINPUT40), .ZN(n995) );
XOR2_X1 U878 ( .A(n1133), .B(n1187), .Z(G30) );
NAND4_X1 U879 ( .A1(KEYINPUT45), .A2(n1155), .A3(n1002), .A4(n1156), .ZN(n1187) );
AND2_X1 U880 ( .A1(n1188), .A2(n1016), .ZN(n1155) );
XNOR2_X1 U881 ( .A(G101), .B(n1189), .ZN(G3) );
NAND2_X1 U882 ( .A1(KEYINPUT43), .A2(n1063), .ZN(n1189) );
AND3_X1 U883 ( .A1(n1014), .A2(n1177), .A3(n986), .ZN(n1063) );
XOR2_X1 U884 ( .A(n1190), .B(n1144), .Z(G27) );
NAND4_X1 U885 ( .A1(n992), .A2(n1188), .A3(n999), .A4(n1017), .ZN(n1144) );
AND2_X1 U886 ( .A1(n1015), .A2(n1184), .ZN(n1188) );
NAND2_X1 U887 ( .A1(n1191), .A2(n1018), .ZN(n1184) );
NAND2_X1 U888 ( .A1(n1192), .A2(n1048), .ZN(n1191) );
INV_X1 U889 ( .A(G900), .ZN(n1048) );
XNOR2_X1 U890 ( .A(G122), .B(n1159), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1178), .A2(n1193), .A3(n993), .A4(n1179), .ZN(n1159) );
NOR2_X1 U892 ( .A1(n1194), .A2(n1025), .ZN(n993) );
XOR2_X1 U893 ( .A(n1195), .B(n1165), .Z(G21) );
NAND3_X1 U894 ( .A1(n986), .A2(n1156), .A3(n1193), .ZN(n1165) );
NAND2_X1 U895 ( .A1(n1196), .A2(n1197), .ZN(n1156) );
NAND2_X1 U896 ( .A1(n999), .A2(n1198), .ZN(n1197) );
INV_X1 U897 ( .A(KEYINPUT7), .ZN(n1198) );
NAND3_X1 U898 ( .A1(n1025), .A2(n1194), .A3(KEYINPUT7), .ZN(n1196) );
INV_X1 U899 ( .A(n1199), .ZN(n1194) );
XNOR2_X1 U900 ( .A(G116), .B(n1200), .ZN(G18) );
NAND4_X1 U901 ( .A1(n1201), .A2(KEYINPUT38), .A3(n1193), .A4(n1014), .ZN(n1200) );
XNOR2_X1 U902 ( .A(n1002), .B(KEYINPUT61), .ZN(n1201) );
NOR2_X1 U903 ( .A1(n1178), .A2(n1030), .ZN(n1002) );
XNOR2_X1 U904 ( .A(G113), .B(n1160), .ZN(G15) );
NAND3_X1 U905 ( .A1(n1014), .A2(n1017), .A3(n1193), .ZN(n1160) );
INV_X1 U906 ( .A(n1167), .ZN(n1193) );
NAND3_X1 U907 ( .A1(n1015), .A2(n1170), .A3(n992), .ZN(n1167) );
AND2_X1 U908 ( .A1(n997), .A2(n1202), .ZN(n992) );
AND2_X1 U909 ( .A1(n1178), .A2(n1030), .ZN(n1017) );
NOR2_X1 U910 ( .A1(n1025), .A2(n1199), .ZN(n1014) );
XOR2_X1 U911 ( .A(G110), .B(n1065), .Z(G12) );
INV_X1 U912 ( .A(n1176), .ZN(n1065) );
NAND3_X1 U913 ( .A1(n999), .A2(n1177), .A3(n986), .ZN(n1176) );
NOR2_X1 U914 ( .A1(n1179), .A2(n1178), .ZN(n986) );
XNOR2_X1 U915 ( .A(n1028), .B(n1203), .ZN(n1178) );
NOR2_X1 U916 ( .A1(G475), .A2(KEYINPUT1), .ZN(n1203) );
NOR2_X1 U917 ( .A1(n1083), .A2(G902), .ZN(n1028) );
XNOR2_X1 U918 ( .A(n1204), .B(n1205), .ZN(n1083) );
XOR2_X1 U919 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U920 ( .A(G125), .B(G122), .Z(n1207) );
XOR2_X1 U921 ( .A(KEYINPUT31), .B(G140), .Z(n1206) );
XOR2_X1 U922 ( .A(n1208), .B(n1209), .Z(n1204) );
XOR2_X1 U923 ( .A(G113), .B(G104), .Z(n1209) );
XOR2_X1 U924 ( .A(n1210), .B(n1211), .Z(n1208) );
AND2_X1 U925 ( .A1(G214), .A2(n1212), .ZN(n1211) );
INV_X1 U926 ( .A(n1030), .ZN(n1179) );
XOR2_X1 U927 ( .A(n1213), .B(G478), .Z(n1030) );
NAND2_X1 U928 ( .A1(n1079), .A2(n1141), .ZN(n1213) );
XNOR2_X1 U929 ( .A(n1214), .B(n1215), .ZN(n1079) );
XNOR2_X1 U930 ( .A(n1216), .B(n1217), .ZN(n1215) );
NOR2_X1 U931 ( .A1(G107), .A2(KEYINPUT53), .ZN(n1217) );
NAND2_X1 U932 ( .A1(n1218), .A2(KEYINPUT39), .ZN(n1216) );
XOR2_X1 U933 ( .A(n1133), .B(n1219), .Z(n1218) );
XOR2_X1 U934 ( .A(G143), .B(G134), .Z(n1219) );
INV_X1 U935 ( .A(G128), .ZN(n1133) );
XOR2_X1 U936 ( .A(n1220), .B(n1221), .Z(n1214) );
XOR2_X1 U937 ( .A(G122), .B(G116), .Z(n1221) );
NAND2_X1 U938 ( .A1(G217), .A2(n1222), .ZN(n1220) );
AND3_X1 U939 ( .A1(n1015), .A2(n1170), .A3(n1016), .ZN(n1177) );
NOR2_X1 U940 ( .A1(n997), .A2(n998), .ZN(n1016) );
INV_X1 U941 ( .A(n1202), .ZN(n998) );
NAND2_X1 U942 ( .A1(G221), .A2(n1223), .ZN(n1202) );
NAND2_X1 U943 ( .A1(G234), .A2(n1141), .ZN(n1223) );
XNOR2_X1 U944 ( .A(n1032), .B(n1224), .ZN(n997) );
NOR2_X1 U945 ( .A1(G469), .A2(KEYINPUT3), .ZN(n1224) );
NAND2_X1 U946 ( .A1(n1225), .A2(n1141), .ZN(n1032) );
XOR2_X1 U947 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U948 ( .A(n1228), .B(n1126), .ZN(n1227) );
XOR2_X1 U949 ( .A(G101), .B(n1229), .Z(n1126) );
NOR2_X1 U950 ( .A1(KEYINPUT49), .A2(n1230), .ZN(n1229) );
XOR2_X1 U951 ( .A(G107), .B(n1231), .Z(n1230) );
NOR2_X1 U952 ( .A1(KEYINPUT16), .A2(n1087), .ZN(n1231) );
INV_X1 U953 ( .A(G104), .ZN(n1087) );
XOR2_X1 U954 ( .A(G128), .B(n1232), .Z(n1226) );
NOR2_X1 U955 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U956 ( .A(KEYINPUT29), .B(n1235), .Z(n1234) );
AND2_X1 U957 ( .A1(n1236), .A2(n1121), .ZN(n1235) );
NOR2_X1 U958 ( .A1(n1236), .A2(n1237), .ZN(n1233) );
XOR2_X1 U959 ( .A(KEYINPUT46), .B(n1121), .Z(n1237) );
AND2_X1 U960 ( .A1(G227), .A2(n1006), .ZN(n1121) );
XNOR2_X1 U961 ( .A(n1238), .B(n1114), .ZN(n1236) );
XOR2_X1 U962 ( .A(G140), .B(KEYINPUT48), .Z(n1114) );
NAND2_X1 U963 ( .A1(KEYINPUT2), .A2(n1117), .ZN(n1238) );
NAND2_X1 U964 ( .A1(n1018), .A2(n1239), .ZN(n1170) );
NAND2_X1 U965 ( .A1(n1192), .A2(n1069), .ZN(n1239) );
INV_X1 U966 ( .A(G898), .ZN(n1069) );
AND3_X1 U967 ( .A1(n1047), .A2(n1240), .A3(G902), .ZN(n1192) );
XOR2_X1 U968 ( .A(G953), .B(KEYINPUT22), .Z(n1047) );
NAND3_X1 U969 ( .A1(n1240), .A2(n1006), .A3(G952), .ZN(n1018) );
NAND2_X1 U970 ( .A1(G237), .A2(G234), .ZN(n1240) );
INV_X1 U971 ( .A(n1171), .ZN(n1015) );
NAND2_X1 U972 ( .A1(n1186), .A2(n1185), .ZN(n1171) );
XOR2_X1 U973 ( .A(n994), .B(KEYINPUT35), .Z(n1185) );
AND2_X1 U974 ( .A1(n1241), .A2(n1242), .ZN(n994) );
XOR2_X1 U975 ( .A(KEYINPUT6), .B(G214), .Z(n1241) );
XOR2_X1 U976 ( .A(n1243), .B(n1029), .Z(n1186) );
XNOR2_X1 U977 ( .A(n1244), .B(n1140), .ZN(n1029) );
AND2_X1 U978 ( .A1(G210), .A2(n1242), .ZN(n1140) );
OR2_X1 U979 ( .A1(G902), .A2(G237), .ZN(n1242) );
NAND2_X1 U980 ( .A1(n1245), .A2(n1141), .ZN(n1244) );
XOR2_X1 U981 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U982 ( .A(KEYINPUT60), .B(KEYINPUT51), .Z(n1247) );
XOR2_X1 U983 ( .A(n1248), .B(n1249), .Z(n1246) );
INV_X1 U984 ( .A(n1139), .ZN(n1249) );
XOR2_X1 U985 ( .A(n1250), .B(n1070), .Z(n1139) );
XNOR2_X1 U986 ( .A(n1251), .B(n1252), .ZN(n1070) );
XOR2_X1 U987 ( .A(G122), .B(G110), .Z(n1252) );
XOR2_X1 U988 ( .A(n1106), .B(n1253), .Z(n1251) );
NOR2_X1 U989 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U990 ( .A(n1256), .B(KEYINPUT21), .Z(n1255) );
NAND2_X1 U991 ( .A1(G101), .A2(n1257), .ZN(n1256) );
NOR2_X1 U992 ( .A1(G101), .A2(n1257), .ZN(n1254) );
XOR2_X1 U993 ( .A(G107), .B(G104), .Z(n1257) );
NAND2_X1 U994 ( .A1(G224), .A2(n1006), .ZN(n1250) );
INV_X1 U995 ( .A(G953), .ZN(n1006) );
NAND2_X1 U996 ( .A1(KEYINPUT17), .A2(n1136), .ZN(n1248) );
XNOR2_X1 U997 ( .A(n1132), .B(n1258), .ZN(n1136) );
XOR2_X1 U998 ( .A(G125), .B(n1259), .Z(n1258) );
XNOR2_X1 U999 ( .A(KEYINPUT8), .B(KEYINPUT23), .ZN(n1243) );
AND2_X1 U1000 ( .A1(n1199), .A2(n1025), .ZN(n999) );
NAND3_X1 U1001 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1025) );
OR2_X1 U1002 ( .A1(n1263), .A2(n1075), .ZN(n1262) );
NAND3_X1 U1003 ( .A1(n1075), .A2(n1263), .A3(n1141), .ZN(n1261) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1264), .ZN(n1263) );
XOR2_X1 U1005 ( .A(n1265), .B(n1266), .Z(n1075) );
XOR2_X1 U1006 ( .A(n1053), .B(n1267), .Z(n1266) );
XNOR2_X1 U1007 ( .A(n1268), .B(n1269), .ZN(n1267) );
NOR2_X1 U1008 ( .A1(KEYINPUT25), .A2(n1190), .ZN(n1269) );
INV_X1 U1009 ( .A(G125), .ZN(n1190) );
NAND2_X1 U1010 ( .A1(KEYINPUT4), .A2(n1195), .ZN(n1268) );
INV_X1 U1011 ( .A(G119), .ZN(n1195) );
XOR2_X1 U1012 ( .A(G140), .B(G128), .Z(n1053) );
XOR2_X1 U1013 ( .A(n1270), .B(n1271), .Z(n1265) );
NOR2_X1 U1014 ( .A1(KEYINPUT58), .A2(n1272), .ZN(n1271) );
XOR2_X1 U1015 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR2_X1 U1016 ( .A1(KEYINPUT33), .A2(n1275), .ZN(n1274) );
NAND2_X1 U1017 ( .A1(n1222), .A2(G221), .ZN(n1273) );
NOR2_X1 U1018 ( .A1(n1264), .A2(G953), .ZN(n1222) );
INV_X1 U1019 ( .A(G234), .ZN(n1264) );
XOR2_X1 U1020 ( .A(G146), .B(n1117), .Z(n1270) );
INV_X1 U1021 ( .A(G110), .ZN(n1117) );
NAND2_X1 U1022 ( .A1(G217), .A2(G902), .ZN(n1260) );
NOR2_X1 U1023 ( .A1(n1031), .A2(n1034), .ZN(n1199) );
NOR2_X1 U1024 ( .A1(n1276), .A2(G472), .ZN(n1034) );
AND2_X1 U1025 ( .A1(n1276), .A2(G472), .ZN(n1031) );
NAND3_X1 U1026 ( .A1(n1277), .A2(n1278), .A3(n1141), .ZN(n1276) );
INV_X1 U1027 ( .A(G902), .ZN(n1141) );
NAND2_X1 U1028 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U1029 ( .A(KEYINPUT63), .ZN(n1280) );
XOR2_X1 U1030 ( .A(n1281), .B(n1282), .Z(n1279) );
NOR2_X1 U1031 ( .A1(KEYINPUT5), .A2(n1092), .ZN(n1281) );
NAND3_X1 U1032 ( .A1(n1283), .A2(n1096), .A3(KEYINPUT63), .ZN(n1277) );
INV_X1 U1033 ( .A(n1092), .ZN(n1096) );
XOR2_X1 U1034 ( .A(n1284), .B(G101), .Z(n1092) );
NAND2_X1 U1035 ( .A1(n1212), .A2(G210), .ZN(n1284) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1212) );
XOR2_X1 U1037 ( .A(KEYINPUT5), .B(n1282), .Z(n1283) );
XOR2_X1 U1038 ( .A(n1285), .B(n1105), .Z(n1282) );
XNOR2_X1 U1039 ( .A(n1259), .B(n1228), .ZN(n1105) );
XNOR2_X1 U1040 ( .A(n1051), .B(n1120), .ZN(n1228) );
NAND2_X1 U1041 ( .A1(KEYINPUT10), .A2(n1052), .ZN(n1120) );
XNOR2_X1 U1042 ( .A(G134), .B(KEYINPUT62), .ZN(n1052) );
XOR2_X1 U1043 ( .A(n1210), .B(n1275), .Z(n1051) );
INV_X1 U1044 ( .A(n1113), .ZN(n1275) );
XNOR2_X1 U1045 ( .A(G137), .B(KEYINPUT55), .ZN(n1113) );
XOR2_X1 U1046 ( .A(n1183), .B(n1132), .Z(n1210) );
XOR2_X1 U1047 ( .A(G143), .B(G146), .Z(n1132) );
INV_X1 U1048 ( .A(G131), .ZN(n1183) );
NOR2_X1 U1049 ( .A1(KEYINPUT59), .A2(G128), .ZN(n1259) );
INV_X1 U1050 ( .A(n1106), .ZN(n1285) );
XNOR2_X1 U1051 ( .A(G113), .B(n1286), .ZN(n1106) );
XOR2_X1 U1052 ( .A(G119), .B(G116), .Z(n1286) );
endmodule


