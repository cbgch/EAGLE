//Key = 1010001100100011101111010010010110001001100001110000111100000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
n1457, n1458, n1459, n1460, n1461;

XOR2_X1 U802 ( .A(G107), .B(n1107), .Z(G9) );
NOR2_X1 U803 ( .A1(n1108), .A2(n1109), .ZN(G75) );
NOR3_X1 U804 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
INV_X1 U805 ( .A(G952), .ZN(n1111) );
NAND3_X1 U806 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1110) );
NAND2_X1 U807 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U808 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U809 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NAND2_X1 U810 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NAND2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1123) );
NAND2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
INV_X1 U816 ( .A(n1135), .ZN(n1131) );
NAND3_X1 U817 ( .A1(n1129), .A2(n1136), .A3(n1125), .ZN(n1118) );
NAND2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U819 ( .A1(n1122), .A2(n1139), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U822 ( .A1(n1120), .A2(n1144), .ZN(n1137) );
NAND2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
INV_X1 U825 ( .A(n1149), .ZN(n1116) );
NOR3_X1 U826 ( .A1(n1150), .A2(G953), .A3(n1151), .ZN(n1108) );
INV_X1 U827 ( .A(n1113), .ZN(n1151) );
NAND4_X1 U828 ( .A1(n1152), .A2(n1129), .A3(n1153), .A4(n1154), .ZN(n1113) );
NOR4_X1 U829 ( .A1(n1147), .A2(n1133), .A3(n1155), .A4(n1156), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U831 ( .A(n1159), .B(KEYINPUT18), .ZN(n1155) );
NOR4_X1 U832 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1153) );
AND2_X1 U833 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1166), .ZN(n1162) );
NOR2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U836 ( .A1(KEYINPUT28), .A2(n1165), .ZN(n1168) );
NOR2_X1 U837 ( .A1(n1169), .A2(KEYINPUT44), .ZN(n1165) );
AND2_X1 U838 ( .A1(n1170), .A2(KEYINPUT28), .ZN(n1167) );
INV_X1 U839 ( .A(n1171), .ZN(n1164) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1161) );
NOR2_X1 U841 ( .A1(KEYINPUT59), .A2(n1174), .ZN(n1172) );
XNOR2_X1 U842 ( .A(KEYINPUT8), .B(n1157), .ZN(n1174) );
AND3_X1 U843 ( .A1(n1173), .A2(n1158), .A3(n1157), .ZN(n1160) );
INV_X1 U844 ( .A(KEYINPUT59), .ZN(n1158) );
XNOR2_X1 U845 ( .A(n1175), .B(KEYINPUT12), .ZN(n1173) );
INV_X1 U846 ( .A(n1143), .ZN(n1152) );
XNOR2_X1 U847 ( .A(G952), .B(KEYINPUT36), .ZN(n1150) );
XOR2_X1 U848 ( .A(n1176), .B(n1177), .Z(G72) );
XOR2_X1 U849 ( .A(n1178), .B(n1179), .Z(n1177) );
NAND2_X1 U850 ( .A1(n1114), .A2(n1180), .ZN(n1179) );
NAND3_X1 U851 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1178) );
INV_X1 U852 ( .A(n1184), .ZN(n1183) );
NAND2_X1 U853 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1185) );
NOR2_X1 U855 ( .A1(KEYINPUT25), .A2(n1189), .ZN(n1188) );
NAND2_X1 U856 ( .A1(n1190), .A2(n1191), .ZN(n1181) );
XOR2_X1 U857 ( .A(n1187), .B(n1192), .Z(n1191) );
NOR2_X1 U858 ( .A1(KEYINPUT25), .A2(n1193), .ZN(n1192) );
INV_X1 U859 ( .A(n1189), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1194), .A2(n1195), .ZN(n1187) );
NAND2_X1 U861 ( .A1(G125), .A2(G140), .ZN(n1194) );
INV_X1 U862 ( .A(n1186), .ZN(n1190) );
NAND2_X1 U863 ( .A1(n1196), .A2(KEYINPUT2), .ZN(n1186) );
XNOR2_X1 U864 ( .A(n1197), .B(n1198), .ZN(n1196) );
NAND3_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1197) );
NAND2_X1 U866 ( .A1(G134), .A2(n1202), .ZN(n1201) );
OR3_X1 U867 ( .A1(n1202), .A2(n1203), .A3(G137), .ZN(n1200) );
INV_X1 U868 ( .A(KEYINPUT19), .ZN(n1202) );
NAND2_X1 U869 ( .A1(G137), .A2(n1203), .ZN(n1199) );
NAND2_X1 U870 ( .A1(KEYINPUT15), .A2(n1204), .ZN(n1203) );
NOR2_X1 U871 ( .A1(n1205), .A2(n1114), .ZN(n1176) );
AND2_X1 U872 ( .A1(G227), .A2(G900), .ZN(n1205) );
XOR2_X1 U873 ( .A(n1206), .B(n1207), .Z(G69) );
XOR2_X1 U874 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U875 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U876 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U877 ( .A(n1214), .B(n1215), .Z(n1212) );
NOR2_X1 U878 ( .A1(G898), .A2(n1216), .ZN(n1210) );
NAND2_X1 U879 ( .A1(n1114), .A2(n1217), .ZN(n1208) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U881 ( .A1(G953), .A2(n1220), .ZN(n1206) );
NAND2_X1 U882 ( .A1(G898), .A2(G224), .ZN(n1220) );
NOR2_X1 U883 ( .A1(n1221), .A2(n1222), .ZN(G66) );
NOR2_X1 U884 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U885 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U886 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U887 ( .A1(n1229), .A2(n1230), .ZN(n1225) );
INV_X1 U888 ( .A(KEYINPUT47), .ZN(n1230) );
XOR2_X1 U889 ( .A(n1231), .B(KEYINPUT32), .Z(n1229) );
NOR2_X1 U890 ( .A1(KEYINPUT47), .A2(n1232), .ZN(n1223) );
XNOR2_X1 U891 ( .A(KEYINPUT32), .B(n1231), .ZN(n1232) );
NOR2_X1 U892 ( .A1(n1221), .A2(n1233), .ZN(G63) );
XOR2_X1 U893 ( .A(n1234), .B(n1235), .Z(n1233) );
AND2_X1 U894 ( .A1(G478), .A2(n1236), .ZN(n1235) );
NAND2_X1 U895 ( .A1(KEYINPUT52), .A2(n1237), .ZN(n1234) );
NOR2_X1 U896 ( .A1(n1221), .A2(n1238), .ZN(G60) );
XOR2_X1 U897 ( .A(n1239), .B(n1240), .Z(n1238) );
AND2_X1 U898 ( .A1(G475), .A2(n1236), .ZN(n1240) );
INV_X1 U899 ( .A(n1228), .ZN(n1236) );
XNOR2_X1 U900 ( .A(G104), .B(n1241), .ZN(G6) );
NAND2_X1 U901 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U902 ( .A(n1244), .B(KEYINPUT29), .Z(n1242) );
NOR2_X1 U903 ( .A1(n1221), .A2(n1245), .ZN(G57) );
XOR2_X1 U904 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U905 ( .A(n1248), .B(n1249), .Z(n1247) );
NOR3_X1 U906 ( .A1(n1228), .A2(KEYINPUT50), .A3(n1250), .ZN(n1248) );
NOR3_X1 U907 ( .A1(n1221), .A2(n1251), .A3(n1252), .ZN(G54) );
NOR2_X1 U908 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U909 ( .A(n1255), .ZN(n1254) );
NOR2_X1 U910 ( .A1(n1256), .A2(n1257), .ZN(n1253) );
NOR2_X1 U911 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U912 ( .A(KEYINPUT45), .ZN(n1259) );
NOR2_X1 U913 ( .A1(KEYINPUT45), .A2(n1260), .ZN(n1256) );
NOR2_X1 U914 ( .A1(n1255), .A2(n1261), .ZN(n1251) );
NOR2_X1 U915 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR2_X1 U916 ( .A1(n1258), .A2(n1264), .ZN(n1263) );
INV_X1 U917 ( .A(KEYINPUT35), .ZN(n1264) );
NAND2_X1 U918 ( .A1(n1265), .A2(n1266), .ZN(n1258) );
NAND2_X1 U919 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U920 ( .A1(n1269), .A2(n1270), .ZN(n1265) );
NOR2_X1 U921 ( .A1(KEYINPUT35), .A2(n1260), .ZN(n1262) );
NAND2_X1 U922 ( .A1(n1271), .A2(n1272), .ZN(n1260) );
NAND2_X1 U923 ( .A1(n1270), .A2(n1268), .ZN(n1272) );
INV_X1 U924 ( .A(n1269), .ZN(n1268) );
NAND2_X1 U925 ( .A1(n1267), .A2(n1269), .ZN(n1271) );
XOR2_X1 U926 ( .A(G110), .B(n1273), .Z(n1269) );
XOR2_X1 U927 ( .A(n1270), .B(KEYINPUT21), .Z(n1267) );
NOR2_X1 U928 ( .A1(n1228), .A2(n1157), .ZN(n1270) );
XNOR2_X1 U929 ( .A(n1274), .B(n1275), .ZN(n1255) );
NAND2_X1 U930 ( .A1(n1276), .A2(n1277), .ZN(n1274) );
OR2_X1 U931 ( .A1(n1278), .A2(n1189), .ZN(n1277) );
XOR2_X1 U932 ( .A(n1279), .B(KEYINPUT57), .Z(n1276) );
NAND2_X1 U933 ( .A1(n1189), .A2(n1278), .ZN(n1279) );
NOR2_X1 U934 ( .A1(n1221), .A2(n1280), .ZN(G51) );
XOR2_X1 U935 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U936 ( .A(n1283), .B(n1284), .ZN(n1282) );
NOR2_X1 U937 ( .A1(n1171), .A2(n1228), .ZN(n1283) );
NAND2_X1 U938 ( .A1(G902), .A2(n1112), .ZN(n1228) );
NAND3_X1 U939 ( .A1(n1218), .A2(n1285), .A3(n1286), .ZN(n1112) );
INV_X1 U940 ( .A(n1180), .ZN(n1286) );
NAND4_X1 U941 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1180) );
NOR4_X1 U942 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1290) );
NOR2_X1 U943 ( .A1(n1295), .A2(n1296), .ZN(n1289) );
NAND2_X1 U944 ( .A1(n1243), .A2(n1297), .ZN(n1288) );
NAND2_X1 U945 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
OR2_X1 U946 ( .A1(n1300), .A2(KEYINPUT48), .ZN(n1299) );
XOR2_X1 U947 ( .A(n1301), .B(KEYINPUT3), .Z(n1298) );
NAND3_X1 U948 ( .A1(KEYINPUT48), .A2(n1302), .A3(n1145), .ZN(n1287) );
INV_X1 U949 ( .A(n1300), .ZN(n1302) );
XNOR2_X1 U950 ( .A(KEYINPUT31), .B(n1219), .ZN(n1285) );
AND4_X1 U951 ( .A1(n1303), .A2(n1304), .A3(n1305), .A4(n1306), .ZN(n1218) );
NOR4_X1 U952 ( .A1(n1107), .A2(n1307), .A3(n1308), .A4(n1309), .ZN(n1306) );
INV_X1 U953 ( .A(n1310), .ZN(n1307) );
AND3_X1 U954 ( .A1(n1311), .A2(n1120), .A3(n1312), .ZN(n1107) );
OR2_X1 U955 ( .A1(n1244), .A2(n1145), .ZN(n1305) );
NAND4_X1 U956 ( .A1(n1313), .A2(n1120), .A3(n1135), .A4(n1314), .ZN(n1244) );
XOR2_X1 U957 ( .A(n1315), .B(n1316), .Z(n1281) );
XNOR2_X1 U958 ( .A(G125), .B(n1317), .ZN(n1316) );
NOR2_X1 U959 ( .A1(KEYINPUT60), .A2(n1318), .ZN(n1317) );
NAND2_X1 U960 ( .A1(KEYINPUT7), .A2(n1319), .ZN(n1315) );
NOR2_X1 U961 ( .A1(n1114), .A2(G952), .ZN(n1221) );
XNOR2_X1 U962 ( .A(n1320), .B(n1296), .ZN(G48) );
AND3_X1 U963 ( .A1(n1243), .A2(n1159), .A3(n1321), .ZN(n1296) );
XOR2_X1 U964 ( .A(G143), .B(n1322), .Z(G45) );
NOR2_X1 U965 ( .A1(n1145), .A2(n1300), .ZN(n1322) );
NAND3_X1 U966 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1300) );
XOR2_X1 U967 ( .A(n1326), .B(n1295), .Z(G42) );
AND3_X1 U968 ( .A1(n1142), .A2(n1122), .A3(n1321), .ZN(n1295) );
AND3_X1 U969 ( .A1(n1313), .A2(n1143), .A3(n1324), .ZN(n1321) );
XNOR2_X1 U970 ( .A(G140), .B(KEYINPUT55), .ZN(n1326) );
XOR2_X1 U971 ( .A(G137), .B(n1294), .Z(G39) );
AND3_X1 U972 ( .A1(n1324), .A2(n1122), .A3(n1327), .ZN(n1294) );
AND3_X1 U973 ( .A1(n1129), .A2(n1159), .A3(n1143), .ZN(n1327) );
XNOR2_X1 U974 ( .A(G134), .B(n1328), .ZN(G36) );
NOR2_X1 U975 ( .A1(n1293), .A2(KEYINPUT27), .ZN(n1328) );
AND2_X1 U976 ( .A1(n1329), .A2(n1311), .ZN(n1293) );
XOR2_X1 U977 ( .A(n1292), .B(n1330), .Z(G33) );
NOR2_X1 U978 ( .A1(KEYINPUT13), .A2(n1198), .ZN(n1330) );
AND2_X1 U979 ( .A1(n1329), .A2(n1313), .ZN(n1292) );
AND3_X1 U980 ( .A1(n1324), .A2(n1122), .A3(n1323), .ZN(n1329) );
NOR2_X1 U981 ( .A1(n1331), .A2(n1147), .ZN(n1122) );
XNOR2_X1 U982 ( .A(n1332), .B(n1333), .ZN(G30) );
NOR2_X1 U983 ( .A1(n1145), .A2(n1301), .ZN(n1333) );
NAND4_X1 U984 ( .A1(n1324), .A2(n1311), .A3(n1143), .A4(n1159), .ZN(n1301) );
AND2_X1 U985 ( .A1(n1135), .A2(n1334), .ZN(n1324) );
INV_X1 U986 ( .A(n1243), .ZN(n1145) );
XNOR2_X1 U987 ( .A(G101), .B(n1303), .ZN(G3) );
NAND3_X1 U988 ( .A1(n1129), .A2(n1312), .A3(n1323), .ZN(n1303) );
XNOR2_X1 U989 ( .A(G125), .B(n1335), .ZN(G27) );
NAND2_X1 U990 ( .A1(KEYINPUT20), .A2(n1291), .ZN(n1335) );
AND4_X1 U991 ( .A1(n1143), .A2(n1334), .A3(n1243), .A4(n1336), .ZN(n1291) );
NOR3_X1 U992 ( .A1(n1127), .A2(n1337), .A3(n1159), .ZN(n1336) );
INV_X1 U993 ( .A(n1313), .ZN(n1127) );
NAND2_X1 U994 ( .A1(n1149), .A2(n1338), .ZN(n1334) );
NAND3_X1 U995 ( .A1(G902), .A2(n1339), .A3(n1184), .ZN(n1338) );
NOR2_X1 U996 ( .A1(n1216), .A2(G900), .ZN(n1184) );
XNOR2_X1 U997 ( .A(n1304), .B(n1340), .ZN(G24) );
NOR2_X1 U998 ( .A1(KEYINPUT41), .A2(n1341), .ZN(n1340) );
NAND3_X1 U999 ( .A1(n1325), .A2(n1120), .A3(n1342), .ZN(n1304) );
NOR2_X1 U1000 ( .A1(n1159), .A2(n1143), .ZN(n1120) );
AND2_X1 U1001 ( .A1(n1343), .A2(n1344), .ZN(n1325) );
XNOR2_X1 U1002 ( .A(n1345), .B(KEYINPUT23), .ZN(n1343) );
XNOR2_X1 U1003 ( .A(G119), .B(n1346), .ZN(G21) );
NOR2_X1 U1004 ( .A1(n1309), .A2(KEYINPUT34), .ZN(n1346) );
AND4_X1 U1005 ( .A1(n1342), .A2(n1129), .A3(n1143), .A4(n1159), .ZN(n1309) );
XOR2_X1 U1006 ( .A(n1347), .B(n1348), .Z(G18) );
NOR2_X1 U1007 ( .A1(KEYINPUT30), .A2(n1349), .ZN(n1348) );
NAND2_X1 U1008 ( .A1(n1350), .A2(n1351), .ZN(n1347) );
NAND4_X1 U1009 ( .A1(n1352), .A2(n1337), .A3(n1353), .A4(n1354), .ZN(n1351) );
NOR2_X1 U1010 ( .A1(n1128), .A2(n1140), .ZN(n1353) );
INV_X1 U1011 ( .A(n1311), .ZN(n1128) );
OR2_X1 U1012 ( .A1(n1219), .A2(n1354), .ZN(n1350) );
INV_X1 U1013 ( .A(KEYINPUT53), .ZN(n1354) );
NAND3_X1 U1014 ( .A1(n1323), .A2(n1311), .A3(n1342), .ZN(n1219) );
NOR2_X1 U1015 ( .A1(n1345), .A2(n1355), .ZN(n1311) );
INV_X1 U1016 ( .A(n1344), .ZN(n1355) );
XOR2_X1 U1017 ( .A(G113), .B(n1308), .Z(G15) );
AND3_X1 U1018 ( .A1(n1323), .A2(n1313), .A3(n1342), .ZN(n1308) );
AND2_X1 U1019 ( .A1(n1125), .A2(n1352), .ZN(n1342) );
INV_X1 U1020 ( .A(n1337), .ZN(n1125) );
NAND2_X1 U1021 ( .A1(n1134), .A2(n1356), .ZN(n1337) );
NOR2_X1 U1022 ( .A1(n1344), .A2(n1357), .ZN(n1313) );
INV_X1 U1023 ( .A(n1345), .ZN(n1357) );
INV_X1 U1024 ( .A(n1140), .ZN(n1323) );
NAND2_X1 U1025 ( .A1(n1358), .A2(n1159), .ZN(n1140) );
XNOR2_X1 U1026 ( .A(n1143), .B(KEYINPUT62), .ZN(n1358) );
XNOR2_X1 U1027 ( .A(G110), .B(n1310), .ZN(G12) );
NAND4_X1 U1028 ( .A1(n1129), .A2(n1312), .A3(n1142), .A4(n1143), .ZN(n1310) );
XOR2_X1 U1029 ( .A(n1359), .B(n1227), .Z(n1143) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1360), .ZN(n1227) );
NAND2_X1 U1031 ( .A1(n1231), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1032 ( .A(n1362), .B(n1363), .Z(n1231) );
XOR2_X1 U1033 ( .A(n1364), .B(n1365), .Z(n1363) );
XNOR2_X1 U1034 ( .A(G137), .B(G110), .ZN(n1365) );
NAND2_X1 U1035 ( .A1(KEYINPUT39), .A2(n1366), .ZN(n1364) );
XNOR2_X1 U1036 ( .A(n1332), .B(G119), .ZN(n1366) );
XOR2_X1 U1037 ( .A(n1367), .B(n1368), .Z(n1362) );
NOR2_X1 U1038 ( .A1(KEYINPUT37), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1039 ( .A(n1370), .B(n1371), .Z(n1367) );
AND3_X1 U1040 ( .A1(G221), .A2(n1114), .A3(G234), .ZN(n1371) );
NAND2_X1 U1041 ( .A1(n1372), .A2(n1373), .ZN(n1370) );
NAND2_X1 U1042 ( .A1(G125), .A2(n1374), .ZN(n1373) );
OR2_X1 U1043 ( .A1(KEYINPUT11), .A2(G140), .ZN(n1374) );
OR2_X1 U1044 ( .A1(n1195), .A2(KEYINPUT11), .ZN(n1372) );
INV_X1 U1045 ( .A(n1159), .ZN(n1142) );
XOR2_X1 U1046 ( .A(n1375), .B(n1250), .Z(n1159) );
INV_X1 U1047 ( .A(G472), .ZN(n1250) );
NAND2_X1 U1048 ( .A1(n1376), .A2(n1361), .ZN(n1375) );
XNOR2_X1 U1049 ( .A(n1246), .B(n1249), .ZN(n1376) );
XNOR2_X1 U1050 ( .A(n1377), .B(G101), .ZN(n1249) );
NAND2_X1 U1051 ( .A1(n1378), .A2(G210), .ZN(n1377) );
XNOR2_X1 U1052 ( .A(n1379), .B(n1380), .ZN(n1246) );
XNOR2_X1 U1053 ( .A(n1284), .B(n1381), .ZN(n1380) );
XNOR2_X1 U1054 ( .A(n1275), .B(KEYINPUT1), .ZN(n1379) );
AND2_X1 U1055 ( .A1(n1135), .A2(n1352), .ZN(n1312) );
AND2_X1 U1056 ( .A1(n1243), .A2(n1314), .ZN(n1352) );
NAND2_X1 U1057 ( .A1(n1149), .A2(n1382), .ZN(n1314) );
OR4_X1 U1058 ( .A1(n1216), .A2(n1361), .A3(n1383), .A4(G898), .ZN(n1382) );
INV_X1 U1059 ( .A(n1339), .ZN(n1383) );
XOR2_X1 U1060 ( .A(G953), .B(KEYINPUT46), .Z(n1216) );
NAND3_X1 U1061 ( .A1(n1339), .A2(n1114), .A3(G952), .ZN(n1149) );
NAND2_X1 U1062 ( .A1(G237), .A2(G234), .ZN(n1339) );
NOR2_X1 U1063 ( .A1(n1148), .A2(n1147), .ZN(n1243) );
AND2_X1 U1064 ( .A1(G214), .A2(n1384), .ZN(n1147) );
INV_X1 U1065 ( .A(n1331), .ZN(n1148) );
XNOR2_X1 U1066 ( .A(n1169), .B(n1171), .ZN(n1331) );
NAND2_X1 U1067 ( .A1(G210), .A2(n1384), .ZN(n1171) );
NAND2_X1 U1068 ( .A1(n1361), .A2(n1385), .ZN(n1384) );
INV_X1 U1069 ( .A(G237), .ZN(n1385) );
INV_X1 U1070 ( .A(n1170), .ZN(n1169) );
NAND2_X1 U1071 ( .A1(n1386), .A2(n1361), .ZN(n1170) );
XOR2_X1 U1072 ( .A(n1387), .B(n1388), .Z(n1386) );
XNOR2_X1 U1073 ( .A(n1389), .B(n1390), .ZN(n1388) );
NOR2_X1 U1074 ( .A1(KEYINPUT33), .A2(n1284), .ZN(n1390) );
XOR2_X1 U1075 ( .A(n1391), .B(n1392), .Z(n1284) );
NOR2_X1 U1076 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
NOR2_X1 U1077 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
NOR2_X1 U1078 ( .A1(n1397), .A2(n1398), .ZN(n1393) );
NOR2_X1 U1079 ( .A1(G146), .A2(n1395), .ZN(n1397) );
INV_X1 U1080 ( .A(KEYINPUT26), .ZN(n1395) );
XNOR2_X1 U1081 ( .A(G128), .B(KEYINPUT38), .ZN(n1391) );
XOR2_X1 U1082 ( .A(n1318), .B(n1319), .Z(n1387) );
AND2_X1 U1083 ( .A1(G224), .A2(n1114), .ZN(n1319) );
XOR2_X1 U1084 ( .A(n1399), .B(n1215), .Z(n1318) );
XNOR2_X1 U1085 ( .A(n1341), .B(G110), .ZN(n1215) );
XOR2_X1 U1086 ( .A(n1400), .B(KEYINPUT14), .Z(n1399) );
NAND3_X1 U1087 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n1400) );
NAND2_X1 U1088 ( .A1(KEYINPUT51), .A2(n1214), .ZN(n1403) );
NAND3_X1 U1089 ( .A1(n1404), .A2(n1405), .A3(n1213), .ZN(n1402) );
INV_X1 U1090 ( .A(KEYINPUT51), .ZN(n1405) );
OR2_X1 U1091 ( .A1(n1213), .A2(n1404), .ZN(n1401) );
NOR2_X1 U1092 ( .A1(KEYINPUT4), .A2(n1214), .ZN(n1404) );
XNOR2_X1 U1093 ( .A(n1381), .B(n1406), .ZN(n1214) );
XOR2_X1 U1094 ( .A(KEYINPUT5), .B(KEYINPUT40), .Z(n1406) );
XOR2_X1 U1095 ( .A(G113), .B(n1407), .Z(n1381) );
XNOR2_X1 U1096 ( .A(G119), .B(n1349), .ZN(n1407) );
XOR2_X1 U1097 ( .A(G101), .B(n1408), .Z(n1213) );
NOR2_X1 U1098 ( .A1(n1134), .A2(n1133), .ZN(n1135) );
INV_X1 U1099 ( .A(n1356), .ZN(n1133) );
NAND2_X1 U1100 ( .A1(G221), .A2(n1360), .ZN(n1356) );
NAND2_X1 U1101 ( .A1(G234), .A2(n1361), .ZN(n1360) );
XNOR2_X1 U1102 ( .A(n1175), .B(n1157), .ZN(n1134) );
INV_X1 U1103 ( .A(G469), .ZN(n1157) );
NAND2_X1 U1104 ( .A1(n1361), .A2(n1409), .ZN(n1175) );
NAND2_X1 U1105 ( .A1(n1410), .A2(n1411), .ZN(n1409) );
NAND2_X1 U1106 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
XOR2_X1 U1107 ( .A(n1414), .B(KEYINPUT58), .Z(n1410) );
OR2_X1 U1108 ( .A1(n1413), .A2(n1412), .ZN(n1414) );
NAND2_X1 U1109 ( .A1(n1415), .A2(n1416), .ZN(n1412) );
OR2_X1 U1110 ( .A1(n1417), .A2(n1273), .ZN(n1416) );
NAND2_X1 U1111 ( .A1(n1418), .A2(n1417), .ZN(n1415) );
INV_X1 U1112 ( .A(G110), .ZN(n1417) );
XNOR2_X1 U1113 ( .A(n1273), .B(KEYINPUT63), .ZN(n1418) );
XOR2_X1 U1114 ( .A(G140), .B(n1419), .Z(n1273) );
AND2_X1 U1115 ( .A1(n1114), .A2(G227), .ZN(n1419) );
XNOR2_X1 U1116 ( .A(n1420), .B(n1275), .ZN(n1413) );
XOR2_X1 U1117 ( .A(n1421), .B(n1198), .Z(n1275) );
NAND2_X1 U1118 ( .A1(KEYINPUT16), .A2(n1422), .ZN(n1421) );
XNOR2_X1 U1119 ( .A(G137), .B(n1204), .ZN(n1422) );
NAND2_X1 U1120 ( .A1(n1423), .A2(KEYINPUT0), .ZN(n1420) );
XNOR2_X1 U1121 ( .A(n1278), .B(n1189), .ZN(n1423) );
XOR2_X1 U1122 ( .A(G128), .B(n1424), .Z(n1189) );
NOR2_X1 U1123 ( .A1(n1425), .A2(n1426), .ZN(n1424) );
XOR2_X1 U1124 ( .A(KEYINPUT22), .B(n1427), .Z(n1426) );
NOR2_X1 U1125 ( .A1(n1398), .A2(n1320), .ZN(n1427) );
INV_X1 U1126 ( .A(n1396), .ZN(n1425) );
NAND2_X1 U1127 ( .A1(n1398), .A2(n1320), .ZN(n1396) );
XOR2_X1 U1128 ( .A(G143), .B(KEYINPUT42), .Z(n1398) );
XNOR2_X1 U1129 ( .A(n1428), .B(n1408), .ZN(n1278) );
XOR2_X1 U1130 ( .A(G104), .B(G107), .Z(n1408) );
XNOR2_X1 U1131 ( .A(KEYINPUT54), .B(n1429), .ZN(n1428) );
NOR2_X1 U1132 ( .A1(KEYINPUT17), .A2(n1430), .ZN(n1429) );
INV_X1 U1133 ( .A(G101), .ZN(n1430) );
NOR2_X1 U1134 ( .A1(n1344), .A2(n1345), .ZN(n1129) );
XOR2_X1 U1135 ( .A(G475), .B(n1431), .Z(n1345) );
NOR2_X1 U1136 ( .A1(G902), .A2(n1239), .ZN(n1431) );
NAND3_X1 U1137 ( .A1(n1432), .A2(n1433), .A3(n1434), .ZN(n1239) );
NAND2_X1 U1138 ( .A1(n1435), .A2(n1436), .ZN(n1434) );
INV_X1 U1139 ( .A(KEYINPUT6), .ZN(n1436) );
NAND3_X1 U1140 ( .A1(KEYINPUT6), .A2(n1437), .A3(n1438), .ZN(n1433) );
OR2_X1 U1141 ( .A1(n1438), .A2(n1437), .ZN(n1432) );
NOR2_X1 U1142 ( .A1(KEYINPUT9), .A2(n1435), .ZN(n1437) );
XOR2_X1 U1143 ( .A(G104), .B(n1439), .Z(n1435) );
XNOR2_X1 U1144 ( .A(n1341), .B(G113), .ZN(n1439) );
INV_X1 U1145 ( .A(G122), .ZN(n1341) );
XOR2_X1 U1146 ( .A(n1440), .B(n1441), .Z(n1438) );
XOR2_X1 U1147 ( .A(n1442), .B(n1369), .Z(n1441) );
XNOR2_X1 U1148 ( .A(n1320), .B(KEYINPUT24), .ZN(n1369) );
INV_X1 U1149 ( .A(G146), .ZN(n1320) );
AND3_X1 U1150 ( .A1(n1378), .A2(n1443), .A3(G214), .ZN(n1442) );
INV_X1 U1151 ( .A(KEYINPUT56), .ZN(n1443) );
NOR2_X1 U1152 ( .A1(G953), .A2(G237), .ZN(n1378) );
XOR2_X1 U1153 ( .A(n1444), .B(n1445), .Z(n1440) );
XNOR2_X1 U1154 ( .A(G143), .B(n1198), .ZN(n1445) );
INV_X1 U1155 ( .A(G131), .ZN(n1198) );
NAND3_X1 U1156 ( .A1(n1446), .A2(n1447), .A3(n1195), .ZN(n1444) );
NAND2_X1 U1157 ( .A1(n1448), .A2(n1389), .ZN(n1195) );
NAND2_X1 U1158 ( .A1(KEYINPUT61), .A2(n1448), .ZN(n1447) );
OR3_X1 U1159 ( .A1(n1389), .A2(KEYINPUT61), .A3(n1448), .ZN(n1446) );
INV_X1 U1160 ( .A(G140), .ZN(n1448) );
INV_X1 U1161 ( .A(G125), .ZN(n1389) );
XOR2_X1 U1162 ( .A(G478), .B(n1449), .Z(n1344) );
AND2_X1 U1163 ( .A1(n1237), .A2(n1361), .ZN(n1449) );
INV_X1 U1164 ( .A(G902), .ZN(n1361) );
NAND2_X1 U1165 ( .A1(n1450), .A2(n1451), .ZN(n1237) );
NAND2_X1 U1166 ( .A1(n1452), .A2(n1453), .ZN(n1451) );
NAND3_X1 U1167 ( .A1(G234), .A2(n1114), .A3(G217), .ZN(n1453) );
INV_X1 U1168 ( .A(n1454), .ZN(n1452) );
XOR2_X1 U1169 ( .A(KEYINPUT10), .B(n1455), .Z(n1450) );
AND4_X1 U1170 ( .A1(n1114), .A2(G234), .A3(G217), .A4(n1454), .ZN(n1455) );
XOR2_X1 U1171 ( .A(n1456), .B(n1457), .Z(n1454) );
XOR2_X1 U1172 ( .A(n1458), .B(n1459), .Z(n1457) );
XNOR2_X1 U1173 ( .A(n1349), .B(G107), .ZN(n1459) );
INV_X1 U1174 ( .A(G116), .ZN(n1349) );
XNOR2_X1 U1175 ( .A(n1332), .B(G122), .ZN(n1458) );
INV_X1 U1176 ( .A(G128), .ZN(n1332) );
XOR2_X1 U1177 ( .A(n1460), .B(n1461), .Z(n1456) );
XNOR2_X1 U1178 ( .A(G143), .B(n1204), .ZN(n1461) );
INV_X1 U1179 ( .A(G134), .ZN(n1204) );
XNOR2_X1 U1180 ( .A(KEYINPUT49), .B(KEYINPUT43), .ZN(n1460) );
INV_X1 U1181 ( .A(G953), .ZN(n1114) );
endmodule


