//Key = 11101001001100110111110011100
module c1355 ( G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, 
        G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, 
        G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, 
        G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, 
        G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, 
        G233gat, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat, 
        G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat, 
        G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat, 
        G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat, 
        G1352gat, G1353gat, G1354gat, G1355gat );
  input G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
         G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
         G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
         G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
         G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat,
         G231gat, G232gat, G233gat, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
         G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
         G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
         G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
         G1352gat, G1353gat, G1354gat, G1355gat;
  wire   n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881;

  XOR2_X1 U556 ( .A(G218gat), .B(n705), .Z(G1355gat) );
  NOR2_X1 U557 ( .A1(n706), .A2(n707), .ZN(n705) );
  XOR2_X1 U558 ( .A(n708), .B(n709), .Z(G1354gat) );
  NOR2_X1 U559 ( .A1(n710), .A2(n707), .ZN(n709) );
  XOR2_X1 U560 ( .A(n711), .B(n712), .Z(G1353gat) );
  NOR2_X1 U561 ( .A1(n707), .A2(n713), .ZN(n712) );
  XOR2_X1 U562 ( .A(G197gat), .B(n714), .Z(G1352gat) );
  NOR2_X1 U563 ( .A1(n707), .A2(n715), .ZN(n714) );
  XOR2_X1 U564 ( .A(n716), .B(keyinput28), .Z(n707) );
  NAND4_X1 U565 ( .A1(n717), .A2(n718), .A3(n719), .A4(n720), .ZN(n716) );
  XOR2_X1 U566 ( .A(G190gat), .B(n721), .Z(G1351gat) );
  NOR2_X1 U567 ( .A1(n706), .A2(n722), .ZN(n721) );
  XOR2_X1 U568 ( .A(n723), .B(n724), .Z(G1350gat) );
  NOR2_X1 U569 ( .A1(n710), .A2(n722), .ZN(n724) );
  XOR2_X1 U570 ( .A(n725), .B(n726), .Z(G1349gat) );
  NOR2_X1 U571 ( .A1(n722), .A2(n713), .ZN(n726) );
  XOR2_X1 U572 ( .A(n727), .B(n728), .Z(G1348gat) );
  NOR2_X1 U573 ( .A1(n722), .A2(n715), .ZN(n727) );
  XOR2_X1 U574 ( .A(n729), .B(keyinput27), .Z(n722) );
  NAND4_X1 U575 ( .A1(n730), .A2(n720), .A3(n731), .A4(n732), .ZN(n729) );
  NOR2_X1 U576 ( .A1(n733), .A2(n719), .ZN(n732) );
  XNOR2_X1 U577 ( .A(G162gat), .B(n734), .ZN(G1347gat) );
  NAND2_X1 U578 ( .A1(n735), .A2(n736), .ZN(n734) );
  XOR2_X1 U579 ( .A(n737), .B(n738), .Z(G1346gat) );
  NAND2_X1 U580 ( .A1(n735), .A2(n739), .ZN(n737) );
  XOR2_X1 U581 ( .A(n740), .B(n741), .Z(G1345gat) );
  NAND2_X1 U582 ( .A1(n735), .A2(n742), .ZN(n740) );
  XOR2_X1 U583 ( .A(n743), .B(n744), .Z(G1344gat) );
  NAND2_X1 U584 ( .A1(n735), .A2(n745), .ZN(n743) );
  XOR2_X1 U585 ( .A(n746), .B(keyinput26), .Z(n735) );
  NAND4_X1 U586 ( .A1(n719), .A2(n720), .A3(n747), .A4(n748), .ZN(n746) );
  NOR2_X1 U587 ( .A1(n718), .A2(n730), .ZN(n748) );
  XNOR2_X1 U588 ( .A(G134gat), .B(n749), .ZN(G1343gat) );
  NAND2_X1 U589 ( .A1(n750), .A2(n736), .ZN(n749) );
  XOR2_X1 U590 ( .A(n751), .B(n752), .Z(G1342gat) );
  NAND2_X1 U591 ( .A1(n750), .A2(n739), .ZN(n751) );
  XOR2_X1 U592 ( .A(n753), .B(n754), .Z(G1341gat) );
  NAND2_X1 U593 ( .A1(n750), .A2(n742), .ZN(n753) );
  XOR2_X1 U594 ( .A(n755), .B(n756), .Z(G1340gat) );
  NAND2_X1 U595 ( .A1(n750), .A2(n745), .ZN(n755) );
  XOR2_X1 U596 ( .A(n757), .B(keyinput25), .Z(n750) );
  NAND4_X1 U597 ( .A1(n758), .A2(n759), .A3(n731), .A4(n720), .ZN(n757) );
  NAND2_X1 U598 ( .A1(n760), .A2(n761), .ZN(n720) );
  OR3_X1 U599 ( .A1(n742), .A2(n762), .A3(n736), .ZN(n761) );
  OR3_X1 U600 ( .A1(n745), .A2(n763), .A3(n739), .ZN(n760) );
  XNOR2_X1 U601 ( .A(G106gat), .B(n764), .ZN(G1339gat) );
  NAND2_X1 U602 ( .A1(n765), .A2(n747), .ZN(n764) );
  XOR2_X1 U603 ( .A(n766), .B(n767), .Z(G1338gat) );
  NAND2_X1 U604 ( .A1(n765), .A2(n768), .ZN(n767) );
  XOR2_X1 U605 ( .A(n769), .B(n770), .Z(G1337gat) );
  NAND2_X1 U606 ( .A1(n765), .A2(n730), .ZN(n769) );
  XOR2_X1 U607 ( .A(n771), .B(n772), .Z(G1336gat) );
  NAND2_X1 U608 ( .A1(n765), .A2(n733), .ZN(n771) );
  XOR2_X1 U609 ( .A(n773), .B(keyinput24), .Z(n765) );
  NAND4_X1 U610 ( .A1(n710), .A2(n763), .A3(n715), .A4(n774), .ZN(n773) );
  NOR2_X1 U611 ( .A1(n713), .A2(n706), .ZN(n763) );
  XOR2_X1 U612 ( .A(G78gat), .B(n775), .Z(G1335gat) );
  NOR2_X1 U613 ( .A1(n776), .A2(n731), .ZN(n775) );
  XOR2_X1 U614 ( .A(G71gat), .B(n777), .Z(G1334gat) );
  NOR2_X1 U615 ( .A1(n776), .A2(n719), .ZN(n777) );
  XNOR2_X1 U616 ( .A(n778), .B(n779), .ZN(G1333gat) );
  NOR2_X1 U617 ( .A1(n758), .A2(n776), .ZN(n778) );
  XOR2_X1 U618 ( .A(n780), .B(n781), .Z(G1332gat) );
  NOR2_X1 U619 ( .A1(n776), .A2(n718), .ZN(n780) );
  XOR2_X1 U620 ( .A(n782), .B(keyinput23), .Z(n776) );
  NAND4_X1 U621 ( .A1(n739), .A2(n774), .A3(n715), .A4(n783), .ZN(n782) );
  NOR2_X1 U622 ( .A1(n736), .A2(n713), .ZN(n783) );
  XOR2_X1 U623 ( .A(n784), .B(n785), .Z(G1331gat) );
  NOR2_X1 U624 ( .A1(n786), .A2(n731), .ZN(n784) );
  XOR2_X1 U625 ( .A(G43gat), .B(n787), .Z(G1330gat) );
  NOR2_X1 U626 ( .A1(n786), .A2(n719), .ZN(n787) );
  XOR2_X1 U627 ( .A(n788), .B(n789), .Z(G1329gat) );
  NOR2_X1 U628 ( .A1(n758), .A2(n786), .ZN(n789) );
  XOR2_X1 U629 ( .A(n790), .B(n791), .Z(G1328gat) );
  NOR2_X1 U630 ( .A1(n786), .A2(n718), .ZN(n790) );
  XOR2_X1 U631 ( .A(n792), .B(keyinput22), .Z(n786) );
  NAND4_X1 U632 ( .A1(n736), .A2(n774), .A3(n713), .A4(n793), .ZN(n792) );
  NOR2_X1 U633 ( .A1(n739), .A2(n715), .ZN(n793) );
  INV_X1 U634 ( .A(n710), .ZN(n739) );
  INV_X1 U635 ( .A(n706), .ZN(n736) );
  XOR2_X1 U636 ( .A(n794), .B(n795), .Z(G1327gat) );
  NAND2_X1 U637 ( .A1(n796), .A2(n747), .ZN(n794) );
  XOR2_X1 U638 ( .A(n797), .B(n798), .Z(G1326gat) );
  NAND2_X1 U639 ( .A1(n796), .A2(n768), .ZN(n797) );
  XNOR2_X1 U640 ( .A(G8gat), .B(n799), .ZN(G1325gat) );
  NAND2_X1 U641 ( .A1(n796), .A2(n730), .ZN(n799) );
  XNOR2_X1 U642 ( .A(n800), .B(n801), .ZN(G1324gat) );
  NAND2_X1 U643 ( .A1(n796), .A2(n733), .ZN(n800) );
  XOR2_X1 U644 ( .A(n802), .B(keyinput21), .Z(n796) );
  NAND4_X1 U645 ( .A1(n706), .A2(n762), .A3(n713), .A4(n774), .ZN(n802) );
  NAND2_X1 U646 ( .A1(n803), .A2(n804), .ZN(n774) );
  OR3_X1 U647 ( .A1(n747), .A2(n759), .A3(n730), .ZN(n804) );
  INV_X1 U648 ( .A(n758), .ZN(n730) );
  NOR2_X1 U649 ( .A1(n718), .A2(n719), .ZN(n759) );
  INV_X1 U650 ( .A(n768), .ZN(n719) );
  INV_X1 U651 ( .A(n733), .ZN(n718) );
  OR3_X1 U652 ( .A1(n768), .A2(n717), .A3(n733), .ZN(n803) );
  XOR2_X1 U653 ( .A(n805), .B(n806), .Z(n733) );
  XOR2_X1 U654 ( .A(n807), .B(n808), .Z(n806) );
  XNOR2_X1 U655 ( .A(n809), .B(n801), .ZN(n808) );
  XOR2_X1 U656 ( .A(n810), .B(n811), .Z(n805) );
  XNOR2_X1 U657 ( .A(n772), .B(n781), .ZN(n811) );
  XOR2_X1 U658 ( .A(n812), .B(n791), .Z(n810) );
  NAND2_X1 U659 ( .A1(G225gat), .A2(G233gat), .ZN(n812) );
  NOR2_X1 U660 ( .A1(n731), .A2(n758), .ZN(n717) );
  XOR2_X1 U661 ( .A(n813), .B(n814), .Z(n758) );
  XOR2_X1 U662 ( .A(n815), .B(n816), .Z(n814) );
  XNOR2_X1 U663 ( .A(n817), .B(n779), .ZN(n816) );
  XOR2_X1 U664 ( .A(n818), .B(n819), .Z(n813) );
  XNOR2_X1 U665 ( .A(n788), .B(n770), .ZN(n819) );
  XOR2_X1 U666 ( .A(n820), .B(G8gat), .Z(n818) );
  NAND2_X1 U667 ( .A1(G226gat), .A2(G233gat), .ZN(n820) );
  INV_X1 U668 ( .A(n747), .ZN(n731) );
  XOR2_X1 U669 ( .A(n821), .B(n822), .Z(n747) );
  XOR2_X1 U670 ( .A(n815), .B(n823), .Z(n822) );
  XOR2_X1 U671 ( .A(n807), .B(n795), .Z(n823) );
  INV_X1 U672 ( .A(n824), .ZN(n795) );
  XOR2_X1 U673 ( .A(n825), .B(n826), .Z(n807) );
  XNOR2_X1 U674 ( .A(n744), .B(n741), .ZN(n826) );
  XNOR2_X1 U675 ( .A(n738), .B(G162gat), .ZN(n825) );
  XOR2_X1 U676 ( .A(n827), .B(n828), .Z(n815) );
  XOR2_X1 U677 ( .A(n708), .B(n711), .Z(n828) );
  XNOR2_X1 U678 ( .A(G197gat), .B(G218gat), .ZN(n827) );
  XOR2_X1 U679 ( .A(n829), .B(n830), .Z(n821) );
  XOR2_X1 U680 ( .A(n831), .B(n832), .Z(n830) );
  NAND2_X1 U681 ( .A1(G228gat), .A2(G233gat), .ZN(n831) );
  XNOR2_X1 U682 ( .A(G106gat), .B(G78gat), .ZN(n829) );
  XOR2_X1 U683 ( .A(n833), .B(n834), .Z(n768) );
  XOR2_X1 U684 ( .A(n817), .B(n835), .Z(n834) );
  XOR2_X1 U685 ( .A(n809), .B(n798), .Z(n835) );
  INV_X1 U686 ( .A(n836), .ZN(n798) );
  XOR2_X1 U687 ( .A(n837), .B(n838), .Z(n809) );
  XOR2_X1 U688 ( .A(n756), .B(n754), .Z(n838) );
  XOR2_X1 U689 ( .A(n752), .B(G134gat), .Z(n837) );
  XOR2_X1 U690 ( .A(n839), .B(n840), .Z(n817) );
  XNOR2_X1 U691 ( .A(n728), .B(n725), .ZN(n840) );
  XOR2_X1 U692 ( .A(n723), .B(G190gat), .Z(n839) );
  XOR2_X1 U693 ( .A(n841), .B(n842), .Z(n833) );
  XOR2_X1 U694 ( .A(G99gat), .B(G71gat), .Z(n842) );
  XOR2_X1 U695 ( .A(n843), .B(G43gat), .Z(n841) );
  NAND2_X1 U696 ( .A1(G227gat), .A2(G233gat), .ZN(n843) );
  INV_X1 U697 ( .A(n742), .ZN(n713) );
  XOR2_X1 U698 ( .A(n844), .B(n845), .Z(n742) );
  XOR2_X1 U699 ( .A(n754), .B(n846), .Z(n845) );
  XNOR2_X1 U700 ( .A(n711), .B(n741), .ZN(n846) );
  XOR2_X1 U701 ( .A(keyinput14), .B(G148gat), .Z(n741) );
  XNOR2_X1 U702 ( .A(keyinput19), .B(G204gat), .ZN(n711) );
  XOR2_X1 U703 ( .A(keyinput7), .B(G120gat), .Z(n754) );
  XOR2_X1 U704 ( .A(n847), .B(n848), .Z(n844) );
  XOR2_X1 U705 ( .A(n849), .B(n725), .Z(n848) );
  XNOR2_X1 U706 ( .A(keyinput17), .B(G176gat), .ZN(n725) );
  XOR2_X1 U707 ( .A(n850), .B(n851), .Z(n847) );
  NAND2_X1 U708 ( .A1(G230gat), .A2(G233gat), .ZN(n850) );
  NOR2_X1 U709 ( .A1(n715), .A2(n710), .ZN(n762) );
  XOR2_X1 U710 ( .A(n852), .B(n853), .Z(n710) );
  XOR2_X1 U711 ( .A(n854), .B(n855), .Z(n853) );
  XOR2_X1 U712 ( .A(n849), .B(n856), .Z(n855) );
  INV_X1 U713 ( .A(n752), .ZN(n856) );
  XNOR2_X1 U714 ( .A(keyinput12), .B(G127gat), .ZN(n752) );
  XOR2_X1 U715 ( .A(n857), .B(n858), .Z(n849) );
  XNOR2_X1 U716 ( .A(n779), .B(n781), .ZN(n858) );
  XOR2_X1 U717 ( .A(keyinput6), .B(G57gat), .Z(n781) );
  XNOR2_X1 U718 ( .A(keyinput8), .B(G64gat), .ZN(n779) );
  XNOR2_X1 U719 ( .A(G71gat), .B(G78gat), .ZN(n857) );
  XOR2_X1 U720 ( .A(n859), .B(n860), .Z(n852) );
  XNOR2_X1 U721 ( .A(n708), .B(n738), .ZN(n860) );
  XOR2_X1 U722 ( .A(keyinput15), .B(G155gat), .Z(n738) );
  XNOR2_X1 U723 ( .A(keyinput20), .B(G211gat), .ZN(n708) );
  XOR2_X1 U724 ( .A(n861), .B(n862), .Z(n859) );
  INV_X1 U725 ( .A(n723), .ZN(n862) );
  XNOR2_X1 U726 ( .A(keyinput18), .B(G183gat), .ZN(n723) );
  NAND2_X1 U727 ( .A1(G231gat), .A2(G233gat), .ZN(n861) );
  INV_X1 U728 ( .A(n745), .ZN(n715) );
  XOR2_X1 U729 ( .A(n863), .B(n864), .Z(n745) );
  XOR2_X1 U730 ( .A(n756), .B(n865), .Z(n864) );
  XNOR2_X1 U731 ( .A(n728), .B(n744), .ZN(n865) );
  XNOR2_X1 U732 ( .A(keyinput13), .B(G141gat), .ZN(n744) );
  XOR2_X1 U733 ( .A(keyinput16), .B(G169gat), .Z(n728) );
  XOR2_X1 U734 ( .A(keyinput11), .B(G113gat), .Z(n756) );
  XOR2_X1 U735 ( .A(n866), .B(n867), .Z(n863) );
  XNOR2_X1 U736 ( .A(G197gat), .B(n868), .ZN(n867) );
  NAND2_X1 U737 ( .A1(G229gat), .A2(G233gat), .ZN(n868) );
  XOR2_X1 U738 ( .A(n854), .B(n869), .Z(n866) );
  XOR2_X1 U739 ( .A(n870), .B(n871), .Z(n854) );
  XOR2_X1 U740 ( .A(n836), .B(n801), .Z(n871) );
  XNOR2_X1 U741 ( .A(keyinput0), .B(G1gat), .ZN(n801) );
  XNOR2_X1 U742 ( .A(keyinput1), .B(G15gat), .ZN(n836) );
  XOR2_X1 U743 ( .A(n824), .B(G8gat), .Z(n870) );
  XNOR2_X1 U744 ( .A(keyinput2), .B(G22gat), .ZN(n824) );
  XOR2_X1 U745 ( .A(n872), .B(n873), .Z(n706) );
  XOR2_X1 U746 ( .A(n874), .B(n875), .Z(n873) );
  XOR2_X1 U747 ( .A(G162gat), .B(G134gat), .Z(n875) );
  XOR2_X1 U748 ( .A(G218gat), .B(G190gat), .Z(n874) );
  XOR2_X1 U749 ( .A(n876), .B(n851), .Z(n872) );
  XNOR2_X1 U750 ( .A(n877), .B(n878), .ZN(n851) );
  XNOR2_X1 U751 ( .A(n770), .B(n772), .ZN(n878) );
  XNOR2_X1 U752 ( .A(keyinput9), .B(G85gat), .ZN(n772) );
  XOR2_X1 U753 ( .A(keyinput10), .B(G92gat), .Z(n770) );
  XOR2_X1 U754 ( .A(G106gat), .B(n766), .Z(n877) );
  INV_X1 U755 ( .A(G99gat), .ZN(n766) );
  XOR2_X1 U756 ( .A(n879), .B(n869), .Z(n876) );
  XNOR2_X1 U757 ( .A(n880), .B(n881), .ZN(n869) );
  XOR2_X1 U758 ( .A(n785), .B(n791), .Z(n881) );
  XOR2_X1 U759 ( .A(keyinput3), .B(G29gat), .Z(n791) );
  INV_X1 U760 ( .A(n832), .ZN(n785) );
  XNOR2_X1 U761 ( .A(keyinput5), .B(G50gat), .ZN(n832) );
  XOR2_X1 U762 ( .A(n788), .B(G43gat), .Z(n880) );
  XNOR2_X1 U763 ( .A(keyinput4), .B(G36gat), .ZN(n788) );
  NAND2_X1 U764 ( .A1(G233gat), .A2(G232gat), .ZN(n879) );
endmodule

