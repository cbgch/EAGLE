//Key = 0100101110101010001010101010101101110010100001001000011010101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373;

XNOR2_X1 U757 ( .A(G107), .B(n1047), .ZN(G9) );
NAND4_X1 U758 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XNOR2_X1 U759 ( .A(KEYINPUT52), .B(n1052), .ZN(n1050) );
NOR2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR3_X1 U761 ( .A1(n1055), .A2(G953), .A3(n1056), .ZN(n1054) );
XOR2_X1 U762 ( .A(n1057), .B(KEYINPUT36), .Z(n1055) );
NAND3_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND4_X1 U764 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1059) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U766 ( .A1(n1067), .A2(n1068), .A3(KEYINPUT3), .ZN(n1065) );
NAND3_X1 U767 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1063) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1076), .ZN(n1069) );
NAND2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U772 ( .A1(n1052), .A2(KEYINPUT3), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND4_X1 U774 ( .A1(n1071), .A2(n1072), .A3(n1067), .A4(n1081), .ZN(n1058) );
NAND3_X1 U775 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1061), .A2(n1085), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U778 ( .A1(n1088), .A2(n1062), .A3(n1089), .ZN(n1082) );
INV_X1 U779 ( .A(n1066), .ZN(n1071) );
NOR3_X1 U780 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1053) );
AND4_X1 U781 ( .A1(n1090), .A2(n1067), .A3(n1091), .A4(n1092), .ZN(n1056) );
NOR4_X1 U782 ( .A1(n1089), .A2(n1079), .A3(n1093), .A4(n1094), .ZN(n1092) );
XNOR2_X1 U783 ( .A(n1095), .B(KEYINPUT18), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1096), .B(n1097), .Z(n1093) );
XOR2_X1 U785 ( .A(KEYINPUT14), .B(G469), .Z(n1097) );
NAND2_X1 U786 ( .A1(KEYINPUT45), .A2(n1098), .ZN(n1096) );
XOR2_X1 U787 ( .A(n1099), .B(n1100), .Z(n1091) );
XNOR2_X1 U788 ( .A(KEYINPUT58), .B(n1101), .ZN(n1100) );
NAND2_X1 U789 ( .A1(KEYINPUT48), .A2(n1102), .ZN(n1099) );
XOR2_X1 U790 ( .A(n1103), .B(n1104), .Z(G72) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1103) );
NAND2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U795 ( .A(KEYINPUT60), .B(n1113), .Z(n1109) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1106), .A2(n1114), .ZN(n1112) );
AND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1108), .ZN(n1116) );
XNOR2_X1 U800 ( .A(G953), .B(KEYINPUT34), .ZN(n1117) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1115) );
NOR2_X1 U802 ( .A1(KEYINPUT11), .A2(n1120), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U804 ( .A(n1123), .B(n1124), .ZN(n1122) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1121) );
NAND2_X1 U806 ( .A1(KEYINPUT4), .A2(n1127), .ZN(n1126) );
NAND2_X1 U807 ( .A1(KEYINPUT12), .A2(n1128), .ZN(n1125) );
NAND2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
OR2_X1 U810 ( .A1(n1106), .A2(G224), .ZN(n1132) );
NAND3_X1 U811 ( .A1(G953), .A2(n1133), .A3(n1134), .ZN(n1129) );
XNOR2_X1 U812 ( .A(n1131), .B(KEYINPUT55), .ZN(n1134) );
XNOR2_X1 U813 ( .A(n1135), .B(n1136), .ZN(n1131) );
NOR4_X1 U814 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
XNOR2_X1 U816 ( .A(n1143), .B(n1144), .ZN(n1142) );
INV_X1 U817 ( .A(n1145), .ZN(n1141) );
NAND2_X1 U818 ( .A1(n1106), .A2(n1146), .ZN(n1135) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1133) );
NOR2_X1 U820 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NOR2_X1 U823 ( .A1(n1147), .A2(n1153), .ZN(G63) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U825 ( .A1(G478), .A2(n1156), .A3(G902), .ZN(n1154) );
XOR2_X1 U826 ( .A(KEYINPUT63), .B(n1060), .Z(n1156) );
NOR2_X1 U827 ( .A1(n1147), .A2(n1157), .ZN(G60) );
XOR2_X1 U828 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U829 ( .A1(n1151), .A2(G475), .ZN(n1158) );
XOR2_X1 U830 ( .A(G104), .B(n1160), .Z(G6) );
NOR2_X1 U831 ( .A1(n1052), .A2(n1161), .ZN(n1160) );
NOR2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(G57) );
XOR2_X1 U833 ( .A(n1164), .B(KEYINPUT6), .Z(n1163) );
NAND2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
INV_X1 U835 ( .A(G952), .ZN(n1166) );
XNOR2_X1 U836 ( .A(G953), .B(KEYINPUT20), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1162) );
XOR2_X1 U838 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U839 ( .A(n1171), .B(n1172), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1151), .A2(G472), .ZN(n1171) );
NOR2_X1 U841 ( .A1(n1147), .A2(n1173), .ZN(G54) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U843 ( .A(n1176), .B(n1177), .ZN(n1175) );
XNOR2_X1 U844 ( .A(n1178), .B(n1179), .ZN(n1177) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR3_X1 U847 ( .A1(n1107), .A2(KEYINPUT19), .A3(G953), .ZN(n1182) );
INV_X1 U848 ( .A(G227), .ZN(n1107) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1180) );
NOR2_X1 U850 ( .A1(KEYINPUT42), .A2(n1186), .ZN(n1185) );
NAND2_X1 U851 ( .A1(n1151), .A2(G469), .ZN(n1184) );
NOR2_X1 U852 ( .A1(n1147), .A2(n1187), .ZN(G51) );
XOR2_X1 U853 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U854 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U855 ( .A1(KEYINPUT39), .A2(n1192), .ZN(n1191) );
XOR2_X1 U856 ( .A(G125), .B(n1193), .Z(n1192) );
NAND2_X1 U857 ( .A1(n1151), .A2(n1194), .ZN(n1188) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1060), .ZN(n1151) );
NOR2_X1 U859 ( .A1(n1114), .A2(n1146), .ZN(n1060) );
NAND4_X1 U860 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1146) );
AND4_X1 U861 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1068), .A2(n1204), .ZN(n1198) );
NAND2_X1 U863 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND3_X1 U864 ( .A1(n1049), .A2(n1051), .A3(n1048), .ZN(n1206) );
XNOR2_X1 U865 ( .A(KEYINPUT30), .B(n1161), .ZN(n1205) );
NAND3_X1 U866 ( .A1(n1049), .A2(n1051), .A3(n1207), .ZN(n1161) );
INV_X1 U867 ( .A(n1083), .ZN(n1049) );
NAND2_X1 U868 ( .A1(n1062), .A2(n1208), .ZN(n1083) );
NAND3_X1 U869 ( .A1(n1209), .A2(n1067), .A3(n1210), .ZN(n1196) );
NAND4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1114) );
NOR4_X1 U871 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR2_X1 U872 ( .A1(KEYINPUT23), .A2(n1219), .ZN(n1218) );
NOR2_X1 U873 ( .A1(n1220), .A2(n1075), .ZN(n1217) );
NOR2_X1 U874 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NOR3_X1 U875 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
XNOR2_X1 U876 ( .A(KEYINPUT44), .B(n1226), .ZN(n1225) );
XOR2_X1 U877 ( .A(KEYINPUT53), .B(n1072), .Z(n1223) );
NOR4_X1 U878 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1052), .ZN(n1221) );
NAND2_X1 U879 ( .A1(KEYINPUT23), .A2(n1230), .ZN(n1227) );
INV_X1 U880 ( .A(n1231), .ZN(n1216) );
NOR2_X1 U881 ( .A1(n1232), .A2(n1233), .ZN(n1213) );
NOR2_X1 U882 ( .A1(n1106), .A2(G952), .ZN(n1147) );
XNOR2_X1 U883 ( .A(G146), .B(n1231), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1207), .A2(n1068), .A3(n1234), .ZN(n1231) );
XOR2_X1 U885 ( .A(G143), .B(n1215), .Z(G45) );
AND3_X1 U886 ( .A1(n1235), .A2(n1068), .A3(n1236), .ZN(n1215) );
NOR3_X1 U887 ( .A1(n1086), .A2(n1237), .A3(n1238), .ZN(n1236) );
INV_X1 U888 ( .A(n1226), .ZN(n1086) );
XNOR2_X1 U889 ( .A(G140), .B(n1211), .ZN(G42) );
NAND4_X1 U890 ( .A1(n1072), .A2(n1235), .A3(n1207), .A4(n1239), .ZN(n1211) );
XNOR2_X1 U891 ( .A(G137), .B(n1212), .ZN(G39) );
NAND3_X1 U892 ( .A1(n1072), .A2(n1067), .A3(n1234), .ZN(n1212) );
XOR2_X1 U893 ( .A(n1240), .B(n1241), .Z(G36) );
NOR2_X1 U894 ( .A1(n1075), .A2(n1242), .ZN(n1241) );
INV_X1 U895 ( .A(n1048), .ZN(n1075) );
NOR2_X1 U896 ( .A1(KEYINPUT59), .A2(n1243), .ZN(n1240) );
INV_X1 U897 ( .A(G134), .ZN(n1243) );
XNOR2_X1 U898 ( .A(n1128), .B(n1233), .ZN(G33) );
NOR2_X1 U899 ( .A1(n1242), .A2(n1074), .ZN(n1233) );
INV_X1 U900 ( .A(n1207), .ZN(n1074) );
NAND3_X1 U901 ( .A1(n1235), .A2(n1226), .A3(n1072), .ZN(n1242) );
AND2_X1 U902 ( .A1(n1080), .A2(n1244), .ZN(n1072) );
INV_X1 U903 ( .A(G131), .ZN(n1128) );
XNOR2_X1 U904 ( .A(G128), .B(n1219), .ZN(G30) );
NAND3_X1 U905 ( .A1(n1048), .A2(n1068), .A3(n1234), .ZN(n1219) );
NOR2_X1 U906 ( .A1(n1228), .A2(n1224), .ZN(n1234) );
INV_X1 U907 ( .A(n1235), .ZN(n1224) );
NOR2_X1 U908 ( .A1(n1229), .A2(n1230), .ZN(n1235) );
INV_X1 U909 ( .A(n1245), .ZN(n1230) );
XNOR2_X1 U910 ( .A(G101), .B(n1197), .ZN(G3) );
NAND2_X1 U911 ( .A1(n1246), .A2(n1226), .ZN(n1197) );
XOR2_X1 U912 ( .A(G125), .B(n1232), .Z(G27) );
AND4_X1 U913 ( .A1(n1068), .A2(n1245), .A3(n1239), .A4(n1247), .ZN(n1232) );
AND2_X1 U914 ( .A1(n1061), .A2(n1207), .ZN(n1247) );
NAND2_X1 U915 ( .A1(n1066), .A2(n1248), .ZN(n1245) );
NAND4_X1 U916 ( .A1(G902), .A2(G953), .A3(n1249), .A4(n1108), .ZN(n1248) );
INV_X1 U917 ( .A(G900), .ZN(n1108) );
XOR2_X1 U918 ( .A(n1203), .B(n1250), .Z(G24) );
XNOR2_X1 U919 ( .A(KEYINPUT8), .B(n1251), .ZN(n1250) );
NAND4_X1 U920 ( .A1(n1210), .A2(n1062), .A3(n1252), .A4(n1253), .ZN(n1203) );
XNOR2_X1 U921 ( .A(G119), .B(n1254), .ZN(G21) );
NAND4_X1 U922 ( .A1(n1255), .A2(n1209), .A3(n1256), .A4(n1061), .ZN(n1254) );
NOR2_X1 U923 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
INV_X1 U924 ( .A(n1228), .ZN(n1209) );
NAND2_X1 U925 ( .A1(n1095), .A2(n1259), .ZN(n1228) );
XNOR2_X1 U926 ( .A(n1068), .B(KEYINPUT54), .ZN(n1255) );
XNOR2_X1 U927 ( .A(G116), .B(n1202), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1048), .A2(n1226), .A3(n1210), .ZN(n1202) );
NOR2_X1 U929 ( .A1(n1253), .A2(n1238), .ZN(n1048) );
INV_X1 U930 ( .A(n1252), .ZN(n1238) );
XNOR2_X1 U931 ( .A(G113), .B(n1201), .ZN(G15) );
NAND3_X1 U932 ( .A1(n1207), .A2(n1226), .A3(n1210), .ZN(n1201) );
AND3_X1 U933 ( .A1(n1068), .A2(n1051), .A3(n1061), .ZN(n1210) );
NOR2_X1 U934 ( .A1(n1260), .A2(n1089), .ZN(n1061) );
NAND2_X1 U935 ( .A1(n1261), .A2(n1262), .ZN(n1226) );
NAND2_X1 U936 ( .A1(n1062), .A2(n1263), .ZN(n1262) );
NOR2_X1 U937 ( .A1(n1259), .A2(n1095), .ZN(n1062) );
OR3_X1 U938 ( .A1(n1264), .A2(n1095), .A3(n1263), .ZN(n1261) );
INV_X1 U939 ( .A(KEYINPUT26), .ZN(n1263) );
NOR2_X1 U940 ( .A1(n1252), .A2(n1237), .ZN(n1207) );
INV_X1 U941 ( .A(n1253), .ZN(n1237) );
XNOR2_X1 U942 ( .A(G110), .B(n1200), .ZN(G12) );
NAND2_X1 U943 ( .A1(n1246), .A2(n1239), .ZN(n1200) );
INV_X1 U944 ( .A(n1087), .ZN(n1239) );
NAND2_X1 U945 ( .A1(n1264), .A2(n1095), .ZN(n1087) );
XNOR2_X1 U946 ( .A(n1265), .B(n1152), .ZN(n1095) );
AND2_X1 U947 ( .A1(G217), .A2(n1266), .ZN(n1152) );
NAND2_X1 U948 ( .A1(n1150), .A2(n1195), .ZN(n1265) );
XNOR2_X1 U949 ( .A(n1267), .B(n1268), .ZN(n1150) );
XOR2_X1 U950 ( .A(n1269), .B(n1270), .Z(n1267) );
NOR2_X1 U951 ( .A1(KEYINPUT62), .A2(n1271), .ZN(n1270) );
XOR2_X1 U952 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U953 ( .A(n1274), .B(n1275), .ZN(n1273) );
XOR2_X1 U954 ( .A(n1276), .B(n1277), .Z(n1272) );
NOR2_X1 U955 ( .A1(KEYINPUT2), .A2(n1278), .ZN(n1277) );
INV_X1 U956 ( .A(G119), .ZN(n1278) );
XNOR2_X1 U957 ( .A(G128), .B(KEYINPUT9), .ZN(n1276) );
NAND2_X1 U958 ( .A1(G221), .A2(n1279), .ZN(n1269) );
INV_X1 U959 ( .A(n1259), .ZN(n1264) );
XOR2_X1 U960 ( .A(n1101), .B(n1102), .Z(n1259) );
INV_X1 U961 ( .A(G472), .ZN(n1102) );
NAND2_X1 U962 ( .A1(n1280), .A2(n1195), .ZN(n1101) );
XOR2_X1 U963 ( .A(n1169), .B(n1281), .Z(n1280) );
XNOR2_X1 U964 ( .A(n1282), .B(n1283), .ZN(n1281) );
NOR2_X1 U965 ( .A1(KEYINPUT50), .A2(n1170), .ZN(n1283) );
XNOR2_X1 U966 ( .A(n1176), .B(n1284), .ZN(n1170) );
NOR2_X1 U967 ( .A1(KEYINPUT17), .A2(n1172), .ZN(n1282) );
XNOR2_X1 U968 ( .A(n1285), .B(n1286), .ZN(n1169) );
XNOR2_X1 U969 ( .A(G116), .B(n1287), .ZN(n1286) );
NAND2_X1 U970 ( .A1(G210), .A2(n1288), .ZN(n1287) );
NOR4_X1 U971 ( .A1(n1258), .A2(n1052), .A3(n1229), .A4(n1257), .ZN(n1246) );
INV_X1 U972 ( .A(n1051), .ZN(n1257) );
NAND2_X1 U973 ( .A1(n1066), .A2(n1289), .ZN(n1051) );
NAND3_X1 U974 ( .A1(n1140), .A2(n1249), .A3(G902), .ZN(n1289) );
NOR2_X1 U975 ( .A1(n1106), .A2(G898), .ZN(n1140) );
NAND3_X1 U976 ( .A1(n1249), .A2(n1106), .A3(G952), .ZN(n1066) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1249) );
INV_X1 U978 ( .A(n1208), .ZN(n1229) );
NOR2_X1 U979 ( .A1(n1088), .A2(n1089), .ZN(n1208) );
AND2_X1 U980 ( .A1(G221), .A2(n1266), .ZN(n1089) );
NAND2_X1 U981 ( .A1(G234), .A2(n1290), .ZN(n1266) );
XNOR2_X1 U982 ( .A(KEYINPUT56), .B(n1195), .ZN(n1290) );
INV_X1 U983 ( .A(n1260), .ZN(n1088) );
XOR2_X1 U984 ( .A(n1098), .B(G469), .Z(n1260) );
AND3_X1 U985 ( .A1(n1291), .A2(n1292), .A3(n1195), .ZN(n1098) );
NAND2_X1 U986 ( .A1(n1293), .A2(n1183), .ZN(n1292) );
NAND2_X1 U987 ( .A1(n1274), .A2(n1294), .ZN(n1291) );
XNOR2_X1 U988 ( .A(n1293), .B(KEYINPUT5), .ZN(n1294) );
XOR2_X1 U989 ( .A(n1179), .B(n1295), .Z(n1293) );
XNOR2_X1 U990 ( .A(G227), .B(n1296), .ZN(n1295) );
NAND3_X1 U991 ( .A1(KEYINPUT35), .A2(n1297), .A3(n1298), .ZN(n1296) );
XOR2_X1 U992 ( .A(n1299), .B(KEYINPUT25), .Z(n1298) );
OR2_X1 U993 ( .A1(n1300), .A2(n1176), .ZN(n1299) );
NAND2_X1 U994 ( .A1(n1176), .A2(n1300), .ZN(n1297) );
NAND2_X1 U995 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U996 ( .A1(n1178), .A2(n1303), .ZN(n1302) );
NAND2_X1 U997 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U998 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U999 ( .A1(n1186), .A2(n1308), .ZN(n1301) );
NAND2_X1 U1000 ( .A1(n1307), .A2(n1309), .ZN(n1308) );
NAND2_X1 U1001 ( .A1(n1123), .A2(n1304), .ZN(n1309) );
INV_X1 U1002 ( .A(KEYINPUT46), .ZN(n1304) );
INV_X1 U1003 ( .A(n1178), .ZN(n1123) );
XOR2_X1 U1004 ( .A(n1310), .B(n1311), .Z(n1178) );
NAND2_X1 U1005 ( .A1(n1312), .A2(KEYINPUT28), .ZN(n1310) );
XOR2_X1 U1006 ( .A(n1313), .B(G143), .Z(n1312) );
NAND2_X1 U1007 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XNOR2_X1 U1008 ( .A(KEYINPUT22), .B(n1316), .ZN(n1315) );
INV_X1 U1009 ( .A(G146), .ZN(n1316) );
XNOR2_X1 U1010 ( .A(KEYINPUT51), .B(KEYINPUT27), .ZN(n1314) );
INV_X1 U1011 ( .A(KEYINPUT57), .ZN(n1307) );
INV_X1 U1012 ( .A(n1306), .ZN(n1186) );
NAND2_X1 U1013 ( .A1(n1317), .A2(n1318), .ZN(n1306) );
NAND2_X1 U1014 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1015 ( .A(KEYINPUT37), .B(G101), .ZN(n1320) );
XNOR2_X1 U1016 ( .A(G104), .B(G107), .ZN(n1319) );
XOR2_X1 U1017 ( .A(n1321), .B(KEYINPUT21), .Z(n1317) );
NAND2_X1 U1018 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XNOR2_X1 U1019 ( .A(KEYINPUT37), .B(n1172), .ZN(n1323) );
INV_X1 U1020 ( .A(G101), .ZN(n1172) );
XNOR2_X1 U1021 ( .A(n1324), .B(G104), .ZN(n1322) );
INV_X1 U1022 ( .A(G107), .ZN(n1324) );
XOR2_X1 U1023 ( .A(n1325), .B(n1127), .Z(n1176) );
INV_X1 U1024 ( .A(n1268), .ZN(n1127) );
XOR2_X1 U1025 ( .A(G137), .B(KEYINPUT0), .Z(n1268) );
XNOR2_X1 U1026 ( .A(G131), .B(n1124), .ZN(n1325) );
XOR2_X1 U1027 ( .A(G140), .B(KEYINPUT61), .Z(n1179) );
INV_X1 U1028 ( .A(n1068), .ZN(n1052) );
NOR2_X1 U1029 ( .A1(n1080), .A2(n1079), .ZN(n1068) );
INV_X1 U1030 ( .A(n1244), .ZN(n1079) );
NAND2_X1 U1031 ( .A1(G214), .A2(n1326), .ZN(n1244) );
XNOR2_X1 U1032 ( .A(n1090), .B(KEYINPUT31), .ZN(n1080) );
XOR2_X1 U1033 ( .A(n1327), .B(n1194), .Z(n1090) );
AND2_X1 U1034 ( .A1(G210), .A2(n1326), .ZN(n1194) );
NAND2_X1 U1035 ( .A1(n1328), .A2(n1195), .ZN(n1326) );
INV_X1 U1036 ( .A(G237), .ZN(n1328) );
NAND2_X1 U1037 ( .A1(n1329), .A2(n1195), .ZN(n1327) );
XOR2_X1 U1038 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1039 ( .A(n1190), .B(KEYINPUT13), .Z(n1331) );
NAND4_X1 U1040 ( .A1(n1332), .A2(n1333), .A3(n1334), .A4(n1335), .ZN(n1190) );
NAND3_X1 U1041 ( .A1(n1145), .A2(n1336), .A3(n1143), .ZN(n1335) );
NAND2_X1 U1042 ( .A1(n1144), .A2(n1337), .ZN(n1336) );
NAND3_X1 U1043 ( .A1(n1338), .A2(n1144), .A3(n1339), .ZN(n1334) );
XNOR2_X1 U1044 ( .A(n1337), .B(n1145), .ZN(n1338) );
INV_X1 U1045 ( .A(n1139), .ZN(n1333) );
NOR3_X1 U1046 ( .A1(n1145), .A2(n1143), .A3(n1144), .ZN(n1139) );
INV_X1 U1047 ( .A(n1339), .ZN(n1143) );
NAND2_X1 U1048 ( .A1(n1137), .A2(n1337), .ZN(n1332) );
INV_X1 U1049 ( .A(KEYINPUT16), .ZN(n1337) );
NOR3_X1 U1050 ( .A1(n1145), .A2(n1340), .A3(n1339), .ZN(n1137) );
XNOR2_X1 U1051 ( .A(n1341), .B(n1342), .ZN(n1339) );
NOR2_X1 U1052 ( .A1(KEYINPUT15), .A2(G104), .ZN(n1342) );
XNOR2_X1 U1053 ( .A(G107), .B(G101), .ZN(n1341) );
INV_X1 U1054 ( .A(n1144), .ZN(n1340) );
XNOR2_X1 U1055 ( .A(n1343), .B(n1285), .ZN(n1144) );
XOR2_X1 U1056 ( .A(G119), .B(n1344), .Z(n1285) );
NAND2_X1 U1057 ( .A1(KEYINPUT24), .A2(n1345), .ZN(n1343) );
INV_X1 U1058 ( .A(G116), .ZN(n1345) );
XNOR2_X1 U1059 ( .A(G122), .B(n1183), .ZN(n1145) );
INV_X1 U1060 ( .A(n1274), .ZN(n1183) );
XOR2_X1 U1061 ( .A(G110), .B(KEYINPUT10), .Z(n1274) );
NAND2_X1 U1062 ( .A1(n1346), .A2(n1347), .ZN(n1330) );
OR2_X1 U1063 ( .A1(n1193), .A2(G125), .ZN(n1347) );
NAND2_X1 U1064 ( .A1(n1348), .A2(G125), .ZN(n1346) );
XOR2_X1 U1065 ( .A(KEYINPUT41), .B(n1193), .Z(n1348) );
XNOR2_X1 U1066 ( .A(n1349), .B(n1284), .ZN(n1193) );
XNOR2_X1 U1067 ( .A(n1350), .B(n1351), .ZN(n1284) );
XNOR2_X1 U1068 ( .A(G146), .B(KEYINPUT40), .ZN(n1350) );
NAND2_X1 U1069 ( .A1(G224), .A2(n1106), .ZN(n1349) );
INV_X1 U1070 ( .A(n1067), .ZN(n1258) );
NOR2_X1 U1071 ( .A1(n1252), .A2(n1253), .ZN(n1067) );
XNOR2_X1 U1072 ( .A(n1352), .B(G475), .ZN(n1253) );
NAND2_X1 U1073 ( .A1(n1159), .A2(n1195), .ZN(n1352) );
XOR2_X1 U1074 ( .A(n1275), .B(n1353), .Z(n1159) );
XNOR2_X1 U1075 ( .A(n1354), .B(n1355), .ZN(n1353) );
NOR2_X1 U1076 ( .A1(KEYINPUT29), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1077 ( .A(n1344), .B(n1357), .Z(n1356) );
XNOR2_X1 U1078 ( .A(n1251), .B(G104), .ZN(n1357) );
XOR2_X1 U1079 ( .A(G113), .B(KEYINPUT1), .Z(n1344) );
NAND2_X1 U1080 ( .A1(KEYINPUT7), .A2(n1358), .ZN(n1354) );
XOR2_X1 U1081 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1082 ( .A(G131), .B(G143), .ZN(n1360) );
NAND2_X1 U1083 ( .A1(G214), .A2(n1288), .ZN(n1359) );
NOR2_X1 U1084 ( .A1(G953), .A2(G237), .ZN(n1288) );
XNOR2_X1 U1085 ( .A(n1361), .B(n1119), .ZN(n1275) );
XOR2_X1 U1086 ( .A(G140), .B(G125), .Z(n1119) );
XNOR2_X1 U1087 ( .A(G146), .B(KEYINPUT47), .ZN(n1361) );
XNOR2_X1 U1088 ( .A(n1362), .B(G478), .ZN(n1252) );
NAND2_X1 U1089 ( .A1(n1155), .A2(n1195), .ZN(n1362) );
INV_X1 U1090 ( .A(G902), .ZN(n1195) );
XOR2_X1 U1091 ( .A(n1363), .B(n1364), .Z(n1155) );
XOR2_X1 U1092 ( .A(n1365), .B(n1366), .Z(n1364) );
NAND2_X1 U1093 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1094 ( .A1(n1369), .A2(n1251), .ZN(n1368) );
INV_X1 U1095 ( .A(G122), .ZN(n1251) );
XNOR2_X1 U1096 ( .A(G116), .B(KEYINPUT32), .ZN(n1369) );
NAND2_X1 U1097 ( .A1(G122), .A2(n1370), .ZN(n1367) );
XNOR2_X1 U1098 ( .A(G116), .B(KEYINPUT33), .ZN(n1370) );
NAND2_X1 U1099 ( .A1(G217), .A2(n1279), .ZN(n1365) );
AND2_X1 U1100 ( .A1(G234), .A2(n1106), .ZN(n1279) );
INV_X1 U1101 ( .A(G953), .ZN(n1106) );
XOR2_X1 U1102 ( .A(n1371), .B(n1372), .Z(n1363) );
NOR2_X1 U1103 ( .A1(KEYINPUT43), .A2(n1373), .ZN(n1372) );
XNOR2_X1 U1104 ( .A(n1124), .B(n1351), .ZN(n1373) );
XNOR2_X1 U1105 ( .A(n1311), .B(G143), .ZN(n1351) );
INV_X1 U1106 ( .A(G128), .ZN(n1311) );
XOR2_X1 U1107 ( .A(G134), .B(KEYINPUT49), .Z(n1124) );
XNOR2_X1 U1108 ( .A(G107), .B(KEYINPUT38), .ZN(n1371) );
endmodule


