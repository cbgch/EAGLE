//Key = 1010001001101111011000101000101110000010001000010101010100111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XNOR2_X1 U733 ( .A(G107), .B(n1011), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
XOR2_X1 U736 ( .A(n1018), .B(KEYINPUT3), .Z(n1017) );
NAND2_X1 U737 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(n1016) );
NOR2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
XOR2_X1 U740 ( .A(KEYINPUT54), .B(n1025), .Z(n1024) );
NOR4_X1 U741 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025) );
NOR4_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1029), .A4(n1032), .ZN(n1023) );
NOR3_X1 U743 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1036), .A2(n1027), .ZN(n1035) );
NOR2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR3_X1 U746 ( .A1(n1039), .A2(KEYINPUT52), .A3(n1028), .ZN(n1034) );
INV_X1 U747 ( .A(n1040), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1030) );
NOR2_X1 U749 ( .A1(n1027), .A2(n1028), .ZN(n1041) );
INV_X1 U750 ( .A(n1043), .ZN(n1027) );
NAND4_X1 U751 ( .A1(n1044), .A2(n1011), .A3(n1045), .A4(n1046), .ZN(n1014) );
NAND4_X1 U752 ( .A1(n1042), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1028), .A2(n1029), .ZN(n1049) );
INV_X1 U754 ( .A(n1050), .ZN(n1028) );
NAND3_X1 U755 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1047) );
NAND3_X1 U756 ( .A1(n1054), .A2(n1022), .A3(n1043), .ZN(n1053) );
OR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1052) );
NAND3_X1 U759 ( .A1(KEYINPUT52), .A2(n1040), .A3(n1022), .ZN(n1051) );
AND3_X1 U760 ( .A1(n1045), .A2(n1046), .A3(n1060), .ZN(n1012) );
NAND4_X1 U761 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1045) );
NOR4_X1 U762 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
XOR2_X1 U763 ( .A(KEYINPUT40), .B(n1032), .Z(n1068) );
XOR2_X1 U764 ( .A(n1069), .B(n1070), .Z(n1067) );
XOR2_X1 U765 ( .A(n1071), .B(n1072), .Z(n1066) );
XOR2_X1 U766 ( .A(KEYINPUT11), .B(n1073), .Z(n1065) );
NOR2_X1 U767 ( .A1(n1033), .A2(n1074), .ZN(n1063) );
XNOR2_X1 U768 ( .A(n1075), .B(n1076), .ZN(n1074) );
NOR2_X1 U769 ( .A1(G478), .A2(KEYINPUT21), .ZN(n1076) );
XOR2_X1 U770 ( .A(n1077), .B(n1078), .Z(n1062) );
XOR2_X1 U771 ( .A(KEYINPUT35), .B(n1079), .Z(n1078) );
NAND2_X1 U772 ( .A1(KEYINPUT6), .A2(G475), .ZN(n1077) );
XOR2_X1 U773 ( .A(n1080), .B(n1081), .Z(n1061) );
NOR2_X1 U774 ( .A1(KEYINPUT57), .A2(n1082), .ZN(n1081) );
XOR2_X1 U775 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1091), .ZN(n1085) );
INV_X1 U780 ( .A(n1087), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1092), .A2(n1090), .ZN(n1087) );
XNOR2_X1 U782 ( .A(KEYINPUT43), .B(n1093), .ZN(n1092) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U784 ( .A(KEYINPUT27), .B(n1096), .Z(n1095) );
AND2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1098), .A2(n1097), .ZN(n1094) );
NOR2_X1 U787 ( .A1(G227), .A2(n1046), .ZN(n1089) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1046), .ZN(n1083) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1019), .ZN(n1099) );
XOR2_X1 U790 ( .A(n1020), .B(KEYINPUT45), .Z(n1100) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(G69) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1046), .ZN(n1104) );
AND2_X1 U794 ( .A1(G224), .A2(G898), .ZN(n1105) );
NAND3_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1103) );
XOR2_X1 U796 ( .A(n1109), .B(KEYINPUT33), .Z(n1108) );
NAND2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
OR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
INV_X1 U799 ( .A(n1112), .ZN(n1111) );
XNOR2_X1 U800 ( .A(n1113), .B(n1114), .ZN(n1110) );
NAND2_X1 U801 ( .A1(KEYINPUT62), .A2(n1115), .ZN(n1113) );
NAND2_X1 U802 ( .A1(G953), .A2(n1116), .ZN(n1106) );
NAND2_X1 U803 ( .A1(n1046), .A2(n1117), .ZN(n1101) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U805 ( .A(KEYINPUT15), .B(n1011), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XOR2_X1 U807 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR3_X1 U808 ( .A1(n1072), .A2(n1124), .A3(n1125), .ZN(n1123) );
NOR2_X1 U809 ( .A1(KEYINPUT60), .A2(n1126), .ZN(n1125) );
NOR2_X1 U810 ( .A1(G902), .A2(n1127), .ZN(n1126) );
AND2_X1 U811 ( .A1(n1128), .A2(KEYINPUT60), .ZN(n1124) );
NAND2_X1 U812 ( .A1(KEYINPUT13), .A2(n1129), .ZN(n1122) );
NOR2_X1 U813 ( .A1(n1120), .A2(n1130), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1075), .A2(n1131), .A3(n1132), .ZN(n1130) );
AND3_X1 U815 ( .A1(n1133), .A2(G478), .A3(n1134), .ZN(n1132) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1133), .ZN(n1131) );
NOR2_X1 U817 ( .A1(n1127), .A2(n1136), .ZN(n1135) );
INV_X1 U818 ( .A(G478), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1120), .A2(n1137), .ZN(G60) );
XOR2_X1 U820 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U821 ( .A1(n1140), .A2(KEYINPUT50), .ZN(n1139) );
NAND2_X1 U822 ( .A1(n1134), .A2(G475), .ZN(n1138) );
XNOR2_X1 U823 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U824 ( .A1(n1120), .A2(n1142), .ZN(G57) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U826 ( .A(n1145), .B(n1146), .ZN(n1144) );
XNOR2_X1 U827 ( .A(n1147), .B(n1148), .ZN(n1143) );
NOR3_X1 U828 ( .A1(n1128), .A2(KEYINPUT20), .A3(n1069), .ZN(n1148) );
INV_X1 U829 ( .A(G472), .ZN(n1069) );
NAND2_X1 U830 ( .A1(KEYINPUT12), .A2(n1149), .ZN(n1147) );
NOR3_X1 U831 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(G54) );
AND2_X1 U832 ( .A1(KEYINPUT53), .A2(n1120), .ZN(n1152) );
NOR3_X1 U833 ( .A1(KEYINPUT53), .A2(n1046), .A3(n1060), .ZN(n1151) );
INV_X1 U834 ( .A(G952), .ZN(n1060) );
XOR2_X1 U835 ( .A(n1153), .B(n1154), .Z(n1150) );
XOR2_X1 U836 ( .A(n1155), .B(n1156), .Z(n1154) );
AND2_X1 U837 ( .A1(G469), .A2(n1134), .ZN(n1156) );
NOR3_X1 U838 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
AND2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR3_X1 U840 ( .A1(n1161), .A2(KEYINPUT8), .A3(n1160), .ZN(n1158) );
NAND2_X1 U841 ( .A1(n1162), .A2(KEYINPUT28), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1157) );
INV_X1 U843 ( .A(KEYINPUT8), .ZN(n1163) );
XOR2_X1 U844 ( .A(n1164), .B(n1165), .Z(n1162) );
NOR2_X1 U845 ( .A1(n1120), .A2(n1166), .ZN(G51) );
XOR2_X1 U846 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U847 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U849 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U850 ( .A(KEYINPUT63), .B(KEYINPUT58), .Z(n1174) );
INV_X1 U851 ( .A(G125), .ZN(n1171) );
XOR2_X1 U852 ( .A(n1175), .B(n1176), .Z(n1167) );
NOR2_X1 U853 ( .A1(n1080), .A2(n1128), .ZN(n1176) );
INV_X1 U854 ( .A(n1134), .ZN(n1128) );
NOR2_X1 U855 ( .A1(n1177), .A2(n1127), .ZN(n1134) );
AND4_X1 U856 ( .A1(n1118), .A2(n1019), .A3(n1011), .A4(n1020), .ZN(n1127) );
NAND3_X1 U857 ( .A1(n1043), .A2(n1178), .A3(n1037), .ZN(n1011) );
AND4_X1 U858 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1019) );
NOR4_X1 U859 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
INV_X1 U860 ( .A(n1187), .ZN(n1185) );
OR2_X1 U861 ( .A1(n1188), .A2(n1022), .ZN(n1181) );
NAND2_X1 U862 ( .A1(n1189), .A2(n1190), .ZN(n1179) );
INV_X1 U863 ( .A(n1191), .ZN(n1190) );
XOR2_X1 U864 ( .A(n1192), .B(KEYINPUT7), .Z(n1189) );
INV_X1 U865 ( .A(n1015), .ZN(n1118) );
NAND4_X1 U866 ( .A1(n1193), .A2(n1194), .A3(n1141), .A4(n1195), .ZN(n1015) );
AND4_X1 U867 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
NAND3_X1 U868 ( .A1(n1043), .A2(n1178), .A3(n1038), .ZN(n1141) );
NOR2_X1 U869 ( .A1(n1046), .A2(G952), .ZN(n1120) );
XNOR2_X1 U870 ( .A(G146), .B(n1180), .ZN(G48) );
NAND3_X1 U871 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1180) );
XOR2_X1 U872 ( .A(G143), .B(n1203), .Z(G45) );
NOR2_X1 U873 ( .A1(n1204), .A2(n1191), .ZN(n1203) );
NAND4_X1 U874 ( .A1(n1040), .A2(n1201), .A3(n1205), .A4(n1206), .ZN(n1191) );
OR2_X1 U875 ( .A1(n1038), .A2(KEYINPUT31), .ZN(n1206) );
NAND2_X1 U876 ( .A1(KEYINPUT31), .A2(n1207), .ZN(n1205) );
NAND2_X1 U877 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U878 ( .A(n1020), .B(n1210), .Z(G42) );
XOR2_X1 U879 ( .A(KEYINPUT22), .B(G140), .Z(n1210) );
NAND4_X1 U880 ( .A1(n1211), .A2(n1038), .A3(n1057), .A4(n1058), .ZN(n1020) );
XNOR2_X1 U881 ( .A(G137), .B(n1212), .ZN(G39) );
NAND2_X1 U882 ( .A1(n1213), .A2(n1059), .ZN(n1212) );
INV_X1 U883 ( .A(n1022), .ZN(n1059) );
XOR2_X1 U884 ( .A(n1188), .B(KEYINPUT9), .Z(n1213) );
NAND3_X1 U885 ( .A1(n1050), .A2(n1214), .A3(n1215), .ZN(n1188) );
INV_X1 U886 ( .A(n1026), .ZN(n1214) );
XOR2_X1 U887 ( .A(n1216), .B(n1217), .Z(G36) );
NOR2_X1 U888 ( .A1(KEYINPUT61), .A2(n1187), .ZN(n1217) );
NAND3_X1 U889 ( .A1(n1040), .A2(n1037), .A3(n1211), .ZN(n1187) );
XNOR2_X1 U890 ( .A(G134), .B(KEYINPUT59), .ZN(n1216) );
XOR2_X1 U891 ( .A(n1184), .B(n1218), .Z(G33) );
NOR2_X1 U892 ( .A1(KEYINPUT34), .A2(n1219), .ZN(n1218) );
AND3_X1 U893 ( .A1(n1038), .A2(n1040), .A3(n1211), .ZN(n1184) );
NOR3_X1 U894 ( .A1(n1026), .A2(n1204), .A3(n1022), .ZN(n1211) );
NAND2_X1 U895 ( .A1(n1056), .A2(n1055), .ZN(n1022) );
INV_X1 U896 ( .A(n1192), .ZN(n1204) );
XOR2_X1 U897 ( .A(G128), .B(n1183), .Z(G30) );
AND3_X1 U898 ( .A1(n1037), .A2(n1201), .A3(n1215), .ZN(n1183) );
AND3_X1 U899 ( .A1(n1058), .A2(n1192), .A3(n1200), .ZN(n1215) );
XOR2_X1 U900 ( .A(n1220), .B(n1193), .Z(G3) );
NAND3_X1 U901 ( .A1(n1050), .A2(n1178), .A3(n1040), .ZN(n1193) );
XOR2_X1 U902 ( .A(G125), .B(n1186), .Z(G27) );
AND3_X1 U903 ( .A1(n1221), .A2(n1057), .A3(n1202), .ZN(n1186) );
AND3_X1 U904 ( .A1(n1058), .A2(n1192), .A3(n1038), .ZN(n1202) );
NAND2_X1 U905 ( .A1(n1222), .A2(n1029), .ZN(n1192) );
NAND3_X1 U906 ( .A1(G902), .A2(n1223), .A3(n1090), .ZN(n1222) );
NOR2_X1 U907 ( .A1(G900), .A2(n1046), .ZN(n1090) );
XOR2_X1 U908 ( .A(n1194), .B(n1224), .Z(G24) );
NAND2_X1 U909 ( .A1(n1225), .A2(KEYINPUT49), .ZN(n1224) );
XNOR2_X1 U910 ( .A(G122), .B(KEYINPUT2), .ZN(n1225) );
NAND4_X1 U911 ( .A1(n1226), .A2(n1227), .A3(n1043), .A4(n1209), .ZN(n1194) );
NOR2_X1 U912 ( .A1(n1058), .A2(n1200), .ZN(n1043) );
XOR2_X1 U913 ( .A(KEYINPUT31), .B(n1228), .Z(n1226) );
XNOR2_X1 U914 ( .A(G119), .B(n1199), .ZN(G21) );
NAND4_X1 U915 ( .A1(n1200), .A2(n1227), .A3(n1050), .A4(n1058), .ZN(n1199) );
XNOR2_X1 U916 ( .A(G116), .B(n1198), .ZN(G18) );
NAND3_X1 U917 ( .A1(n1227), .A2(n1037), .A3(n1040), .ZN(n1198) );
NOR2_X1 U918 ( .A1(n1209), .A2(n1228), .ZN(n1037) );
NAND2_X1 U919 ( .A1(n1229), .A2(n1230), .ZN(G15) );
NAND2_X1 U920 ( .A1(G113), .A2(n1197), .ZN(n1230) );
XOR2_X1 U921 ( .A(n1231), .B(KEYINPUT26), .Z(n1229) );
OR2_X1 U922 ( .A1(n1197), .A2(G113), .ZN(n1231) );
NAND3_X1 U923 ( .A1(n1040), .A2(n1227), .A3(n1038), .ZN(n1197) );
AND2_X1 U924 ( .A1(n1228), .A2(n1209), .ZN(n1038) );
INV_X1 U925 ( .A(n1208), .ZN(n1228) );
AND2_X1 U926 ( .A1(n1221), .A2(n1232), .ZN(n1227) );
NOR4_X1 U927 ( .A1(n1032), .A2(n1056), .A3(n1033), .A4(n1073), .ZN(n1221) );
INV_X1 U928 ( .A(n1042), .ZN(n1033) );
NOR2_X1 U929 ( .A1(n1057), .A2(n1058), .ZN(n1040) );
XOR2_X1 U930 ( .A(n1233), .B(n1196), .Z(G12) );
NAND4_X1 U931 ( .A1(n1050), .A2(n1178), .A3(n1057), .A4(n1058), .ZN(n1196) );
XNOR2_X1 U932 ( .A(n1071), .B(n1234), .ZN(n1058) );
NOR2_X1 U933 ( .A1(KEYINPUT46), .A2(n1072), .ZN(n1234) );
NAND2_X1 U934 ( .A1(G217), .A2(n1235), .ZN(n1072) );
NAND2_X1 U935 ( .A1(n1129), .A2(n1177), .ZN(n1071) );
XNOR2_X1 U936 ( .A(n1236), .B(n1237), .ZN(n1129) );
XOR2_X1 U937 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U938 ( .A(n1240), .B(n1241), .ZN(n1239) );
NOR2_X1 U939 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1241) );
NAND2_X1 U940 ( .A1(KEYINPUT0), .A2(n1242), .ZN(n1240) );
AND2_X1 U941 ( .A1(n1243), .A2(G221), .ZN(n1238) );
XOR2_X1 U942 ( .A(n1244), .B(n1245), .Z(n1236) );
NOR2_X1 U943 ( .A1(KEYINPUT23), .A2(n1246), .ZN(n1245) );
NOR2_X1 U944 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NOR2_X1 U945 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NOR2_X1 U946 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
INV_X1 U947 ( .A(KEYINPUT55), .ZN(n1251) );
NOR2_X1 U948 ( .A1(n1253), .A2(n1254), .ZN(n1247) );
XNOR2_X1 U949 ( .A(G146), .B(KEYINPUT42), .ZN(n1254) );
NOR2_X1 U950 ( .A1(n1255), .A2(n1252), .ZN(n1253) );
XOR2_X1 U951 ( .A(G146), .B(KEYINPUT1), .Z(n1252) );
AND2_X1 U952 ( .A1(n1250), .A2(KEYINPUT55), .ZN(n1255) );
XNOR2_X1 U953 ( .A(n1256), .B(G140), .ZN(n1250) );
NAND2_X1 U954 ( .A1(KEYINPUT51), .A2(G125), .ZN(n1256) );
XOR2_X1 U955 ( .A(G119), .B(n1233), .Z(n1244) );
INV_X1 U956 ( .A(n1200), .ZN(n1057) );
XOR2_X1 U957 ( .A(n1070), .B(n1257), .Z(n1200) );
NOR2_X1 U958 ( .A1(G472), .A2(KEYINPUT44), .ZN(n1257) );
NAND2_X1 U959 ( .A1(n1258), .A2(n1177), .ZN(n1070) );
XOR2_X1 U960 ( .A(n1259), .B(n1145), .Z(n1258) );
XOR2_X1 U961 ( .A(n1260), .B(n1220), .Z(n1145) );
NAND2_X1 U962 ( .A1(G210), .A2(n1261), .ZN(n1260) );
XOR2_X1 U963 ( .A(n1262), .B(n1114), .Z(n1259) );
INV_X1 U964 ( .A(n1149), .ZN(n1114) );
NAND2_X1 U965 ( .A1(KEYINPUT30), .A2(n1146), .ZN(n1262) );
XNOR2_X1 U966 ( .A(n1169), .B(n1161), .ZN(n1146) );
AND2_X1 U967 ( .A1(n1201), .A2(n1232), .ZN(n1178) );
NAND2_X1 U968 ( .A1(n1029), .A2(n1263), .ZN(n1232) );
NAND4_X1 U969 ( .A1(G902), .A2(G953), .A3(n1223), .A4(n1116), .ZN(n1263) );
INV_X1 U970 ( .A(G898), .ZN(n1116) );
NAND3_X1 U971 ( .A1(n1223), .A2(n1046), .A3(G952), .ZN(n1029) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1223) );
NOR3_X1 U973 ( .A1(n1056), .A2(n1073), .A3(n1026), .ZN(n1201) );
NAND2_X1 U974 ( .A1(n1032), .A2(n1042), .ZN(n1026) );
NAND2_X1 U975 ( .A1(G221), .A2(n1235), .ZN(n1042) );
NAND2_X1 U976 ( .A1(G234), .A2(n1177), .ZN(n1235) );
INV_X1 U977 ( .A(n1048), .ZN(n1032) );
XOR2_X1 U978 ( .A(n1264), .B(G469), .Z(n1048) );
NAND2_X1 U979 ( .A1(n1265), .A2(n1177), .ZN(n1264) );
XOR2_X1 U980 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U981 ( .A(n1153), .B(n1097), .ZN(n1267) );
XNOR2_X1 U982 ( .A(n1161), .B(n1165), .ZN(n1097) );
XOR2_X1 U983 ( .A(n1268), .B(n1269), .Z(n1165) );
NAND2_X1 U984 ( .A1(KEYINPUT17), .A2(G128), .ZN(n1268) );
XOR2_X1 U985 ( .A(n1219), .B(n1270), .Z(n1161) );
XOR2_X1 U986 ( .A(G137), .B(G134), .Z(n1270) );
XNOR2_X1 U987 ( .A(n1271), .B(n1272), .ZN(n1153) );
XOR2_X1 U988 ( .A(G140), .B(G110), .Z(n1272) );
NAND2_X1 U989 ( .A1(G227), .A2(n1046), .ZN(n1271) );
XOR2_X1 U990 ( .A(n1164), .B(KEYINPUT29), .Z(n1266) );
NAND3_X1 U991 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1164) );
NAND2_X1 U992 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U993 ( .A1(KEYINPUT41), .A2(n1278), .ZN(n1274) );
NAND3_X1 U994 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
NAND2_X1 U995 ( .A1(n1277), .A2(G101), .ZN(n1280) );
NAND3_X1 U996 ( .A1(G107), .A2(n1282), .A3(n1220), .ZN(n1279) );
NAND2_X1 U997 ( .A1(n1283), .A2(n1284), .ZN(n1273) );
INV_X1 U998 ( .A(KEYINPUT41), .ZN(n1284) );
INV_X1 U999 ( .A(n1055), .ZN(n1073) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1285), .ZN(n1055) );
XNOR2_X1 U1001 ( .A(n1286), .B(n1080), .ZN(n1056) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1285), .ZN(n1080) );
NAND2_X1 U1003 ( .A1(n1287), .A2(n1177), .ZN(n1285) );
INV_X1 U1004 ( .A(G237), .ZN(n1287) );
XOR2_X1 U1005 ( .A(n1082), .B(KEYINPUT19), .Z(n1286) );
NAND2_X1 U1006 ( .A1(n1288), .A2(n1177), .ZN(n1082) );
INV_X1 U1007 ( .A(G902), .ZN(n1177) );
XOR2_X1 U1008 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1009 ( .A(n1291), .B(n1175), .Z(n1290) );
XOR2_X1 U1010 ( .A(n1149), .B(n1292), .Z(n1175) );
XNOR2_X1 U1011 ( .A(n1293), .B(n1294), .ZN(n1292) );
NOR2_X1 U1012 ( .A1(KEYINPUT25), .A2(n1295), .ZN(n1294) );
INV_X1 U1013 ( .A(n1115), .ZN(n1295) );
NOR2_X1 U1014 ( .A1(n1283), .A2(n1296), .ZN(n1115) );
NOR2_X1 U1015 ( .A1(n1281), .A2(n1282), .ZN(n1296) );
INV_X1 U1016 ( .A(n1276), .ZN(n1281) );
NOR2_X1 U1017 ( .A1(n1220), .A2(G107), .ZN(n1276) );
NAND2_X1 U1018 ( .A1(n1297), .A2(n1298), .ZN(n1283) );
NAND2_X1 U1019 ( .A1(n1299), .A2(G107), .ZN(n1298) );
XOR2_X1 U1020 ( .A(n1220), .B(n1282), .Z(n1299) );
INV_X1 U1021 ( .A(n1277), .ZN(n1282) );
INV_X1 U1022 ( .A(G101), .ZN(n1220) );
OR3_X1 U1023 ( .A1(n1277), .A2(G101), .A3(G107), .ZN(n1297) );
XNOR2_X1 U1024 ( .A(G104), .B(KEYINPUT18), .ZN(n1277) );
NAND2_X1 U1025 ( .A1(KEYINPUT14), .A2(n1112), .ZN(n1293) );
XOR2_X1 U1026 ( .A(n1233), .B(n1300), .Z(n1112) );
NOR2_X1 U1027 ( .A1(G122), .A2(KEYINPUT16), .ZN(n1300) );
XOR2_X1 U1028 ( .A(n1301), .B(n1302), .Z(n1149) );
XNOR2_X1 U1029 ( .A(G116), .B(G119), .ZN(n1301) );
NAND2_X1 U1030 ( .A1(KEYINPUT24), .A2(n1169), .ZN(n1291) );
NAND2_X1 U1031 ( .A1(n1303), .A2(n1304), .ZN(n1169) );
NAND2_X1 U1032 ( .A1(G128), .A2(n1305), .ZN(n1304) );
INV_X1 U1033 ( .A(n1269), .ZN(n1305) );
XOR2_X1 U1034 ( .A(n1306), .B(KEYINPUT5), .Z(n1303) );
NAND2_X1 U1035 ( .A1(n1269), .A2(n1242), .ZN(n1306) );
XOR2_X1 U1036 ( .A(n1173), .B(G125), .Z(n1289) );
NAND2_X1 U1037 ( .A1(G224), .A2(n1307), .ZN(n1173) );
XOR2_X1 U1038 ( .A(KEYINPUT32), .B(G953), .Z(n1307) );
NOR2_X1 U1039 ( .A1(n1208), .A2(n1209), .ZN(n1050) );
XOR2_X1 U1040 ( .A(n1079), .B(G475), .Z(n1209) );
NOR2_X1 U1041 ( .A1(n1140), .A2(G902), .ZN(n1079) );
AND2_X1 U1042 ( .A1(n1308), .A2(n1309), .ZN(n1140) );
NAND2_X1 U1043 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1044 ( .A(KEYINPUT47), .B(n1312), .Z(n1308) );
NOR2_X1 U1045 ( .A1(n1310), .A2(n1311), .ZN(n1312) );
XNOR2_X1 U1046 ( .A(n1313), .B(n1302), .ZN(n1311) );
XOR2_X1 U1047 ( .A(G113), .B(KEYINPUT37), .Z(n1302) );
XNOR2_X1 U1048 ( .A(G104), .B(G122), .ZN(n1313) );
XOR2_X1 U1049 ( .A(n1314), .B(n1315), .Z(n1310) );
XOR2_X1 U1050 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1051 ( .A(KEYINPUT38), .B(KEYINPUT10), .ZN(n1317) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1261), .ZN(n1316) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1261) );
XNOR2_X1 U1054 ( .A(n1318), .B(n1098), .ZN(n1314) );
XNOR2_X1 U1055 ( .A(G125), .B(G140), .ZN(n1098) );
XOR2_X1 U1056 ( .A(n1269), .B(n1319), .Z(n1318) );
NOR2_X1 U1057 ( .A1(KEYINPUT4), .A2(n1219), .ZN(n1319) );
INV_X1 U1058 ( .A(G131), .ZN(n1219) );
XNOR2_X1 U1059 ( .A(G146), .B(n1320), .ZN(n1269) );
XOR2_X1 U1060 ( .A(n1075), .B(G478), .Z(n1208) );
NOR2_X1 U1061 ( .A1(n1133), .A2(G902), .ZN(n1075) );
XOR2_X1 U1062 ( .A(n1321), .B(n1322), .Z(n1133) );
XOR2_X1 U1063 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1064 ( .A(G107), .B(n1325), .ZN(n1324) );
NOR2_X1 U1065 ( .A1(KEYINPUT48), .A2(G134), .ZN(n1325) );
XOR2_X1 U1066 ( .A(G122), .B(n1242), .Z(n1323) );
INV_X1 U1067 ( .A(G128), .ZN(n1242) );
XOR2_X1 U1068 ( .A(n1326), .B(n1320), .Z(n1321) );
XOR2_X1 U1069 ( .A(G143), .B(KEYINPUT36), .Z(n1320) );
XOR2_X1 U1070 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1071 ( .A1(G116), .A2(KEYINPUT39), .ZN(n1328) );
NAND2_X1 U1072 ( .A1(G217), .A2(n1243), .ZN(n1327) );
AND2_X1 U1073 ( .A1(G234), .A2(n1046), .ZN(n1243) );
INV_X1 U1074 ( .A(G953), .ZN(n1046) );
INV_X1 U1075 ( .A(G110), .ZN(n1233) );
endmodule


