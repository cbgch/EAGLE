//Key = 0001100001010111111001100101011111110000110110100111101111000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399;

XNOR2_X1 U767 ( .A(G107), .B(n1071), .ZN(G9) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(G75) );
NOR4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(G953), .A4(n1076), .ZN(n1073) );
NOR3_X1 U770 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1075) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1080) );
NAND4_X1 U774 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1074) );
NAND3_X1 U775 ( .A1(n1090), .A2(n1091), .A3(n1085), .ZN(n1089) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
OR2_X1 U777 ( .A1(n1091), .A2(n1085), .ZN(n1088) );
INV_X1 U778 ( .A(KEYINPUT55), .ZN(n1085) );
NAND2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND3_X1 U783 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
XNOR2_X1 U784 ( .A(KEYINPUT1), .B(n1079), .ZN(n1103) );
NAND3_X1 U785 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1100) );
NAND2_X1 U786 ( .A1(n1092), .A2(n1108), .ZN(n1096) );
NAND2_X1 U787 ( .A1(n1094), .A2(n1109), .ZN(n1087) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND3_X1 U789 ( .A1(n1112), .A2(n1099), .A3(n1106), .ZN(n1111) );
NAND2_X1 U790 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U791 ( .A1(n1104), .A2(n1115), .A3(n1116), .ZN(n1114) );
NAND2_X1 U792 ( .A1(n1105), .A2(n1117), .ZN(n1113) );
NAND3_X1 U793 ( .A1(n1092), .A2(n1118), .A3(n1119), .ZN(n1110) );
INV_X1 U794 ( .A(n1077), .ZN(n1092) );
NAND3_X1 U795 ( .A1(n1104), .A2(n1099), .A3(n1105), .ZN(n1077) );
NOR3_X1 U796 ( .A1(n1076), .A2(G953), .A3(G952), .ZN(n1072) );
AND4_X1 U797 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1076) );
NOR4_X1 U798 ( .A1(n1124), .A2(n1079), .A3(n1125), .A4(n1126), .ZN(n1123) );
XNOR2_X1 U799 ( .A(G472), .B(n1127), .ZN(n1126) );
XOR2_X1 U800 ( .A(n1128), .B(n1129), .Z(n1125) );
XNOR2_X1 U801 ( .A(G469), .B(KEYINPUT6), .ZN(n1129) );
XOR2_X1 U802 ( .A(n1130), .B(KEYINPUT56), .Z(n1124) );
NOR3_X1 U803 ( .A1(n1131), .A2(n1132), .A3(n1116), .ZN(n1122) );
NOR2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
XOR2_X1 U805 ( .A(KEYINPUT16), .B(G475), .Z(n1134) );
INV_X1 U806 ( .A(n1135), .ZN(n1133) );
XNOR2_X1 U807 ( .A(n1136), .B(n1137), .ZN(n1120) );
XNOR2_X1 U808 ( .A(n1138), .B(KEYINPUT34), .ZN(n1137) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(G72) );
NOR2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NAND2_X1 U812 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NAND2_X1 U813 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U814 ( .A1(n1149), .A2(n1142), .ZN(n1148) );
XOR2_X1 U815 ( .A(n1150), .B(KEYINPUT47), .Z(n1145) );
NAND3_X1 U816 ( .A1(n1149), .A2(n1142), .A3(n1151), .ZN(n1150) );
XNOR2_X1 U817 ( .A(n1147), .B(KEYINPUT20), .ZN(n1151) );
AND2_X1 U818 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
NAND2_X1 U819 ( .A1(n1154), .A2(n1144), .ZN(n1153) );
XOR2_X1 U820 ( .A(n1155), .B(n1156), .Z(n1152) );
XOR2_X1 U821 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U822 ( .A(n1159), .B(n1160), .ZN(n1158) );
NAND2_X1 U823 ( .A1(KEYINPUT41), .A2(n1161), .ZN(n1160) );
NAND2_X1 U824 ( .A1(KEYINPUT27), .A2(n1162), .ZN(n1159) );
XNOR2_X1 U825 ( .A(G137), .B(KEYINPUT31), .ZN(n1157) );
XOR2_X1 U826 ( .A(n1163), .B(n1164), .Z(n1155) );
XNOR2_X1 U827 ( .A(n1165), .B(n1166), .ZN(n1163) );
NOR2_X1 U828 ( .A1(KEYINPUT59), .A2(n1167), .ZN(n1166) );
XOR2_X1 U829 ( .A(n1168), .B(n1169), .Z(G69) );
XOR2_X1 U830 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U831 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U832 ( .A(KEYINPUT5), .B(n1142), .ZN(n1173) );
INV_X1 U833 ( .A(n1174), .ZN(n1172) );
NAND2_X1 U834 ( .A1(G953), .A2(n1175), .ZN(n1170) );
NAND2_X1 U835 ( .A1(G898), .A2(G224), .ZN(n1175) );
OR2_X1 U836 ( .A1(n1176), .A2(n1177), .ZN(n1168) );
NOR3_X1 U837 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(G66) );
AND2_X1 U838 ( .A1(KEYINPUT63), .A2(n1181), .ZN(n1180) );
NOR3_X1 U839 ( .A1(KEYINPUT63), .A2(G953), .A3(G952), .ZN(n1179) );
XOR2_X1 U840 ( .A(n1182), .B(n1183), .Z(n1178) );
NAND2_X1 U841 ( .A1(n1184), .A2(n1138), .ZN(n1182) );
INV_X1 U842 ( .A(n1185), .ZN(n1138) );
NOR2_X1 U843 ( .A1(n1181), .A2(n1186), .ZN(G63) );
XOR2_X1 U844 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U845 ( .A1(KEYINPUT45), .A2(n1189), .ZN(n1188) );
NAND2_X1 U846 ( .A1(n1184), .A2(G478), .ZN(n1187) );
NOR2_X1 U847 ( .A1(n1181), .A2(n1190), .ZN(G60) );
XOR2_X1 U848 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U849 ( .A1(n1184), .A2(G475), .ZN(n1191) );
XOR2_X1 U850 ( .A(n1193), .B(n1194), .Z(G6) );
XOR2_X1 U851 ( .A(KEYINPUT23), .B(G104), .Z(n1194) );
NAND2_X1 U852 ( .A1(KEYINPUT49), .A2(n1195), .ZN(n1193) );
NOR2_X1 U853 ( .A1(n1181), .A2(n1196), .ZN(G57) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U855 ( .A(n1199), .B(n1200), .Z(n1197) );
NOR2_X1 U856 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XOR2_X1 U857 ( .A(n1203), .B(KEYINPUT57), .Z(n1202) );
NAND2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U859 ( .A(KEYINPUT22), .B(n1206), .ZN(n1204) );
NOR2_X1 U860 ( .A1(n1206), .A2(n1205), .ZN(n1201) );
XOR2_X1 U861 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND2_X1 U862 ( .A1(KEYINPUT15), .A2(n1209), .ZN(n1207) );
NAND2_X1 U863 ( .A1(n1184), .A2(G472), .ZN(n1199) );
NOR2_X1 U864 ( .A1(n1181), .A2(n1210), .ZN(G54) );
XOR2_X1 U865 ( .A(n1211), .B(n1212), .Z(n1210) );
XNOR2_X1 U866 ( .A(n1208), .B(n1213), .ZN(n1212) );
NAND2_X1 U867 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
INV_X1 U869 ( .A(KEYINPUT28), .ZN(n1217) );
NAND3_X1 U870 ( .A1(n1167), .A2(n1218), .A3(KEYINPUT28), .ZN(n1214) );
XOR2_X1 U871 ( .A(n1219), .B(n1220), .Z(n1211) );
XOR2_X1 U872 ( .A(n1221), .B(n1222), .Z(n1220) );
NAND2_X1 U873 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
NAND2_X1 U874 ( .A1(n1184), .A2(G469), .ZN(n1219) );
NOR3_X1 U875 ( .A1(n1181), .A2(n1225), .A3(n1226), .ZN(G51) );
NOR2_X1 U876 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U877 ( .A(n1229), .B(n1230), .Z(n1228) );
NOR2_X1 U878 ( .A1(KEYINPUT48), .A2(n1231), .ZN(n1229) );
INV_X1 U879 ( .A(n1232), .ZN(n1231) );
NOR2_X1 U880 ( .A1(n1233), .A2(n1234), .ZN(n1225) );
XOR2_X1 U881 ( .A(n1235), .B(n1230), .Z(n1234) );
XNOR2_X1 U882 ( .A(n1236), .B(n1176), .ZN(n1230) );
NAND2_X1 U883 ( .A1(n1184), .A2(G210), .ZN(n1236) );
NOR2_X1 U884 ( .A1(n1237), .A2(n1086), .ZN(n1184) );
NOR2_X1 U885 ( .A1(n1174), .A2(n1149), .ZN(n1086) );
NAND4_X1 U886 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1149) );
AND4_X1 U887 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1241) );
NAND2_X1 U888 ( .A1(n1108), .A2(n1246), .ZN(n1240) );
NAND2_X1 U889 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XOR2_X1 U890 ( .A(n1249), .B(KEYINPUT42), .Z(n1247) );
NAND2_X1 U891 ( .A1(n1250), .A2(n1251), .ZN(n1174) );
AND4_X1 U892 ( .A1(n1252), .A2(n1253), .A3(n1071), .A4(n1254), .ZN(n1251) );
NAND3_X1 U893 ( .A1(n1094), .A2(n1117), .A3(n1255), .ZN(n1071) );
AND4_X1 U894 ( .A1(n1256), .A2(n1257), .A3(n1195), .A4(n1258), .ZN(n1250) );
NAND3_X1 U895 ( .A1(n1255), .A2(n1094), .A3(n1107), .ZN(n1195) );
NOR2_X1 U896 ( .A1(n1232), .A2(KEYINPUT48), .ZN(n1235) );
NOR2_X1 U897 ( .A1(n1259), .A2(n1260), .ZN(n1232) );
XNOR2_X1 U898 ( .A(KEYINPUT4), .B(n1261), .ZN(n1259) );
NOR2_X1 U899 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U900 ( .A(KEYINPUT40), .B(n1209), .ZN(n1263) );
XNOR2_X1 U901 ( .A(n1165), .B(KEYINPUT54), .ZN(n1262) );
INV_X1 U902 ( .A(n1227), .ZN(n1233) );
NOR2_X1 U903 ( .A1(n1142), .A2(G952), .ZN(n1181) );
XNOR2_X1 U904 ( .A(G146), .B(n1238), .ZN(G48) );
NAND3_X1 U905 ( .A1(n1107), .A2(n1108), .A3(n1264), .ZN(n1238) );
XOR2_X1 U906 ( .A(G143), .B(n1265), .Z(G45) );
NOR2_X1 U907 ( .A1(n1266), .A2(n1248), .ZN(n1265) );
NAND4_X1 U908 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1248) );
XNOR2_X1 U909 ( .A(n1108), .B(KEYINPUT26), .ZN(n1266) );
XNOR2_X1 U910 ( .A(G140), .B(n1239), .ZN(G42) );
NAND3_X1 U911 ( .A1(n1271), .A2(n1106), .A3(n1267), .ZN(n1239) );
XNOR2_X1 U912 ( .A(G137), .B(n1245), .ZN(G39) );
NAND3_X1 U913 ( .A1(n1106), .A2(n1104), .A3(n1264), .ZN(n1245) );
XOR2_X1 U914 ( .A(G134), .B(n1272), .Z(G36) );
NOR2_X1 U915 ( .A1(KEYINPUT58), .A2(n1244), .ZN(n1272) );
NAND3_X1 U916 ( .A1(n1093), .A2(n1117), .A3(n1267), .ZN(n1244) );
NAND3_X1 U917 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(G33) );
NAND2_X1 U918 ( .A1(n1276), .A2(n1243), .ZN(n1275) );
NAND2_X1 U919 ( .A1(n1277), .A2(n1278), .ZN(n1274) );
INV_X1 U920 ( .A(KEYINPUT3), .ZN(n1278) );
NAND2_X1 U921 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
INV_X1 U922 ( .A(n1276), .ZN(n1280) );
XNOR2_X1 U923 ( .A(n1243), .B(n1281), .ZN(n1279) );
NAND2_X1 U924 ( .A1(KEYINPUT3), .A2(n1282), .ZN(n1273) );
NAND2_X1 U925 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U926 ( .A1(n1243), .A2(n1281), .ZN(n1284) );
OR3_X1 U927 ( .A1(n1243), .A2(n1276), .A3(n1281), .ZN(n1283) );
INV_X1 U928 ( .A(KEYINPUT21), .ZN(n1281) );
XOR2_X1 U929 ( .A(G131), .B(KEYINPUT24), .Z(n1276) );
NAND3_X1 U930 ( .A1(n1093), .A2(n1107), .A3(n1267), .ZN(n1243) );
NOR2_X1 U931 ( .A1(n1084), .A2(n1079), .ZN(n1093) );
INV_X1 U932 ( .A(n1106), .ZN(n1079) );
NOR2_X1 U933 ( .A1(n1285), .A2(n1119), .ZN(n1106) );
XNOR2_X1 U934 ( .A(n1286), .B(n1287), .ZN(G30) );
NOR2_X1 U935 ( .A1(n1288), .A2(n1249), .ZN(n1287) );
NAND2_X1 U936 ( .A1(n1264), .A2(n1117), .ZN(n1249) );
AND3_X1 U937 ( .A1(n1083), .A2(n1289), .A3(n1267), .ZN(n1264) );
AND2_X1 U938 ( .A1(n1290), .A2(n1102), .ZN(n1267) );
INV_X1 U939 ( .A(n1108), .ZN(n1288) );
XNOR2_X1 U940 ( .A(G101), .B(n1257), .ZN(G3) );
NAND3_X1 U941 ( .A1(n1255), .A2(n1104), .A3(n1268), .ZN(n1257) );
XNOR2_X1 U942 ( .A(G125), .B(n1242), .ZN(G27) );
NAND4_X1 U943 ( .A1(n1290), .A2(n1271), .A3(n1105), .A4(n1108), .ZN(n1242) );
AND3_X1 U944 ( .A1(n1291), .A2(n1289), .A3(n1107), .ZN(n1271) );
AND2_X1 U945 ( .A1(n1292), .A2(n1099), .ZN(n1290) );
NAND2_X1 U946 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND3_X1 U947 ( .A1(G902), .A2(n1144), .A3(n1154), .ZN(n1294) );
INV_X1 U948 ( .A(n1295), .ZN(n1154) );
INV_X1 U949 ( .A(G900), .ZN(n1144) );
XNOR2_X1 U950 ( .A(G122), .B(n1256), .ZN(G24) );
NAND4_X1 U951 ( .A1(n1296), .A2(n1094), .A3(n1269), .A4(n1270), .ZN(n1256) );
AND2_X1 U952 ( .A1(n1291), .A2(n1297), .ZN(n1094) );
XNOR2_X1 U953 ( .A(G119), .B(n1254), .ZN(G21) );
NAND4_X1 U954 ( .A1(n1083), .A2(n1296), .A3(n1104), .A4(n1289), .ZN(n1254) );
XNOR2_X1 U955 ( .A(G116), .B(n1298), .ZN(G18) );
NOR2_X1 U956 ( .A1(KEYINPUT36), .A2(n1299), .ZN(n1298) );
INV_X1 U957 ( .A(n1258), .ZN(n1299) );
NAND3_X1 U958 ( .A1(n1296), .A2(n1117), .A3(n1268), .ZN(n1258) );
NAND2_X1 U959 ( .A1(n1300), .A2(n1301), .ZN(n1117) );
NAND2_X1 U960 ( .A1(n1104), .A2(n1302), .ZN(n1301) );
INV_X1 U961 ( .A(KEYINPUT62), .ZN(n1302) );
NAND3_X1 U962 ( .A1(n1303), .A2(n1269), .A3(KEYINPUT62), .ZN(n1300) );
XNOR2_X1 U963 ( .A(G113), .B(n1253), .ZN(G15) );
NAND3_X1 U964 ( .A1(n1268), .A2(n1296), .A3(n1107), .ZN(n1253) );
NOR2_X1 U965 ( .A1(n1269), .A2(n1303), .ZN(n1107) );
AND2_X1 U966 ( .A1(n1105), .A2(n1304), .ZN(n1296) );
AND2_X1 U967 ( .A1(n1115), .A2(n1305), .ZN(n1105) );
INV_X1 U968 ( .A(n1084), .ZN(n1268) );
NAND2_X1 U969 ( .A1(n1083), .A2(n1297), .ZN(n1084) );
XNOR2_X1 U970 ( .A(n1082), .B(KEYINPUT17), .ZN(n1297) );
INV_X1 U971 ( .A(n1289), .ZN(n1082) );
INV_X1 U972 ( .A(n1291), .ZN(n1083) );
XNOR2_X1 U973 ( .A(G110), .B(n1252), .ZN(G12) );
NAND4_X1 U974 ( .A1(n1255), .A2(n1104), .A3(n1291), .A4(n1289), .ZN(n1252) );
XOR2_X1 U975 ( .A(n1306), .B(n1185), .Z(n1289) );
NAND2_X1 U976 ( .A1(G217), .A2(n1307), .ZN(n1185) );
NAND2_X1 U977 ( .A1(KEYINPUT13), .A2(n1136), .ZN(n1306) );
AND2_X1 U978 ( .A1(n1183), .A2(n1237), .ZN(n1136) );
XNOR2_X1 U979 ( .A(n1308), .B(n1309), .ZN(n1183) );
NOR2_X1 U980 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
AND2_X1 U981 ( .A1(KEYINPUT14), .A2(n1312), .ZN(n1311) );
NOR2_X1 U982 ( .A1(KEYINPUT51), .A2(n1312), .ZN(n1310) );
XOR2_X1 U983 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U984 ( .A(n1315), .B(n1316), .ZN(n1314) );
XOR2_X1 U985 ( .A(G119), .B(n1317), .Z(n1316) );
NOR2_X1 U986 ( .A1(G110), .A2(KEYINPUT60), .ZN(n1317) );
INV_X1 U987 ( .A(n1165), .ZN(n1315) );
XNOR2_X1 U988 ( .A(G128), .B(n1318), .ZN(n1313) );
XNOR2_X1 U989 ( .A(n1319), .B(G140), .ZN(n1318) );
XOR2_X1 U990 ( .A(n1320), .B(G137), .Z(n1308) );
NAND2_X1 U991 ( .A1(n1321), .A2(G221), .ZN(n1320) );
XOR2_X1 U992 ( .A(n1322), .B(n1127), .Z(n1291) );
NAND2_X1 U993 ( .A1(n1323), .A2(n1237), .ZN(n1127) );
XOR2_X1 U994 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U995 ( .A(n1205), .B(n1198), .Z(n1325) );
XNOR2_X1 U996 ( .A(n1326), .B(G101), .ZN(n1198) );
NAND3_X1 U997 ( .A1(G210), .A2(n1142), .A3(n1327), .ZN(n1326) );
XNOR2_X1 U998 ( .A(n1328), .B(G113), .ZN(n1205) );
NAND2_X1 U999 ( .A1(n1329), .A2(KEYINPUT43), .ZN(n1328) );
XNOR2_X1 U1000 ( .A(G116), .B(n1330), .ZN(n1329) );
NOR2_X1 U1001 ( .A1(G119), .A2(KEYINPUT53), .ZN(n1330) );
XNOR2_X1 U1002 ( .A(n1331), .B(n1332), .ZN(n1324) );
XOR2_X1 U1003 ( .A(n1209), .B(KEYINPUT29), .Z(n1331) );
NAND2_X1 U1004 ( .A1(KEYINPUT46), .A2(n1333), .ZN(n1322) );
INV_X1 U1005 ( .A(G472), .ZN(n1333) );
NOR2_X1 U1006 ( .A1(n1269), .A2(n1270), .ZN(n1104) );
INV_X1 U1007 ( .A(n1303), .ZN(n1270) );
NOR2_X1 U1008 ( .A1(n1334), .A2(n1132), .ZN(n1303) );
NOR2_X1 U1009 ( .A1(n1135), .A2(G475), .ZN(n1132) );
AND2_X1 U1010 ( .A1(G475), .A2(n1135), .ZN(n1334) );
NAND2_X1 U1011 ( .A1(n1192), .A2(n1237), .ZN(n1135) );
XNOR2_X1 U1012 ( .A(n1335), .B(n1336), .ZN(n1192) );
XOR2_X1 U1013 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1014 ( .A(n1339), .B(G104), .ZN(n1338) );
INV_X1 U1015 ( .A(G131), .ZN(n1339) );
XNOR2_X1 U1016 ( .A(n1319), .B(G143), .ZN(n1337) );
INV_X1 U1017 ( .A(G146), .ZN(n1319) );
XNOR2_X1 U1018 ( .A(n1340), .B(n1341), .ZN(n1335) );
XOR2_X1 U1019 ( .A(n1342), .B(n1343), .Z(n1341) );
NAND2_X1 U1020 ( .A1(KEYINPUT44), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1021 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1022 ( .A1(n1347), .A2(G140), .ZN(n1346) );
XOR2_X1 U1023 ( .A(KEYINPUT32), .B(n1348), .Z(n1345) );
NOR2_X1 U1024 ( .A1(G140), .A2(n1347), .ZN(n1348) );
XNOR2_X1 U1025 ( .A(KEYINPUT33), .B(n1165), .ZN(n1347) );
NAND3_X1 U1026 ( .A1(G214), .A2(n1142), .A3(n1327), .ZN(n1342) );
XNOR2_X1 U1027 ( .A(G237), .B(KEYINPUT7), .ZN(n1327) );
NAND2_X1 U1028 ( .A1(n1130), .A2(n1121), .ZN(n1269) );
NAND2_X1 U1029 ( .A1(G478), .A2(n1349), .ZN(n1121) );
OR2_X1 U1030 ( .A1(n1349), .A2(G478), .ZN(n1130) );
OR2_X1 U1031 ( .A1(n1189), .A2(G902), .ZN(n1349) );
XOR2_X1 U1032 ( .A(n1350), .B(n1351), .Z(n1189) );
XOR2_X1 U1033 ( .A(n1352), .B(n1353), .Z(n1351) );
NAND2_X1 U1034 ( .A1(n1321), .A2(G217), .ZN(n1353) );
AND2_X1 U1035 ( .A1(G234), .A2(n1142), .ZN(n1321) );
NAND3_X1 U1036 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1352) );
NAND2_X1 U1037 ( .A1(n1162), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1038 ( .A1(KEYINPUT25), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1039 ( .A(KEYINPUT61), .B(n1359), .Z(n1358) );
NAND3_X1 U1040 ( .A1(KEYINPUT25), .A2(n1360), .A3(n1359), .ZN(n1355) );
OR2_X1 U1041 ( .A1(n1359), .A2(KEYINPUT25), .ZN(n1354) );
XOR2_X1 U1042 ( .A(G128), .B(G143), .Z(n1359) );
XNOR2_X1 U1043 ( .A(G107), .B(n1361), .ZN(n1350) );
XNOR2_X1 U1044 ( .A(G122), .B(n1362), .ZN(n1361) );
AND2_X1 U1045 ( .A1(n1304), .A2(n1102), .ZN(n1255) );
NOR2_X1 U1046 ( .A1(n1115), .A2(n1116), .ZN(n1102) );
INV_X1 U1047 ( .A(n1305), .ZN(n1116) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1237), .ZN(n1307) );
XNOR2_X1 U1050 ( .A(n1128), .B(n1363), .ZN(n1115) );
NOR2_X1 U1051 ( .A1(G469), .A2(KEYINPUT2), .ZN(n1363) );
NAND2_X1 U1052 ( .A1(n1364), .A2(n1237), .ZN(n1128) );
INV_X1 U1053 ( .A(G902), .ZN(n1237) );
XOR2_X1 U1054 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1055 ( .A(n1332), .B(n1216), .ZN(n1366) );
XOR2_X1 U1056 ( .A(n1218), .B(n1167), .Z(n1216) );
XNOR2_X1 U1057 ( .A(n1367), .B(n1286), .ZN(n1167) );
NAND2_X1 U1058 ( .A1(KEYINPUT18), .A2(n1368), .ZN(n1367) );
XNOR2_X1 U1059 ( .A(G104), .B(n1369), .ZN(n1218) );
INV_X1 U1060 ( .A(n1208), .ZN(n1332) );
XOR2_X1 U1061 ( .A(n1164), .B(n1370), .Z(n1208) );
XNOR2_X1 U1062 ( .A(n1371), .B(n1162), .ZN(n1370) );
INV_X1 U1063 ( .A(n1360), .ZN(n1162) );
XOR2_X1 U1064 ( .A(G134), .B(KEYINPUT12), .Z(n1360) );
NOR2_X1 U1065 ( .A1(G137), .A2(KEYINPUT8), .ZN(n1371) );
XOR2_X1 U1066 ( .A(G131), .B(KEYINPUT37), .Z(n1164) );
XNOR2_X1 U1067 ( .A(n1222), .B(n1372), .ZN(n1365) );
NAND2_X1 U1068 ( .A1(n1373), .A2(n1224), .ZN(n1372) );
NAND2_X1 U1069 ( .A1(G140), .A2(n1374), .ZN(n1224) );
INV_X1 U1070 ( .A(G110), .ZN(n1374) );
XOR2_X1 U1071 ( .A(n1223), .B(KEYINPUT38), .Z(n1373) );
NAND2_X1 U1072 ( .A1(G110), .A2(n1161), .ZN(n1223) );
INV_X1 U1073 ( .A(G140), .ZN(n1161) );
NOR2_X1 U1074 ( .A1(n1143), .A2(G953), .ZN(n1222) );
INV_X1 U1075 ( .A(G227), .ZN(n1143) );
AND3_X1 U1076 ( .A1(n1375), .A2(n1099), .A3(n1108), .ZN(n1304) );
NOR2_X1 U1077 ( .A1(n1118), .A2(n1119), .ZN(n1108) );
AND2_X1 U1078 ( .A1(G214), .A2(n1376), .ZN(n1119) );
OR2_X1 U1079 ( .A1(G902), .A2(G237), .ZN(n1376) );
INV_X1 U1080 ( .A(n1285), .ZN(n1118) );
NAND3_X1 U1081 ( .A1(n1377), .A2(n1378), .A3(n1379), .ZN(n1285) );
NAND2_X1 U1082 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
OR3_X1 U1083 ( .A1(n1381), .A2(n1380), .A3(G902), .ZN(n1378) );
AND2_X1 U1084 ( .A1(G237), .A2(G210), .ZN(n1380) );
XOR2_X1 U1085 ( .A(n1176), .B(n1382), .Z(n1381) );
XNOR2_X1 U1086 ( .A(n1383), .B(n1227), .ZN(n1382) );
NAND2_X1 U1087 ( .A1(G224), .A2(n1142), .ZN(n1227) );
NOR3_X1 U1088 ( .A1(n1384), .A2(KEYINPUT0), .A3(n1260), .ZN(n1383) );
AND2_X1 U1089 ( .A1(n1209), .A2(n1165), .ZN(n1260) );
NOR2_X1 U1090 ( .A1(n1209), .A2(n1385), .ZN(n1384) );
XNOR2_X1 U1091 ( .A(n1165), .B(KEYINPUT11), .ZN(n1385) );
XOR2_X1 U1092 ( .A(G125), .B(KEYINPUT50), .Z(n1165) );
XOR2_X1 U1093 ( .A(n1386), .B(n1368), .Z(n1209) );
XOR2_X1 U1094 ( .A(G143), .B(G146), .Z(n1368) );
NAND2_X1 U1095 ( .A1(KEYINPUT52), .A2(n1286), .ZN(n1386) );
INV_X1 U1096 ( .A(G128), .ZN(n1286) );
XNOR2_X1 U1097 ( .A(n1387), .B(n1388), .ZN(n1176) );
XOR2_X1 U1098 ( .A(n1389), .B(n1390), .Z(n1388) );
XNOR2_X1 U1099 ( .A(n1362), .B(G110), .ZN(n1390) );
INV_X1 U1100 ( .A(G116), .ZN(n1362) );
XOR2_X1 U1101 ( .A(KEYINPUT30), .B(KEYINPUT10), .Z(n1389) );
XOR2_X1 U1102 ( .A(n1391), .B(n1392), .Z(n1387) );
XOR2_X1 U1103 ( .A(n1393), .B(n1340), .Z(n1392) );
XOR2_X1 U1104 ( .A(G113), .B(G122), .Z(n1340) );
NOR2_X1 U1105 ( .A1(G119), .A2(KEYINPUT39), .ZN(n1393) );
NAND2_X1 U1106 ( .A1(n1394), .A2(n1395), .ZN(n1391) );
OR2_X1 U1107 ( .A1(n1369), .A2(G104), .ZN(n1395) );
NAND2_X1 U1108 ( .A1(n1396), .A2(G104), .ZN(n1394) );
XOR2_X1 U1109 ( .A(KEYINPUT19), .B(n1369), .Z(n1396) );
XNOR2_X1 U1110 ( .A(G101), .B(n1397), .ZN(n1369) );
INV_X1 U1111 ( .A(G107), .ZN(n1397) );
NAND2_X1 U1112 ( .A1(G902), .A2(G210), .ZN(n1377) );
NAND2_X1 U1113 ( .A1(G234), .A2(G237), .ZN(n1099) );
NAND2_X1 U1114 ( .A1(n1293), .A2(n1398), .ZN(n1375) );
NAND2_X1 U1115 ( .A1(n1177), .A2(G902), .ZN(n1398) );
NOR2_X1 U1116 ( .A1(n1295), .A2(G898), .ZN(n1177) );
XOR2_X1 U1117 ( .A(G953), .B(KEYINPUT35), .Z(n1295) );
NAND2_X1 U1118 ( .A1(G952), .A2(n1399), .ZN(n1293) );
XNOR2_X1 U1119 ( .A(KEYINPUT9), .B(n1142), .ZN(n1399) );
INV_X1 U1120 ( .A(G953), .ZN(n1142) );
endmodule


