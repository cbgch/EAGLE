//Key = 1100000111101001100011011101101011111000001111001111011111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;

XNOR2_X1 U667 ( .A(G107), .B(n925), .ZN(G9) );
NOR2_X1 U668 ( .A1(n926), .A2(n927), .ZN(G75) );
NOR3_X1 U669 ( .A1(n928), .A2(n929), .A3(n930), .ZN(n927) );
NAND3_X1 U670 ( .A1(n931), .A2(n932), .A3(n933), .ZN(n928) );
NAND2_X1 U671 ( .A1(n934), .A2(n935), .ZN(n933) );
NAND2_X1 U672 ( .A1(n936), .A2(n937), .ZN(n935) );
NAND3_X1 U673 ( .A1(n938), .A2(n939), .A3(n940), .ZN(n937) );
NAND2_X1 U674 ( .A1(n941), .A2(n942), .ZN(n939) );
NAND2_X1 U675 ( .A1(KEYINPUT3), .A2(n943), .ZN(n941) );
NAND4_X1 U676 ( .A1(n944), .A2(n945), .A3(n946), .A4(n947), .ZN(n938) );
NAND2_X1 U677 ( .A1(n948), .A2(n949), .ZN(n946) );
NAND2_X1 U678 ( .A1(n950), .A2(n951), .ZN(n945) );
OR2_X1 U679 ( .A1(n952), .A2(n953), .ZN(n951) );
NAND2_X1 U680 ( .A1(n943), .A2(n954), .ZN(n944) );
INV_X1 U681 ( .A(KEYINPUT3), .ZN(n954) );
NAND3_X1 U682 ( .A1(n950), .A2(n955), .A3(n948), .ZN(n936) );
NAND2_X1 U683 ( .A1(n956), .A2(n957), .ZN(n955) );
NAND2_X1 U684 ( .A1(n940), .A2(n958), .ZN(n957) );
NAND2_X1 U685 ( .A1(n959), .A2(n960), .ZN(n958) );
NAND2_X1 U686 ( .A1(n961), .A2(n962), .ZN(n960) );
NAND2_X1 U687 ( .A1(n947), .A2(n963), .ZN(n956) );
NAND2_X1 U688 ( .A1(n964), .A2(n965), .ZN(n963) );
NAND2_X1 U689 ( .A1(n966), .A2(n967), .ZN(n965) );
INV_X1 U690 ( .A(n968), .ZN(n934) );
NOR3_X1 U691 ( .A1(n969), .A2(G953), .A3(n970), .ZN(n926) );
INV_X1 U692 ( .A(n931), .ZN(n970) );
NAND2_X1 U693 ( .A1(n971), .A2(n972), .ZN(n931) );
NOR4_X1 U694 ( .A1(n962), .A2(n967), .A3(n973), .A4(n974), .ZN(n972) );
XOR2_X1 U695 ( .A(n975), .B(n976), .Z(n973) );
XOR2_X1 U696 ( .A(n977), .B(KEYINPUT11), .Z(n975) );
NOR4_X1 U697 ( .A1(n978), .A2(n979), .A3(n980), .A4(n981), .ZN(n971) );
XOR2_X1 U698 ( .A(n982), .B(n983), .Z(n981) );
XNOR2_X1 U699 ( .A(n984), .B(KEYINPUT17), .ZN(n983) );
XNOR2_X1 U700 ( .A(KEYINPUT63), .B(n929), .ZN(n969) );
INV_X1 U701 ( .A(G952), .ZN(n929) );
XOR2_X1 U702 ( .A(n985), .B(n986), .Z(G72) );
XOR2_X1 U703 ( .A(n987), .B(n988), .Z(n986) );
NOR2_X1 U704 ( .A1(n989), .A2(n990), .ZN(n988) );
XOR2_X1 U705 ( .A(n991), .B(n992), .Z(n990) );
XNOR2_X1 U706 ( .A(n993), .B(n994), .ZN(n992) );
NAND2_X1 U707 ( .A1(KEYINPUT34), .A2(n995), .ZN(n993) );
XNOR2_X1 U708 ( .A(G125), .B(n996), .ZN(n991) );
NAND2_X1 U709 ( .A1(KEYINPUT51), .A2(n997), .ZN(n996) );
NAND2_X1 U710 ( .A1(n998), .A2(n999), .ZN(n987) );
XNOR2_X1 U711 ( .A(KEYINPUT45), .B(n932), .ZN(n998) );
NAND2_X1 U712 ( .A1(G953), .A2(n1000), .ZN(n985) );
NAND2_X1 U713 ( .A1(G900), .A2(G227), .ZN(n1000) );
XOR2_X1 U714 ( .A(n1001), .B(n1002), .Z(G69) );
NOR2_X1 U715 ( .A1(n1003), .A2(n932), .ZN(n1002) );
NOR2_X1 U716 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U717 ( .A1(n1006), .A2(n1007), .ZN(n1001) );
NAND2_X1 U718 ( .A1(n1008), .A2(n932), .ZN(n1007) );
XOR2_X1 U719 ( .A(n1009), .B(n1010), .Z(n1008) );
NOR2_X1 U720 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
XOR2_X1 U721 ( .A(n1013), .B(KEYINPUT4), .Z(n1009) );
NAND2_X1 U722 ( .A1(KEYINPUT54), .A2(n1014), .ZN(n1013) );
NAND4_X1 U723 ( .A1(n1014), .A2(G898), .A3(KEYINPUT54), .A4(G953), .ZN(n1006) );
NOR2_X1 U724 ( .A1(n1015), .A2(n1016), .ZN(G66) );
XOR2_X1 U725 ( .A(n1017), .B(n1018), .Z(n1016) );
XNOR2_X1 U726 ( .A(n1019), .B(KEYINPUT43), .ZN(n1018) );
NAND3_X1 U727 ( .A1(n1020), .A2(G217), .A3(KEYINPUT1), .ZN(n1019) );
XNOR2_X1 U728 ( .A(n1021), .B(KEYINPUT15), .ZN(n1015) );
NOR2_X1 U729 ( .A1(n1021), .A2(n1022), .ZN(G63) );
XOR2_X1 U730 ( .A(n1023), .B(n1024), .Z(n1022) );
NAND2_X1 U731 ( .A1(n1020), .A2(G478), .ZN(n1023) );
NOR3_X1 U732 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(G60) );
NOR3_X1 U733 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n1027) );
AND2_X1 U734 ( .A1(n1028), .A2(n1021), .ZN(n1026) );
INV_X1 U735 ( .A(KEYINPUT5), .ZN(n1028) );
XOR2_X1 U736 ( .A(n1029), .B(n1030), .Z(n1025) );
NAND3_X1 U737 ( .A1(n1020), .A2(G475), .A3(KEYINPUT30), .ZN(n1029) );
XOR2_X1 U738 ( .A(n1031), .B(n1032), .Z(G6) );
XOR2_X1 U739 ( .A(KEYINPUT12), .B(G104), .Z(n1032) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1033), .ZN(G57) );
XOR2_X1 U741 ( .A(n1034), .B(n1035), .Z(n1033) );
XOR2_X1 U742 ( .A(n1036), .B(n1037), .Z(n1035) );
XOR2_X1 U743 ( .A(n1038), .B(n1039), .Z(n1034) );
NOR2_X1 U744 ( .A1(KEYINPUT46), .A2(n1040), .ZN(n1039) );
XNOR2_X1 U745 ( .A(n1041), .B(KEYINPUT28), .ZN(n1040) );
NAND2_X1 U746 ( .A1(n1020), .A2(G472), .ZN(n1038) );
NOR2_X1 U747 ( .A1(n1021), .A2(n1042), .ZN(G54) );
XOR2_X1 U748 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U749 ( .A1(KEYINPUT22), .A2(n1045), .ZN(n1044) );
XNOR2_X1 U750 ( .A(n1046), .B(n1047), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U752 ( .A(n1050), .B(KEYINPUT53), .Z(n1049) );
NAND2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U754 ( .A(KEYINPUT58), .B(n1053), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1053), .ZN(n1048) );
XOR2_X1 U756 ( .A(n1054), .B(G110), .Z(n1051) );
NAND2_X1 U757 ( .A1(KEYINPUT49), .A2(n997), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1020), .A2(G469), .ZN(n1043) );
NOR2_X1 U759 ( .A1(n1021), .A2(n1055), .ZN(G51) );
XOR2_X1 U760 ( .A(n1056), .B(n1057), .Z(n1055) );
NOR2_X1 U761 ( .A1(KEYINPUT14), .A2(n1058), .ZN(n1057) );
XNOR2_X1 U762 ( .A(n1059), .B(n1014), .ZN(n1058) );
XNOR2_X1 U763 ( .A(n1060), .B(n1061), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1020), .A2(n1062), .ZN(n1056) );
AND2_X1 U765 ( .A1(G902), .A2(n930), .ZN(n1020) );
OR3_X1 U766 ( .A1(n1012), .A2(n1063), .A3(n999), .ZN(n930) );
NAND4_X1 U767 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n999) );
NOR4_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U770 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1066) );
AND2_X1 U771 ( .A1(KEYINPUT56), .A2(n1077), .ZN(n1076) );
NOR4_X1 U772 ( .A1(KEYINPUT56), .A2(n1078), .A3(n1072), .A4(n1079), .ZN(n1075) );
NOR3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1074) );
XNOR2_X1 U774 ( .A(n940), .B(KEYINPUT29), .ZN(n1081) );
XOR2_X1 U775 ( .A(KEYINPUT39), .B(n1011), .Z(n1063) );
NAND4_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1011) );
NAND4_X1 U777 ( .A1(n1087), .A2(n1031), .A3(n1088), .A4(n925), .ZN(n1012) );
NAND3_X1 U778 ( .A1(n953), .A2(n950), .A3(n1089), .ZN(n925) );
NAND3_X1 U779 ( .A1(n1089), .A2(n950), .A3(n952), .ZN(n1031) );
NAND2_X1 U780 ( .A1(n943), .A2(n1089), .ZN(n1087) );
NOR2_X1 U781 ( .A1(n932), .A2(G952), .ZN(n1021) );
XNOR2_X1 U782 ( .A(n1070), .B(n1090), .ZN(G48) );
NAND2_X1 U783 ( .A1(KEYINPUT27), .A2(G146), .ZN(n1090) );
AND2_X1 U784 ( .A1(n952), .A2(n1091), .ZN(n1070) );
XOR2_X1 U785 ( .A(G143), .B(n1069), .Z(G45) );
AND4_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1069) );
NOR2_X1 U787 ( .A1(n1096), .A2(n964), .ZN(n1094) );
XNOR2_X1 U788 ( .A(G140), .B(n1064), .ZN(G42) );
NAND2_X1 U789 ( .A1(n1097), .A2(n949), .ZN(n1064) );
XOR2_X1 U790 ( .A(G137), .B(n1098), .Z(G39) );
NOR3_X1 U791 ( .A1(n1080), .A2(n1082), .A3(n1099), .ZN(n1098) );
XOR2_X1 U792 ( .A(G134), .B(n1077), .Z(G36) );
NOR2_X1 U793 ( .A1(n1078), .A2(n1082), .ZN(n1077) );
NAND3_X1 U794 ( .A1(n1093), .A2(n953), .A3(n940), .ZN(n1078) );
XNOR2_X1 U795 ( .A(G131), .B(n1065), .ZN(G33) );
NAND2_X1 U796 ( .A1(n1097), .A2(n1093), .ZN(n1065) );
AND3_X1 U797 ( .A1(n952), .A2(n1095), .A3(n940), .ZN(n1097) );
INV_X1 U798 ( .A(n1099), .ZN(n940) );
NAND2_X1 U799 ( .A1(n1100), .A2(n966), .ZN(n1099) );
INV_X1 U800 ( .A(n980), .ZN(n966) );
XOR2_X1 U801 ( .A(G128), .B(n1068), .Z(G30) );
AND2_X1 U802 ( .A1(n1091), .A2(n953), .ZN(n1068) );
NOR4_X1 U803 ( .A1(n1101), .A2(n1082), .A3(n1102), .A4(n964), .ZN(n1091) );
INV_X1 U804 ( .A(n1095), .ZN(n1082) );
NOR2_X1 U805 ( .A1(n959), .A2(n1072), .ZN(n1095) );
INV_X1 U806 ( .A(n1103), .ZN(n1072) );
XNOR2_X1 U807 ( .A(G101), .B(n1104), .ZN(G3) );
NAND4_X1 U808 ( .A1(n1105), .A2(n943), .A3(n1079), .A4(n1106), .ZN(n1104) );
AND2_X1 U809 ( .A1(n948), .A2(n1093), .ZN(n943) );
XOR2_X1 U810 ( .A(n1107), .B(KEYINPUT33), .Z(n1105) );
XNOR2_X1 U811 ( .A(n1108), .B(n1109), .ZN(G27) );
NOR2_X1 U812 ( .A1(n1073), .A2(n1110), .ZN(n1109) );
XNOR2_X1 U813 ( .A(KEYINPUT40), .B(n1103), .ZN(n1110) );
NAND2_X1 U814 ( .A1(n968), .A2(n1111), .ZN(n1103) );
NAND3_X1 U815 ( .A1(G902), .A2(n1112), .A3(n989), .ZN(n1111) );
AND2_X1 U816 ( .A1(G953), .A2(n1113), .ZN(n989) );
XOR2_X1 U817 ( .A(KEYINPUT57), .B(G900), .Z(n1113) );
NAND4_X1 U818 ( .A1(n949), .A2(n952), .A3(n947), .A4(n1114), .ZN(n1073) );
INV_X1 U819 ( .A(n942), .ZN(n947) );
XNOR2_X1 U820 ( .A(G122), .B(n1083), .ZN(G24) );
NAND4_X1 U821 ( .A1(n1092), .A2(n1115), .A3(n950), .A4(n978), .ZN(n1083) );
NOR2_X1 U822 ( .A1(n1116), .A2(n1117), .ZN(n950) );
XOR2_X1 U823 ( .A(n1084), .B(n1118), .Z(G21) );
NAND2_X1 U824 ( .A1(KEYINPUT35), .A2(G119), .ZN(n1118) );
NAND2_X1 U825 ( .A1(n1115), .A2(n1119), .ZN(n1084) );
INV_X1 U826 ( .A(n1080), .ZN(n1119) );
NAND3_X1 U827 ( .A1(n1116), .A2(n1117), .A3(n948), .ZN(n1080) );
XNOR2_X1 U828 ( .A(n1085), .B(n1120), .ZN(G18) );
NOR2_X1 U829 ( .A1(KEYINPUT13), .A2(n1121), .ZN(n1120) );
NAND3_X1 U830 ( .A1(n1093), .A2(n953), .A3(n1115), .ZN(n1085) );
NOR3_X1 U831 ( .A1(n964), .A2(n1122), .A3(n942), .ZN(n1115) );
INV_X1 U832 ( .A(n1114), .ZN(n964) );
XNOR2_X1 U833 ( .A(n1107), .B(KEYINPUT47), .ZN(n1114) );
NOR2_X1 U834 ( .A1(n1092), .A2(n1096), .ZN(n953) );
XNOR2_X1 U835 ( .A(G113), .B(n1086), .ZN(G15) );
NAND3_X1 U836 ( .A1(n952), .A2(n1093), .A3(n1123), .ZN(n1086) );
NOR3_X1 U837 ( .A1(n1107), .A2(n1122), .A3(n942), .ZN(n1123) );
NOR2_X1 U838 ( .A1(n1102), .A2(n1117), .ZN(n1093) );
INV_X1 U839 ( .A(n1101), .ZN(n1117) );
NOR2_X1 U840 ( .A1(n1124), .A2(n1125), .ZN(n952) );
INV_X1 U841 ( .A(n1092), .ZN(n1124) );
XNOR2_X1 U842 ( .A(G110), .B(n1088), .ZN(G12) );
NAND3_X1 U843 ( .A1(n949), .A2(n1089), .A3(n948), .ZN(n1088) );
NOR2_X1 U844 ( .A1(n1125), .A2(n1092), .ZN(n948) );
XNOR2_X1 U845 ( .A(n979), .B(KEYINPUT8), .ZN(n1092) );
XNOR2_X1 U846 ( .A(n1126), .B(G475), .ZN(n979) );
NAND2_X1 U847 ( .A1(n1030), .A2(n1127), .ZN(n1126) );
XNOR2_X1 U848 ( .A(n1128), .B(n1129), .ZN(n1030) );
XNOR2_X1 U849 ( .A(n1130), .B(n1131), .ZN(n1129) );
NOR2_X1 U850 ( .A1(G104), .A2(KEYINPUT18), .ZN(n1131) );
NAND2_X1 U851 ( .A1(KEYINPUT32), .A2(G113), .ZN(n1130) );
XOR2_X1 U852 ( .A(n1132), .B(G122), .Z(n1128) );
NAND2_X1 U853 ( .A1(n1133), .A2(KEYINPUT24), .ZN(n1132) );
XOR2_X1 U854 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U855 ( .A(G125), .B(n1136), .ZN(n1135) );
NAND2_X1 U856 ( .A1(KEYINPUT48), .A2(n1137), .ZN(n1136) );
XOR2_X1 U857 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U858 ( .A(n1140), .B(G131), .Z(n1139) );
NAND2_X1 U859 ( .A1(n1141), .A2(G214), .ZN(n1140) );
XNOR2_X1 U860 ( .A(G143), .B(KEYINPUT62), .ZN(n1138) );
XOR2_X1 U861 ( .A(n1096), .B(KEYINPUT20), .Z(n1125) );
INV_X1 U862 ( .A(n978), .ZN(n1096) );
XNOR2_X1 U863 ( .A(n1142), .B(n1143), .ZN(n978) );
XOR2_X1 U864 ( .A(KEYINPUT37), .B(G478), .Z(n1143) );
NAND2_X1 U865 ( .A1(n1024), .A2(n1127), .ZN(n1142) );
XNOR2_X1 U866 ( .A(n1144), .B(n1145), .ZN(n1024) );
XNOR2_X1 U867 ( .A(n1146), .B(n1147), .ZN(n1145) );
INV_X1 U868 ( .A(n1148), .ZN(n1147) );
XOR2_X1 U869 ( .A(n1149), .B(n1150), .Z(n1144) );
AND2_X1 U870 ( .A1(n1151), .A2(G217), .ZN(n1150) );
NAND2_X1 U871 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
OR2_X1 U872 ( .A1(n1154), .A2(G128), .ZN(n1153) );
XOR2_X1 U873 ( .A(n1155), .B(KEYINPUT26), .Z(n1152) );
NAND2_X1 U874 ( .A1(G128), .A2(n1154), .ZN(n1155) );
XOR2_X1 U875 ( .A(G143), .B(KEYINPUT36), .Z(n1154) );
NOR3_X1 U876 ( .A1(n959), .A2(n1122), .A3(n1107), .ZN(n1089) );
NAND2_X1 U877 ( .A1(n1100), .A2(n980), .ZN(n1107) );
XNOR2_X1 U878 ( .A(n1156), .B(n1062), .ZN(n980) );
AND2_X1 U879 ( .A1(G210), .A2(n1157), .ZN(n1062) );
NAND2_X1 U880 ( .A1(n1158), .A2(n1127), .ZN(n1156) );
XOR2_X1 U881 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U882 ( .A(n1161), .B(n1014), .Z(n1160) );
XOR2_X1 U883 ( .A(n1162), .B(n1163), .Z(n1014) );
XOR2_X1 U884 ( .A(G110), .B(n1164), .Z(n1163) );
XOR2_X1 U885 ( .A(G119), .B(G113), .Z(n1164) );
XNOR2_X1 U886 ( .A(n1148), .B(n1165), .ZN(n1162) );
XOR2_X1 U887 ( .A(G107), .B(n1166), .Z(n1148) );
XNOR2_X1 U888 ( .A(G122), .B(n1121), .ZN(n1166) );
INV_X1 U889 ( .A(G116), .ZN(n1121) );
NAND2_X1 U890 ( .A1(KEYINPUT44), .A2(n1061), .ZN(n1161) );
NOR2_X1 U891 ( .A1(n1004), .A2(G953), .ZN(n1061) );
INV_X1 U892 ( .A(G224), .ZN(n1004) );
NOR2_X1 U893 ( .A1(n1167), .A2(n1168), .ZN(n1159) );
NOR3_X1 U894 ( .A1(KEYINPUT16), .A2(n1041), .A3(n1108), .ZN(n1168) );
INV_X1 U895 ( .A(G125), .ZN(n1108) );
NOR2_X1 U896 ( .A1(n1060), .A2(n1169), .ZN(n1167) );
INV_X1 U897 ( .A(KEYINPUT16), .ZN(n1169) );
XOR2_X1 U898 ( .A(n1041), .B(G125), .Z(n1060) );
XNOR2_X1 U899 ( .A(KEYINPUT52), .B(n967), .ZN(n1100) );
AND2_X1 U900 ( .A1(G214), .A2(n1157), .ZN(n967) );
OR2_X1 U901 ( .A1(G902), .A2(G237), .ZN(n1157) );
INV_X1 U902 ( .A(n1106), .ZN(n1122) );
NAND2_X1 U903 ( .A1(n968), .A2(n1170), .ZN(n1106) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1112), .A4(n1005), .ZN(n1170) );
INV_X1 U905 ( .A(G898), .ZN(n1005) );
NAND3_X1 U906 ( .A1(n1112), .A2(n932), .A3(G952), .ZN(n968) );
NAND2_X1 U907 ( .A1(G237), .A2(G234), .ZN(n1112) );
INV_X1 U908 ( .A(n1079), .ZN(n959) );
NAND2_X1 U909 ( .A1(n1171), .A2(n1172), .ZN(n1079) );
OR2_X1 U910 ( .A1(n942), .A2(KEYINPUT7), .ZN(n1172) );
NAND2_X1 U911 ( .A1(n961), .A2(n1173), .ZN(n942) );
INV_X1 U912 ( .A(n974), .ZN(n961) );
NAND3_X1 U913 ( .A1(n974), .A2(n1173), .A3(KEYINPUT7), .ZN(n1171) );
XNOR2_X1 U914 ( .A(n962), .B(KEYINPUT59), .ZN(n1173) );
AND2_X1 U915 ( .A1(G221), .A2(n1174), .ZN(n962) );
XNOR2_X1 U916 ( .A(n1175), .B(G469), .ZN(n974) );
NAND2_X1 U917 ( .A1(n1176), .A2(n1127), .ZN(n1175) );
XOR2_X1 U918 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U919 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U920 ( .A1(KEYINPUT6), .A2(n1046), .ZN(n1180) );
XNOR2_X1 U921 ( .A(n1181), .B(n1182), .ZN(n1046) );
XNOR2_X1 U922 ( .A(n1183), .B(n1184), .ZN(n1182) );
XOR2_X1 U923 ( .A(KEYINPUT0), .B(G107), .Z(n1184) );
XOR2_X1 U924 ( .A(n995), .B(n1165), .Z(n1181) );
XOR2_X1 U925 ( .A(G101), .B(G104), .Z(n1165) );
XNOR2_X1 U926 ( .A(n1185), .B(n1186), .ZN(n995) );
NOR2_X1 U927 ( .A1(KEYINPUT38), .A2(n1187), .ZN(n1186) );
NAND2_X1 U928 ( .A1(KEYINPUT55), .A2(n1188), .ZN(n1179) );
INV_X1 U929 ( .A(n1053), .ZN(n1188) );
NAND2_X1 U930 ( .A1(G227), .A2(n932), .ZN(n1053) );
XNOR2_X1 U931 ( .A(n997), .B(G110), .ZN(n1177) );
INV_X1 U932 ( .A(G140), .ZN(n997) );
NOR2_X1 U933 ( .A1(n1101), .A2(n1116), .ZN(n949) );
INV_X1 U934 ( .A(n1102), .ZN(n1116) );
XOR2_X1 U935 ( .A(n1189), .B(n977), .Z(n1102) );
NAND3_X1 U936 ( .A1(n1190), .A2(n1191), .A3(n1127), .ZN(n977) );
NAND2_X1 U937 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
INV_X1 U938 ( .A(KEYINPUT2), .ZN(n1193) );
NAND3_X1 U939 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1192) );
OR2_X1 U940 ( .A1(n1037), .A2(n1197), .ZN(n1196) );
NAND3_X1 U941 ( .A1(n1198), .A2(n1197), .A3(n1199), .ZN(n1195) );
OR2_X1 U942 ( .A1(n1199), .A2(n1198), .ZN(n1194) );
AND2_X1 U943 ( .A1(KEYINPUT10), .A2(n1037), .ZN(n1198) );
NAND4_X1 U944 ( .A1(n1200), .A2(n1201), .A3(n1199), .A4(KEYINPUT2), .ZN(n1190) );
XOR2_X1 U945 ( .A(n1036), .B(n1202), .Z(n1199) );
INV_X1 U946 ( .A(n1041), .ZN(n1202) );
XNOR2_X1 U947 ( .A(n1187), .B(n1203), .ZN(n1041) );
XNOR2_X1 U948 ( .A(KEYINPUT23), .B(n1204), .ZN(n1203) );
INV_X1 U949 ( .A(n1185), .ZN(n1204) );
XOR2_X1 U950 ( .A(G128), .B(KEYINPUT21), .Z(n1185) );
XNOR2_X1 U951 ( .A(G146), .B(G143), .ZN(n1187) );
XNOR2_X1 U952 ( .A(n1205), .B(n1183), .ZN(n1036) );
INV_X1 U953 ( .A(n994), .ZN(n1183) );
XNOR2_X1 U954 ( .A(n1206), .B(n1146), .ZN(n994) );
XOR2_X1 U955 ( .A(G134), .B(KEYINPUT50), .Z(n1146) );
XNOR2_X1 U956 ( .A(G131), .B(G137), .ZN(n1206) );
XOR2_X1 U957 ( .A(n1207), .B(G113), .Z(n1205) );
NAND2_X1 U958 ( .A1(n1208), .A2(KEYINPUT9), .ZN(n1207) );
XNOR2_X1 U959 ( .A(G116), .B(G119), .ZN(n1208) );
NAND2_X1 U960 ( .A1(KEYINPUT41), .A2(n1209), .ZN(n1201) );
NAND2_X1 U961 ( .A1(KEYINPUT10), .A2(n1037), .ZN(n1209) );
NAND2_X1 U962 ( .A1(n1037), .A2(n1197), .ZN(n1200) );
INV_X1 U963 ( .A(KEYINPUT41), .ZN(n1197) );
XNOR2_X1 U964 ( .A(n1210), .B(G101), .ZN(n1037) );
NAND2_X1 U965 ( .A1(n1141), .A2(G210), .ZN(n1210) );
NOR2_X1 U966 ( .A1(G953), .A2(G237), .ZN(n1141) );
NAND2_X1 U967 ( .A1(KEYINPUT42), .A2(n976), .ZN(n1189) );
XOR2_X1 U968 ( .A(G472), .B(KEYINPUT25), .Z(n976) );
XNOR2_X1 U969 ( .A(n982), .B(n1211), .ZN(n1101) );
NOR2_X1 U970 ( .A1(n984), .A2(KEYINPUT19), .ZN(n1211) );
AND2_X1 U971 ( .A1(G217), .A2(n1174), .ZN(n984) );
NAND2_X1 U972 ( .A1(G234), .A2(n1127), .ZN(n1174) );
NAND2_X1 U973 ( .A1(n1017), .A2(n1127), .ZN(n982) );
INV_X1 U974 ( .A(G902), .ZN(n1127) );
XOR2_X1 U975 ( .A(n1212), .B(n1213), .Z(n1017) );
XOR2_X1 U976 ( .A(n1134), .B(n1214), .Z(n1213) );
XOR2_X1 U977 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U978 ( .A1(G125), .A2(KEYINPUT31), .ZN(n1216) );
NAND2_X1 U979 ( .A1(n1151), .A2(G221), .ZN(n1215) );
AND2_X1 U980 ( .A1(G234), .A2(n932), .ZN(n1151) );
INV_X1 U981 ( .A(G953), .ZN(n932) );
XNOR2_X1 U982 ( .A(G146), .B(G140), .ZN(n1134) );
XOR2_X1 U983 ( .A(n1217), .B(n1218), .Z(n1212) );
XOR2_X1 U984 ( .A(G137), .B(G128), .Z(n1218) );
XOR2_X1 U985 ( .A(n1219), .B(G110), .Z(n1217) );
NAND2_X1 U986 ( .A1(n1220), .A2(KEYINPUT60), .ZN(n1219) );
XNOR2_X1 U987 ( .A(G119), .B(KEYINPUT61), .ZN(n1220) );
endmodule


