//Key = 0011001110011011010000101111001000011010110010110001010110100110


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204;

XOR2_X2 U1239 ( .A(RESTART), .B(KEYINPUT35), .Z(n1942) );
INV_X2 U1240 ( .A(n1814), .ZN(n1797) );
XOR2_X1 U1241 ( .A(U280), .B(KEYINPUT21), .Z(n1802) );
INV_X1 U1242 ( .A(n1802), .ZN(n1657) );
INV_X1 U1243 ( .A(n1802), .ZN(n1658) );
INV_X1 U1244 ( .A(n1659), .ZN(U375) );
NAND2_X1 U1245 ( .A1(n1660), .A2(n1661), .ZN(U344) );
NAND2_X1 U1246 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1662), .ZN(n1661) );
NAND2_X1 U1247 ( .A1(n1663), .A2(DATA_IN_7_), .ZN(n1660) );
NAND2_X1 U1248 ( .A1(n1664), .A2(n1665), .ZN(U343) );
NAND2_X1 U1249 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1662), .ZN(n1665) );
NAND2_X1 U1250 ( .A1(n1663), .A2(DATA_IN_6_), .ZN(n1664) );
NAND2_X1 U1251 ( .A1(n1666), .A2(n1667), .ZN(U342) );
NAND2_X1 U1252 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1662), .ZN(n1667) );
NAND2_X1 U1253 ( .A1(n1663), .A2(DATA_IN_5_), .ZN(n1666) );
NAND2_X1 U1254 ( .A1(n1668), .A2(n1669), .ZN(U341) );
NAND2_X1 U1255 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1662), .ZN(n1669) );
XOR2_X1 U1256 ( .A(KEYINPUT24), .B(n1670), .Z(n1668) );
NOR2_X1 U1257 ( .A1(n1671), .A2(n1662), .ZN(n1670) );
NAND2_X1 U1258 ( .A1(n1672), .A2(n1673), .ZN(U340) );
NAND2_X1 U1259 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1662), .ZN(n1673) );
NAND2_X1 U1260 ( .A1(n1663), .A2(DATA_IN_3_), .ZN(n1672) );
NAND2_X1 U1261 ( .A1(n1674), .A2(n1675), .ZN(U339) );
NAND2_X1 U1262 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1662), .ZN(n1675) );
NAND2_X1 U1263 ( .A1(n1663), .A2(DATA_IN_2_), .ZN(n1674) );
NAND2_X1 U1264 ( .A1(n1676), .A2(n1677), .ZN(U338) );
NAND2_X1 U1265 ( .A1(n1678), .A2(n1662), .ZN(n1677) );
XOR2_X1 U1266 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT37), .Z(n1678) );
NAND2_X1 U1267 ( .A1(n1679), .A2(n1663), .ZN(n1676) );
XOR2_X1 U1268 ( .A(KEYINPUT20), .B(DATA_IN_1_), .Z(n1679) );
NAND2_X1 U1269 ( .A1(n1680), .A2(n1681), .ZN(U337) );
NAND2_X1 U1270 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1662), .ZN(n1681) );
NAND2_X1 U1271 ( .A1(n1682), .A2(n1663), .ZN(n1680) );
INV_X1 U1272 ( .A(n1662), .ZN(n1663) );
NAND2_X1 U1273 ( .A1(n1659), .A2(n1683), .ZN(n1662) );
NAND2_X1 U1274 ( .A1(n1684), .A2(n1685), .ZN(n1683) );
XOR2_X1 U1275 ( .A(n1686), .B(KEYINPUT56), .Z(n1682) );
NAND2_X1 U1276 ( .A1(n1687), .A2(n1688), .ZN(U336) );
NAND2_X1 U1277 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1689), .ZN(n1688) );
NAND2_X1 U1278 ( .A1(n1690), .A2(DATA_IN_7_), .ZN(n1687) );
NAND2_X1 U1279 ( .A1(n1691), .A2(n1692), .ZN(U335) );
NAND2_X1 U1280 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1689), .ZN(n1692) );
NAND2_X1 U1281 ( .A1(n1690), .A2(DATA_IN_6_), .ZN(n1691) );
NAND2_X1 U1282 ( .A1(n1693), .A2(n1694), .ZN(U334) );
NAND2_X1 U1283 ( .A1(DATA_IN_5_), .A2(n1695), .ZN(n1694) );
XOR2_X1 U1284 ( .A(KEYINPUT4), .B(n1690), .Z(n1695) );
NAND2_X1 U1285 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1689), .ZN(n1693) );
NAND2_X1 U1286 ( .A1(n1696), .A2(n1697), .ZN(U333) );
NAND2_X1 U1287 ( .A1(n1690), .A2(DATA_IN_4_), .ZN(n1697) );
XOR2_X1 U1288 ( .A(n1698), .B(KEYINPUT60), .Z(n1696) );
NAND2_X1 U1289 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1689), .ZN(n1698) );
NAND2_X1 U1290 ( .A1(n1699), .A2(n1700), .ZN(U332) );
NAND2_X1 U1291 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1689), .ZN(n1700) );
NAND2_X1 U1292 ( .A1(n1690), .A2(DATA_IN_3_), .ZN(n1699) );
NAND2_X1 U1293 ( .A1(n1701), .A2(n1702), .ZN(U331) );
NAND2_X1 U1294 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1689), .ZN(n1702) );
NAND2_X1 U1295 ( .A1(n1690), .A2(DATA_IN_2_), .ZN(n1701) );
NAND2_X1 U1296 ( .A1(n1703), .A2(n1704), .ZN(U330) );
NAND2_X1 U1297 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1689), .ZN(n1704) );
NAND2_X1 U1298 ( .A1(n1690), .A2(DATA_IN_1_), .ZN(n1703) );
NAND2_X1 U1299 ( .A1(n1705), .A2(n1706), .ZN(U329) );
NAND2_X1 U1300 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1689), .ZN(n1706) );
NAND2_X1 U1301 ( .A1(n1690), .A2(DATA_IN_0_), .ZN(n1705) );
INV_X1 U1302 ( .A(n1689), .ZN(n1690) );
NAND2_X1 U1303 ( .A1(n1659), .A2(n1707), .ZN(n1689) );
NAND2_X1 U1304 ( .A1(n1708), .A2(n1685), .ZN(n1707) );
NAND2_X1 U1305 ( .A1(n1709), .A2(n1710), .ZN(n1708) );
NAND2_X1 U1306 ( .A1(n1711), .A2(n1712), .ZN(n1710) );
NAND3_X1 U1307 ( .A1(n1713), .A2(n1714), .A3(n1715), .ZN(n1712) );
NAND2_X1 U1308 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1716), .ZN(n1715) );
NAND3_X1 U1309 ( .A1(n1717), .A2(n1718), .A3(n1719), .ZN(n1714) );
NAND2_X1 U1310 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1720), .ZN(n1719) );
NAND3_X1 U1311 ( .A1(n1721), .A2(n1722), .A3(n1723), .ZN(n1718) );
XOR2_X1 U1312 ( .A(KEYINPUT15), .B(n1724), .Z(n1723) );
NOR2_X1 U1313 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1720), .ZN(n1724) );
NAND3_X1 U1314 ( .A1(n1725), .A2(n1726), .A3(n1727), .ZN(n1722) );
NAND2_X1 U1315 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1671), .ZN(n1727) );
NAND3_X1 U1316 ( .A1(n1728), .A2(n1729), .A3(n1730), .ZN(n1726) );
NAND2_X1 U1317 ( .A1(DATA_IN_2_), .A2(n1731), .ZN(n1730) );
NAND3_X1 U1318 ( .A1(n1732), .A2(n1733), .A3(n1734), .ZN(n1729) );
OR2_X1 U1319 ( .A1(n1731), .A2(DATA_IN_2_), .ZN(n1734) );
NAND3_X1 U1320 ( .A1(n1735), .A2(n1686), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1733) );
NAND2_X1 U1321 ( .A1(n1736), .A2(n1737), .ZN(n1735) );
XOR2_X1 U1322 ( .A(KEYINPUT50), .B(DATA_IN_1_), .Z(n1736) );
NAND2_X1 U1323 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1738), .ZN(n1732) );
NAND2_X1 U1324 ( .A1(DATA_IN_3_), .A2(n1739), .ZN(n1728) );
XOR2_X1 U1325 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT12), .Z(n1739) );
NAND2_X1 U1326 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1740), .ZN(n1725) );
NAND2_X1 U1327 ( .A1(n1741), .A2(DATA_IN_4_), .ZN(n1721) );
XNOR2_X1 U1328 ( .A(RMIN_REG_4__SCAN_IN), .B(KEYINPUT39), .ZN(n1741) );
NAND2_X1 U1329 ( .A1(n1742), .A2(n1743), .ZN(n1717) );
XOR2_X1 U1330 ( .A(n1744), .B(KEYINPUT22), .Z(n1742) );
NAND2_X1 U1331 ( .A1(DATA_IN_6_), .A2(n1744), .ZN(n1713) );
OR2_X1 U1332 ( .A1(n1716), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1711) );
XOR2_X1 U1333 ( .A(KEYINPUT9), .B(n1684), .Z(n1709) );
AND2_X1 U1334 ( .A1(n1745), .A2(n1746), .ZN(n1684) );
NAND3_X1 U1335 ( .A1(n1747), .A2(n1748), .A3(n1749), .ZN(n1746) );
OR2_X1 U1336 ( .A1(n1716), .A2(RMAX_REG_7__SCAN_IN), .ZN(n1749) );
NAND3_X1 U1337 ( .A1(n1750), .A2(n1751), .A3(n1752), .ZN(n1748) );
NAND2_X1 U1338 ( .A1(DATA_IN_6_), .A2(n1753), .ZN(n1752) );
NAND3_X1 U1339 ( .A1(n1754), .A2(n1755), .A3(n1756), .ZN(n1751) );
NAND2_X1 U1340 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1720), .ZN(n1756) );
NAND3_X1 U1341 ( .A1(n1757), .A2(n1758), .A3(n1759), .ZN(n1755) );
OR2_X1 U1342 ( .A1(n1671), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1759) );
NAND3_X1 U1343 ( .A1(n1760), .A2(n1761), .A3(n1762), .ZN(n1758) );
XOR2_X1 U1344 ( .A(KEYINPUT27), .B(n1763), .Z(n1762) );
NOR2_X1 U1345 ( .A1(DATA_IN_2_), .A2(n1764), .ZN(n1763) );
NAND3_X1 U1346 ( .A1(n1765), .A2(n1766), .A3(n1767), .ZN(n1761) );
XOR2_X1 U1347 ( .A(n1768), .B(KEYINPUT18), .Z(n1767) );
NAND2_X1 U1348 ( .A1(DATA_IN_2_), .A2(n1769), .ZN(n1768) );
XOR2_X1 U1349 ( .A(RMAX_REG_2__SCAN_IN), .B(KEYINPUT47), .Z(n1769) );
NAND3_X1 U1350 ( .A1(n1770), .A2(n1771), .A3(DATA_IN_0_), .ZN(n1766) );
INV_X1 U1351 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1771) );
NAND2_X1 U1352 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1738), .ZN(n1770) );
INV_X1 U1353 ( .A(DATA_IN_1_), .ZN(n1738) );
NAND2_X1 U1354 ( .A1(DATA_IN_1_), .A2(n1772), .ZN(n1765) );
NAND2_X1 U1355 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1740), .ZN(n1760) );
OR2_X1 U1356 ( .A1(n1740), .A2(RMAX_REG_3__SCAN_IN), .ZN(n1757) );
INV_X1 U1357 ( .A(DATA_IN_3_), .ZN(n1740) );
NAND2_X1 U1358 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1671), .ZN(n1754) );
OR2_X1 U1359 ( .A1(n1720), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1750) );
INV_X1 U1360 ( .A(DATA_IN_5_), .ZN(n1720) );
NAND2_X1 U1361 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1743), .ZN(n1747) );
INV_X1 U1362 ( .A(DATA_IN_6_), .ZN(n1743) );
NAND2_X1 U1363 ( .A1(n1773), .A2(n1716), .ZN(n1745) );
INV_X1 U1364 ( .A(DATA_IN_7_), .ZN(n1716) );
XNOR2_X1 U1365 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT53), .ZN(n1773) );
NAND2_X1 U1366 ( .A1(n1774), .A2(n1775), .ZN(U328) );
NAND2_X1 U1367 ( .A1(DATA_IN_7_), .A2(n1776), .ZN(n1775) );
NAND2_X1 U1368 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1777), .ZN(n1774) );
NAND2_X1 U1369 ( .A1(n1778), .A2(n1779), .ZN(U327) );
NAND2_X1 U1370 ( .A1(DATA_IN_6_), .A2(n1776), .ZN(n1779) );
NAND2_X1 U1371 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1777), .ZN(n1778) );
NAND2_X1 U1372 ( .A1(n1780), .A2(n1781), .ZN(U326) );
NAND2_X1 U1373 ( .A1(DATA_IN_5_), .A2(n1776), .ZN(n1781) );
NAND2_X1 U1374 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1777), .ZN(n1780) );
NAND2_X1 U1375 ( .A1(n1782), .A2(n1783), .ZN(U325) );
NAND2_X1 U1376 ( .A1(DATA_IN_4_), .A2(n1776), .ZN(n1783) );
NAND2_X1 U1377 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1777), .ZN(n1782) );
NAND2_X1 U1378 ( .A1(n1784), .A2(n1785), .ZN(U324) );
NAND2_X1 U1379 ( .A1(n1786), .A2(n1776), .ZN(n1785) );
XOR2_X1 U1380 ( .A(KEYINPUT5), .B(DATA_IN_3_), .Z(n1786) );
NAND2_X1 U1381 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1777), .ZN(n1784) );
NAND2_X1 U1382 ( .A1(n1787), .A2(n1788), .ZN(U323) );
NAND2_X1 U1383 ( .A1(DATA_IN_2_), .A2(n1776), .ZN(n1788) );
NAND2_X1 U1384 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1777), .ZN(n1787) );
NAND2_X1 U1385 ( .A1(n1789), .A2(n1790), .ZN(U322) );
NAND2_X1 U1386 ( .A1(DATA_IN_1_), .A2(n1776), .ZN(n1790) );
NAND2_X1 U1387 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1777), .ZN(n1789) );
NAND2_X1 U1388 ( .A1(n1791), .A2(n1792), .ZN(U321) );
NAND2_X1 U1389 ( .A1(DATA_IN_0_), .A2(n1776), .ZN(n1792) );
NAND2_X1 U1390 ( .A1(n1793), .A2(n1794), .ZN(n1776) );
NAND3_X1 U1391 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1795), .A3(n1796), .ZN(n1794) );
INV_X1 U1392 ( .A(KEYINPUT31), .ZN(n1796) );
NAND3_X1 U1393 ( .A1(n1797), .A2(n1798), .A3(KEYINPUT31), .ZN(n1793) );
NAND2_X1 U1394 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1777), .ZN(n1791) );
NAND2_X1 U1395 ( .A1(n1659), .A2(n1795), .ZN(n1777) );
NAND2_X1 U1396 ( .A1(n1685), .A2(n1798), .ZN(n1795) );
NAND2_X1 U1397 ( .A1(n1685), .A2(n1799), .ZN(n1659) );
NAND2_X1 U1398 ( .A1(n1800), .A2(n1801), .ZN(U320) );
NAND2_X1 U1399 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1658), .ZN(n1801) );
NAND2_X1 U1400 ( .A1(n1797), .A2(DATA_IN_7_), .ZN(n1800) );
NAND2_X1 U1401 ( .A1(n1803), .A2(n1804), .ZN(U319) );
NAND2_X1 U1402 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1658), .ZN(n1804) );
NAND2_X1 U1403 ( .A1(n1797), .A2(DATA_IN_6_), .ZN(n1803) );
NAND2_X1 U1404 ( .A1(n1805), .A2(n1806), .ZN(U318) );
NAND2_X1 U1405 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1658), .ZN(n1806) );
NAND2_X1 U1406 ( .A1(n1797), .A2(DATA_IN_5_), .ZN(n1805) );
NAND2_X1 U1407 ( .A1(n1807), .A2(n1808), .ZN(U317) );
NAND2_X1 U1408 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1658), .ZN(n1808) );
NAND2_X1 U1409 ( .A1(n1797), .A2(DATA_IN_4_), .ZN(n1807) );
NAND2_X1 U1410 ( .A1(n1809), .A2(n1810), .ZN(U316) );
NAND2_X1 U1411 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1658), .ZN(n1810) );
NAND2_X1 U1412 ( .A1(n1797), .A2(DATA_IN_3_), .ZN(n1809) );
NAND2_X1 U1413 ( .A1(n1811), .A2(n1812), .ZN(U315) );
NAND2_X1 U1414 ( .A1(n1813), .A2(DATA_IN_2_), .ZN(n1812) );
XOR2_X1 U1415 ( .A(n1814), .B(KEYINPUT8), .Z(n1813) );
NAND2_X1 U1416 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1658), .ZN(n1811) );
NAND2_X1 U1417 ( .A1(n1815), .A2(n1816), .ZN(U314) );
NAND2_X1 U1418 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1658), .ZN(n1816) );
NAND2_X1 U1419 ( .A1(n1797), .A2(DATA_IN_1_), .ZN(n1815) );
NAND2_X1 U1420 ( .A1(n1817), .A2(n1818), .ZN(U313) );
NAND2_X1 U1421 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1658), .ZN(n1818) );
NAND2_X1 U1422 ( .A1(n1797), .A2(DATA_IN_0_), .ZN(n1817) );
NAND2_X1 U1423 ( .A1(n1819), .A2(n1820), .ZN(U312) );
NAND2_X1 U1424 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1658), .ZN(n1820) );
NAND2_X1 U1425 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1797), .ZN(n1819) );
NAND2_X1 U1426 ( .A1(n1821), .A2(n1822), .ZN(U311) );
NAND2_X1 U1427 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1658), .ZN(n1822) );
NAND2_X1 U1428 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1797), .ZN(n1821) );
NAND2_X1 U1429 ( .A1(n1823), .A2(n1824), .ZN(U310) );
NAND2_X1 U1430 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1658), .ZN(n1824) );
XOR2_X1 U1431 ( .A(n1825), .B(KEYINPUT28), .Z(n1823) );
NAND2_X1 U1432 ( .A1(n1797), .A2(n1826), .ZN(n1825) );
XOR2_X1 U1433 ( .A(REG1_REG_5__SCAN_IN), .B(KEYINPUT43), .Z(n1826) );
NAND2_X1 U1434 ( .A1(n1827), .A2(n1828), .ZN(U309) );
NAND2_X1 U1435 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1658), .ZN(n1828) );
NAND2_X1 U1436 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1797), .ZN(n1827) );
NAND2_X1 U1437 ( .A1(n1829), .A2(n1830), .ZN(U308) );
NAND2_X1 U1438 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1797), .ZN(n1830) );
XOR2_X1 U1439 ( .A(KEYINPUT44), .B(n1831), .Z(n1829) );
AND2_X1 U1440 ( .A1(n1658), .A2(REG2_REG_3__SCAN_IN), .ZN(n1831) );
NAND2_X1 U1441 ( .A1(n1832), .A2(n1833), .ZN(U307) );
NAND2_X1 U1442 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1658), .ZN(n1833) );
NAND2_X1 U1443 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1797), .ZN(n1832) );
NAND2_X1 U1444 ( .A1(n1834), .A2(n1835), .ZN(U306) );
NAND2_X1 U1445 ( .A1(n1797), .A2(n1836), .ZN(n1835) );
XOR2_X1 U1446 ( .A(REG1_REG_1__SCAN_IN), .B(KEYINPUT19), .Z(n1836) );
NAND2_X1 U1447 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1658), .ZN(n1834) );
NAND2_X1 U1448 ( .A1(n1837), .A2(n1838), .ZN(U305) );
NAND2_X1 U1449 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1839), .ZN(n1838) );
XOR2_X1 U1450 ( .A(KEYINPUT45), .B(n1797), .Z(n1839) );
NAND2_X1 U1451 ( .A1(n1840), .A2(REG2_REG_0__SCAN_IN), .ZN(n1837) );
XNOR2_X1 U1452 ( .A(n1657), .B(KEYINPUT38), .ZN(n1840) );
NAND2_X1 U1453 ( .A1(n1841), .A2(n1842), .ZN(U304) );
NAND2_X1 U1454 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1843), .ZN(n1842) );
XOR2_X1 U1455 ( .A(KEYINPUT63), .B(n1657), .Z(n1843) );
NAND2_X1 U1456 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1797), .ZN(n1841) );
NAND2_X1 U1457 ( .A1(n1844), .A2(n1845), .ZN(U303) );
NAND2_X1 U1458 ( .A1(n1846), .A2(n1658), .ZN(n1845) );
XOR2_X1 U1459 ( .A(REG3_REG_6__SCAN_IN), .B(KEYINPUT54), .Z(n1846) );
NAND2_X1 U1460 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1797), .ZN(n1844) );
NAND2_X1 U1461 ( .A1(n1847), .A2(n1848), .ZN(U302) );
NAND2_X1 U1462 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1658), .ZN(n1848) );
NAND2_X1 U1463 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1797), .ZN(n1847) );
NAND2_X1 U1464 ( .A1(n1849), .A2(n1850), .ZN(U301) );
NAND2_X1 U1465 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1658), .ZN(n1850) );
NAND2_X1 U1466 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1797), .ZN(n1849) );
NAND2_X1 U1467 ( .A1(n1851), .A2(n1852), .ZN(U300) );
NAND2_X1 U1468 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1658), .ZN(n1852) );
NAND2_X1 U1469 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1797), .ZN(n1851) );
NAND2_X1 U1470 ( .A1(n1853), .A2(n1854), .ZN(U299) );
NAND2_X1 U1471 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1658), .ZN(n1854) );
NAND2_X1 U1472 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1797), .ZN(n1853) );
NAND2_X1 U1473 ( .A1(n1855), .A2(n1856), .ZN(U298) );
NAND2_X1 U1474 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1657), .ZN(n1856) );
NAND2_X1 U1475 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1797), .ZN(n1855) );
NAND2_X1 U1476 ( .A1(n1857), .A2(n1858), .ZN(U297) );
NAND2_X1 U1477 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1657), .ZN(n1858) );
NAND2_X1 U1478 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1797), .ZN(n1857) );
NAND2_X1 U1479 ( .A1(n1859), .A2(n1860), .ZN(U296) );
NAND2_X1 U1480 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1657), .ZN(n1860) );
NAND2_X1 U1481 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1797), .ZN(n1859) );
NAND2_X1 U1482 ( .A1(n1861), .A2(n1862), .ZN(U295) );
NAND2_X1 U1483 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1657), .ZN(n1862) );
NAND2_X1 U1484 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1797), .ZN(n1861) );
NAND2_X1 U1485 ( .A1(n1863), .A2(n1864), .ZN(U294) );
NAND2_X1 U1486 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1657), .ZN(n1864) );
NAND2_X1 U1487 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1797), .ZN(n1863) );
NAND2_X1 U1488 ( .A1(n1865), .A2(n1866), .ZN(U293) );
NAND2_X1 U1489 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1657), .ZN(n1866) );
NAND2_X1 U1490 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1797), .ZN(n1865) );
NAND2_X1 U1491 ( .A1(n1867), .A2(n1868), .ZN(U292) );
NAND2_X1 U1492 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1657), .ZN(n1868) );
NAND2_X1 U1493 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1797), .ZN(n1867) );
NAND2_X1 U1494 ( .A1(n1869), .A2(n1870), .ZN(U291) );
NAND2_X1 U1495 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1657), .ZN(n1870) );
NAND2_X1 U1496 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1797), .ZN(n1869) );
NAND2_X1 U1497 ( .A1(n1871), .A2(n1872), .ZN(U290) );
NAND2_X1 U1498 ( .A1(n1797), .A2(n1873), .ZN(n1872) );
XOR2_X1 U1499 ( .A(REG3_REG_1__SCAN_IN), .B(KEYINPUT1), .Z(n1873) );
NAND2_X1 U1500 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1657), .ZN(n1871) );
NAND2_X1 U1501 ( .A1(n1874), .A2(n1875), .ZN(U289) );
NAND2_X1 U1502 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1657), .ZN(n1875) );
NAND2_X1 U1503 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1797), .ZN(n1874) );
NAND4_X1 U1504 ( .A1(n1876), .A2(n1877), .A3(n1878), .A4(n1879), .ZN(U288));
NAND2_X1 U1505 ( .A1(n1880), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1879) );
NAND2_X1 U1506 ( .A1(n1881), .A2(REG4_REG_7__SCAN_IN), .ZN(n1878) );
NAND2_X1 U1507 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1657), .ZN(n1877) );
NAND4_X1 U1508 ( .A1(n1882), .A2(n1883), .A3(n1876), .A4(n1884), .ZN(U287));
NOR3_X1 U1509 ( .A1(n1885), .A2(n1886), .A3(n1887), .ZN(n1884) );
NOR3_X1 U1510 ( .A1(n1888), .A2(n1889), .A3(n1890), .ZN(n1887) );
NOR3_X1 U1511 ( .A1(n1891), .A2(n1892), .A3(n1893), .ZN(n1886) );
XOR2_X1 U1512 ( .A(n1894), .B(KEYINPUT29), .Z(n1893) );
NOR2_X1 U1513 ( .A1(n1895), .A2(n1896), .ZN(n1885) );
XNOR2_X1 U1514 ( .A(RLAST_REG_6__SCAN_IN), .B(KEYINPUT16), .ZN(n1895) );
NAND2_X1 U1515 ( .A1(n1881), .A2(REG4_REG_6__SCAN_IN), .ZN(n1883) );
NAND2_X1 U1516 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1657), .ZN(n1882) );
NAND4_X1 U1517 ( .A1(n1897), .A2(n1898), .A3(n1876), .A4(n1899), .ZN(U286));
NOR4_X1 U1518 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(n1899));
AND2_X1 U1519 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1880), .ZN(n1903) );
NOR2_X1 U1520 ( .A1(n1904), .A2(n1905), .ZN(n1902) );
NOR3_X1 U1521 ( .A1(n1891), .A2(n1906), .A3(n1907), .ZN(n1901) );
NOR2_X1 U1522 ( .A1(n1908), .A2(n1909), .ZN(n1907) );
INV_X1 U1523 ( .A(n1894), .ZN(n1906) );
NOR3_X1 U1524 ( .A1(n1890), .A2(n1910), .A3(n1911), .ZN(n1900) );
NOR2_X1 U1525 ( .A1(n1908), .A2(n1912), .ZN(n1911) );
INV_X1 U1526 ( .A(n1888), .ZN(n1910) );
AND2_X1 U1527 ( .A1(n1913), .A2(n1914), .ZN(n1876) );
NAND3_X1 U1528 ( .A1(n1915), .A2(n1888), .A3(n1889), .ZN(n1914) );
NAND2_X1 U1529 ( .A1(n1916), .A2(n1917), .ZN(n1888) );
OR2_X1 U1530 ( .A1(n1889), .A2(n1908), .ZN(n1917) );
AND2_X1 U1531 ( .A1(n1918), .A2(n1919), .ZN(n1889) );
XNOR2_X1 U1532 ( .A(KEYINPUT2), .B(n1904), .ZN(n1919) );
XOR2_X1 U1533 ( .A(n1920), .B(KEYINPUT41), .Z(n1918) );
XOR2_X1 U1534 ( .A(KEYINPUT52), .B(n1912), .Z(n1916) );
NAND3_X1 U1535 ( .A1(n1892), .A2(n1894), .A3(n1921), .ZN(n1913) );
INV_X1 U1536 ( .A(n1891), .ZN(n1921) );
NAND2_X1 U1537 ( .A1(n1909), .A2(n1922), .ZN(n1894) );
OR2_X1 U1538 ( .A1(n1892), .A2(n1908), .ZN(n1922) );
NOR2_X1 U1539 ( .A1(n1904), .A2(n1923), .ZN(n1908) );
AND2_X1 U1540 ( .A1(n1923), .A2(n1904), .ZN(n1892) );
NAND2_X1 U1541 ( .A1(n1924), .A2(n1925), .ZN(n1904) );
NAND4_X1 U1542 ( .A1(n1926), .A2(n1927), .A3(n1928), .A4(n1929), .ZN(n1925));
NAND2_X1 U1543 ( .A1(n1930), .A2(n1931), .ZN(n1929) );
INV_X1 U1544 ( .A(n1932), .ZN(n1930) );
NAND2_X1 U1545 ( .A1(n1933), .A2(n1932), .ZN(n1928) );
XOR2_X1 U1546 ( .A(KEYINPUT36), .B(n1934), .Z(n1933) );
NAND2_X1 U1547 ( .A1(n1935), .A2(n1936), .ZN(n1927) );
NAND4_X1 U1548 ( .A1(n1935), .A2(n1937), .A3(n1938), .A4(n1939), .ZN(n1924));
NAND2_X1 U1549 ( .A1(n1934), .A2(n1932), .ZN(n1939) );
XNOR2_X1 U1550 ( .A(n1931), .B(KEYINPUT40), .ZN(n1934) );
OR2_X1 U1551 ( .A1(n1932), .A2(n1931), .ZN(n1938) );
NAND2_X1 U1552 ( .A1(n1940), .A2(n1941), .ZN(n1931) );
NAND2_X1 U1553 ( .A1(DATA_IN_6_), .A2(n1942), .ZN(n1941) );
NAND2_X1 U1554 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1940) );
NAND2_X1 U1555 ( .A1(n1943), .A2(n1944), .ZN(n1932) );
NAND2_X1 U1556 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1942), .ZN(n1944) );
NAND2_X1 U1557 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1943) );
NAND2_X1 U1558 ( .A1(n1945), .A2(n1926), .ZN(n1937) );
NAND2_X1 U1559 ( .A1(n1946), .A2(n1947), .ZN(n1926) );
NAND2_X1 U1560 ( .A1(n1948), .A2(n1949), .ZN(n1935) );
INV_X1 U1561 ( .A(n1920), .ZN(n1923) );
NAND2_X1 U1562 ( .A1(n1881), .A2(REG4_REG_5__SCAN_IN), .ZN(n1898) );
NAND2_X1 U1563 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1657), .ZN(n1897) );
NAND4_X1 U1564 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(U285));
NOR3_X1 U1565 ( .A1(n1954), .A2(n1955), .A3(n1956), .ZN(n1953) );
NOR3_X1 U1566 ( .A1(n1890), .A2(n1912), .A3(n1957), .ZN(n1956) );
NOR2_X1 U1567 ( .A1(n1958), .A2(n1959), .ZN(n1957) );
NOR2_X1 U1568 ( .A1(n1960), .A2(n1961), .ZN(n1958) );
AND3_X1 U1569 ( .A1(n1959), .A2(n1962), .A3(n1963), .ZN(n1912) );
NOR3_X1 U1570 ( .A1(n1891), .A2(n1909), .A3(n1964), .ZN(n1955) );
NOR2_X1 U1571 ( .A1(n1965), .A2(n1966), .ZN(n1964) );
NOR2_X1 U1572 ( .A1(n1967), .A2(n1968), .ZN(n1965) );
NOR3_X1 U1573 ( .A1(n1968), .A2(n1967), .A3(n1969), .ZN(n1909) );
NOR3_X1 U1574 ( .A1(n1970), .A2(KEYINPUT6), .A3(n1971), .ZN(n1967) );
NOR2_X1 U1575 ( .A1(n1972), .A2(n1959), .ZN(n1968) );
NAND2_X1 U1576 ( .A1(n1920), .A2(n1973), .ZN(n1959) );
NAND2_X1 U1577 ( .A1(n1974), .A2(n1975), .ZN(n1973) );
NAND2_X1 U1578 ( .A1(n1970), .A2(n1971), .ZN(n1920) );
INV_X1 U1579 ( .A(KEYINPUT6), .ZN(n1972) );
NOR2_X1 U1580 ( .A1(n1971), .A2(n1905), .ZN(n1954) );
INV_X1 U1581 ( .A(n1974), .ZN(n1971) );
NAND2_X1 U1582 ( .A1(n1976), .A2(n1977), .ZN(n1974) );
NAND4_X1 U1583 ( .A1(n1978), .A2(n1979), .A3(n1980), .A4(n1949), .ZN(n1977));
NAND2_X1 U1584 ( .A1(n1948), .A2(n1981), .ZN(n1980) );
OR3_X1 U1585 ( .A1(n1981), .A2(n1948), .A3(KEYINPUT48), .ZN(n1979) );
INV_X1 U1586 ( .A(n1982), .ZN(n1981) );
NAND2_X1 U1587 ( .A1(KEYINPUT48), .A2(n1945), .ZN(n1978) );
NAND2_X1 U1588 ( .A1(n1983), .A2(n1946), .ZN(n1976) );
INV_X1 U1589 ( .A(n1949), .ZN(n1946) );
NAND2_X1 U1590 ( .A1(n1984), .A2(n1985), .ZN(n1949) );
NAND2_X1 U1591 ( .A1(n1986), .A2(n1987), .ZN(n1985) );
NAND2_X1 U1592 ( .A1(n1988), .A2(n1989), .ZN(n1987) );
NAND2_X1 U1593 ( .A1(n1990), .A2(n1991), .ZN(n1984) );
XOR2_X1 U1594 ( .A(n1948), .B(n1982), .Z(n1983) );
NOR2_X1 U1595 ( .A1(n1945), .A2(KEYINPUT49), .ZN(n1982) );
INV_X1 U1596 ( .A(n1936), .ZN(n1945) );
NAND2_X1 U1597 ( .A1(n1992), .A2(n1993), .ZN(n1936) );
NAND2_X1 U1598 ( .A1(DATA_IN_5_), .A2(n1942), .ZN(n1993) );
NAND2_X1 U1599 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1992) );
INV_X1 U1600 ( .A(n1947), .ZN(n1948) );
NAND2_X1 U1601 ( .A1(n1994), .A2(n1995), .ZN(n1947) );
NAND2_X1 U1602 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1942), .ZN(n1995) );
NAND2_X1 U1603 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1994) );
NAND2_X1 U1604 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1657), .ZN(n1952) );
NAND2_X1 U1605 ( .A1(n1880), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1951) );
NAND2_X1 U1606 ( .A1(n1881), .A2(REG4_REG_4__SCAN_IN), .ZN(n1950) );
NAND4_X1 U1607 ( .A1(n1996), .A2(n1997), .A3(n1998), .A4(n1999), .ZN(U284));
NOR3_X1 U1608 ( .A1(n2000), .A2(n2001), .A3(n2002), .ZN(n1999) );
NOR2_X1 U1609 ( .A1(n1890), .A2(n2003), .ZN(n2002) );
XOR2_X1 U1610 ( .A(n1961), .B(n1962), .Z(n2003) );
NOR3_X1 U1611 ( .A1(n1891), .A2(n1966), .A3(n2004), .ZN(n2001) );
XOR2_X1 U1612 ( .A(n2005), .B(KEYINPUT26), .Z(n2004) );
NAND2_X1 U1613 ( .A1(n1960), .A2(n2006), .ZN(n2005) );
XOR2_X1 U1614 ( .A(KEYINPUT62), .B(n2007), .Z(n2006) );
INV_X1 U1615 ( .A(n1962), .ZN(n1960) );
INV_X1 U1616 ( .A(n1969), .ZN(n1966) );
NAND2_X1 U1617 ( .A1(n2007), .A2(n1962), .ZN(n1969) );
NAND2_X1 U1618 ( .A1(n1975), .A2(n2008), .ZN(n1962) );
NAND2_X1 U1619 ( .A1(n2009), .A2(n2010), .ZN(n2008) );
INV_X1 U1620 ( .A(n1970), .ZN(n1975) );
NOR2_X1 U1621 ( .A1(n2010), .A2(n2009), .ZN(n1970) );
NOR2_X1 U1622 ( .A1(n2011), .A2(n1905), .ZN(n2000) );
INV_X1 U1623 ( .A(n2009), .ZN(n2011) );
NAND2_X1 U1624 ( .A1(n2012), .A2(n2013), .ZN(n2009) );
NAND2_X1 U1625 ( .A1(n2014), .A2(n1991), .ZN(n2013) );
NAND2_X1 U1626 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
NAND2_X1 U1627 ( .A1(n1986), .A2(n1989), .ZN(n2016) );
XOR2_X1 U1628 ( .A(KEYINPUT46), .B(n2017), .Z(n2015) );
NOR2_X1 U1629 ( .A1(n1986), .A2(n2018), .ZN(n2017) );
NAND2_X1 U1630 ( .A1(n2019), .A2(n1988), .ZN(n2012) );
INV_X1 U1631 ( .A(n1991), .ZN(n1988) );
NAND2_X1 U1632 ( .A1(n2020), .A2(n2021), .ZN(n1991) );
NAND2_X1 U1633 ( .A1(n2022), .A2(n2023), .ZN(n2021) );
NAND2_X1 U1634 ( .A1(n2024), .A2(n2025), .ZN(n2023) );
OR2_X1 U1635 ( .A1(n2024), .A2(n2025), .ZN(n2020) );
NAND2_X1 U1636 ( .A1(n2026), .A2(n2027), .ZN(n2019) );
NAND2_X1 U1637 ( .A1(n1986), .A2(n2028), .ZN(n2027) );
NAND2_X1 U1638 ( .A1(KEYINPUT58), .A2(n1989), .ZN(n2028) );
INV_X1 U1639 ( .A(n2029), .ZN(n1986) );
NAND3_X1 U1640 ( .A1(n2030), .A2(n2031), .A3(n2029), .ZN(n2026) );
NAND2_X1 U1641 ( .A1(n2032), .A2(n2033), .ZN(n2029) );
NAND2_X1 U1642 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1942), .ZN(n2033) );
NAND2_X1 U1643 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2032) );
OR2_X1 U1644 ( .A1(n1990), .A2(KEYINPUT58), .ZN(n2031) );
XNOR2_X1 U1645 ( .A(KEYINPUT55), .B(n2018), .ZN(n2030) );
XNOR2_X1 U1646 ( .A(n1990), .B(KEYINPUT42), .ZN(n2018) );
INV_X1 U1647 ( .A(n1989), .ZN(n1990) );
NAND2_X1 U1648 ( .A1(n2034), .A2(n2035), .ZN(n1989) );
NAND2_X1 U1649 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2035) );
XOR2_X1 U1650 ( .A(KEYINPUT61), .B(n2036), .Z(n2034) );
AND2_X1 U1651 ( .A1(n1942), .A2(DATA_IN_4_), .ZN(n2036) );
NAND2_X1 U1652 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1657), .ZN(n1998) );
NAND2_X1 U1653 ( .A1(n1880), .A2(RLAST_REG_3__SCAN_IN), .ZN(n1997) );
NAND2_X1 U1654 ( .A1(n1881), .A2(REG4_REG_3__SCAN_IN), .ZN(n1996) );
NAND4_X1 U1655 ( .A1(n2037), .A2(n2038), .A3(n2039), .A4(n2040), .ZN(U283));
NOR3_X1 U1656 ( .A1(n2041), .A2(n2042), .A3(n2043), .ZN(n2040) );
NOR3_X1 U1657 ( .A1(n1891), .A2(n2007), .A3(n2044), .ZN(n2043) );
NOR2_X1 U1658 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
AND2_X1 U1659 ( .A1(n2047), .A2(n2048), .ZN(n2045) );
AND3_X1 U1660 ( .A1(n2047), .A2(n2046), .A3(n2048), .ZN(n2007) );
NOR3_X1 U1661 ( .A1(n1890), .A2(n1963), .A3(n2049), .ZN(n2042) );
NOR2_X1 U1662 ( .A1(n2050), .A2(n2046), .ZN(n2049) );
NOR2_X1 U1663 ( .A1(n2051), .A2(n2052), .ZN(n2050) );
INV_X1 U1664 ( .A(n1961), .ZN(n1963) );
NAND3_X1 U1665 ( .A1(n2053), .A2(n2054), .A3(n2046), .ZN(n1961) );
NAND2_X1 U1666 ( .A1(n2010), .A2(n2055), .ZN(n2046) );
NAND2_X1 U1667 ( .A1(n2056), .A2(n2057), .ZN(n2055) );
OR2_X1 U1668 ( .A1(n2057), .A2(n2056), .ZN(n2010) );
NOR2_X1 U1669 ( .A1(n2058), .A2(n1905), .ZN(n2041) );
INV_X1 U1670 ( .A(n2056), .ZN(n2058) );
XOR2_X1 U1671 ( .A(n2025), .B(n2059), .Z(n2056) );
XNOR2_X1 U1672 ( .A(n2024), .B(n2022), .ZN(n2059) );
AND2_X1 U1673 ( .A1(n2060), .A2(n2061), .ZN(n2022) );
NAND2_X1 U1674 ( .A1(DATA_IN_3_), .A2(n1942), .ZN(n2061) );
NAND2_X1 U1675 ( .A1(RESTART), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2060) );
NAND2_X1 U1676 ( .A1(n2062), .A2(n2063), .ZN(n2024) );
NAND2_X1 U1677 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1942), .ZN(n2063) );
NAND2_X1 U1678 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2062) );
NAND2_X1 U1679 ( .A1(n2064), .A2(n2065), .ZN(n2025) );
NAND2_X1 U1680 ( .A1(n2066), .A2(n2067), .ZN(n2065) );
NAND2_X1 U1681 ( .A1(n2068), .A2(n2069), .ZN(n2066) );
NAND2_X1 U1682 ( .A1(n2070), .A2(n2071), .ZN(n2064) );
NAND2_X1 U1683 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1657), .ZN(n2039) );
NAND2_X1 U1684 ( .A1(n1880), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2038) );
NAND2_X1 U1685 ( .A1(n1881), .A2(REG4_REG_2__SCAN_IN), .ZN(n2037) );
NAND4_X1 U1686 ( .A1(n2072), .A2(n2073), .A3(n2074), .A4(n2075), .ZN(U282));
NOR3_X1 U1687 ( .A1(n2076), .A2(n2077), .A3(n2078), .ZN(n2075) );
NOR2_X1 U1688 ( .A1(n2079), .A2(n1890), .ZN(n2078) );
NOR2_X1 U1689 ( .A1(n2080), .A2(n2081), .ZN(n2079) );
XOR2_X1 U1690 ( .A(KEYINPUT34), .B(n2082), .Z(n2081) );
NOR2_X1 U1691 ( .A1(n2052), .A2(n2054), .ZN(n2082) );
INV_X1 U1692 ( .A(n2053), .ZN(n2052) );
NOR2_X1 U1693 ( .A1(n2051), .A2(n2053), .ZN(n2080) );
NAND2_X1 U1694 ( .A1(n2057), .A2(n2083), .ZN(n2053) );
NAND2_X1 U1695 ( .A1(n2084), .A2(n2085), .ZN(n2083) );
NOR2_X1 U1696 ( .A1(n2086), .A2(n1891), .ZN(n2077) );
XNOR2_X1 U1697 ( .A(n2048), .B(n2047), .ZN(n2086) );
NAND3_X1 U1698 ( .A1(n2087), .A2(n2088), .A3(n2057), .ZN(n2048) );
NAND2_X1 U1699 ( .A1(n2089), .A2(n2090), .ZN(n2057) );
NAND3_X1 U1700 ( .A1(KEYINPUT3), .A2(n2084), .A3(n2085), .ZN(n2088) );
INV_X1 U1701 ( .A(n2090), .ZN(n2084) );
OR2_X1 U1702 ( .A1(n2085), .A2(KEYINPUT3), .ZN(n2087) );
NOR2_X1 U1703 ( .A1(n2090), .A2(n1905), .ZN(n2076) );
XOR2_X1 U1704 ( .A(n2067), .B(n2091), .Z(n2090) );
NOR2_X1 U1705 ( .A1(n2092), .A2(n2093), .ZN(n2091) );
NOR3_X1 U1706 ( .A1(n2071), .A2(KEYINPUT59), .A3(n2069), .ZN(n2093) );
NOR2_X1 U1707 ( .A1(n2068), .A2(n2070), .ZN(n2092) );
INV_X1 U1708 ( .A(n2069), .ZN(n2070) );
NAND2_X1 U1709 ( .A1(n2094), .A2(n2095), .ZN(n2069) );
NAND2_X1 U1710 ( .A1(n2096), .A2(n2097), .ZN(n2095) );
NAND2_X1 U1711 ( .A1(n2098), .A2(n2099), .ZN(n2097) );
OR2_X1 U1712 ( .A1(n2099), .A2(n2098), .ZN(n2094) );
INV_X1 U1713 ( .A(n2071), .ZN(n2068) );
NAND2_X1 U1714 ( .A1(n2100), .A2(n2101), .ZN(n2071) );
NAND2_X1 U1715 ( .A1(DATA_IN_2_), .A2(n1942), .ZN(n2101) );
NAND2_X1 U1716 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2100) );
NAND2_X1 U1717 ( .A1(n2102), .A2(n2103), .ZN(n2067) );
NAND2_X1 U1718 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1942), .ZN(n2103) );
XOR2_X1 U1719 ( .A(n2104), .B(KEYINPUT57), .Z(n2102) );
NAND2_X1 U1720 ( .A1(n2105), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2104) );
XNOR2_X1 U1721 ( .A(RESTART), .B(KEYINPUT51), .ZN(n2105) );
NAND2_X1 U1722 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1657), .ZN(n2074) );
NAND2_X1 U1723 ( .A1(n1880), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2073) );
NAND2_X1 U1724 ( .A1(n1881), .A2(REG4_REG_1__SCAN_IN), .ZN(n2072) );
INV_X1 U1725 ( .A(n2106), .ZN(n1881) );
NAND4_X1 U1726 ( .A1(n2107), .A2(n2108), .A3(n2109), .A4(n2110), .ZN(U281));
NOR3_X1 U1727 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n2110) );
NOR2_X1 U1728 ( .A1(n2114), .A2(n1905), .ZN(n2113) );
NAND3_X1 U1729 ( .A1(n2115), .A2(n2116), .A3(n2117), .ZN(n1905) );
NAND2_X1 U1730 ( .A1(n2118), .A2(n2119), .ZN(n2116) );
XNOR2_X1 U1731 ( .A(RESTART), .B(KEYINPUT11), .ZN(n2118) );
NAND2_X1 U1732 ( .A1(n1942), .A2(n2120), .ZN(n2115) );
NAND4_X1 U1733 ( .A1(n2121), .A2(ENABLE), .A3(n2122), .A4(n2123), .ZN(n2120));
AND2_X1 U1734 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1880), .ZN(n2112) );
INV_X1 U1735 ( .A(n1896), .ZN(n1880) );
NAND3_X1 U1736 ( .A1(n1942), .A2(n1798), .A3(n2117), .ZN(n1896) );
INV_X1 U1737 ( .A(ENABLE), .ZN(n1798) );
NOR2_X1 U1738 ( .A1(n2124), .A2(n2106), .ZN(n2111) );
NAND2_X1 U1739 ( .A1(AVERAGE), .A2(n2125), .ZN(n2106) );
OR2_X1 U1740 ( .A1(n2047), .A2(n1891), .ZN(n2109) );
NAND3_X1 U1741 ( .A1(n2126), .A2(n2123), .A3(n2125), .ZN(n1891) );
AND3_X1 U1742 ( .A1(n2117), .A2(n1942), .A3(ENABLE), .ZN(n2125) );
INV_X1 U1743 ( .A(AVERAGE), .ZN(n2123) );
NAND2_X1 U1744 ( .A1(n2121), .A2(n2122), .ZN(n2126) );
NAND3_X1 U1745 ( .A1(n2127), .A2(n2128), .A3(n2129), .ZN(n2122) );
OR2_X1 U1746 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2129) );
NAND2_X1 U1747 ( .A1(n2130), .A2(n2131), .ZN(n2128) );
OR2_X1 U1748 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2131) );
NAND2_X1 U1749 ( .A1(n2132), .A2(n2133), .ZN(n2130) );
NAND2_X1 U1750 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2133) );
NAND2_X1 U1751 ( .A1(n2134), .A2(n2135), .ZN(n2132) );
NAND2_X1 U1752 ( .A1(n2136), .A2(n2137), .ZN(n2135) );
NAND3_X1 U1753 ( .A1(n2138), .A2(n2139), .A3(n2140), .ZN(n2137) );
OR2_X1 U1754 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2140) );
NAND3_X1 U1755 ( .A1(n2141), .A2(n2142), .A3(n2143), .ZN(n2139) );
XOR2_X1 U1756 ( .A(KEYINPUT25), .B(n2144), .Z(n2143) );
NOR3_X1 U1757 ( .A1(n2145), .A2(n2146), .A3(n2147), .ZN(n2144) );
NOR2_X1 U1758 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2148), .ZN(n2147) );
XOR2_X1 U1759 ( .A(KEYINPUT23), .B(DATA_IN_1_), .Z(n2148) );
NOR2_X1 U1760 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2146) );
NOR2_X1 U1761 ( .A1(n2149), .A2(n2150), .ZN(n2145) );
AND2_X1 U1762 ( .A1(DATA_IN_1_), .A2(REG4_REG_1__SCAN_IN), .ZN(n2150) );
NOR2_X1 U1763 ( .A1(n1686), .A2(n2124), .ZN(n2149) );
INV_X1 U1764 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2124) );
INV_X1 U1765 ( .A(DATA_IN_0_), .ZN(n1686) );
NAND2_X1 U1766 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2142) );
NAND2_X1 U1767 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2141) );
OR2_X1 U1768 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2138) );
NAND2_X1 U1769 ( .A1(n2151), .A2(REG4_REG_4__SCAN_IN), .ZN(n2136) );
XOR2_X1 U1770 ( .A(n1671), .B(KEYINPUT30), .Z(n2151) );
INV_X1 U1771 ( .A(DATA_IN_4_), .ZN(n1671) );
OR2_X1 U1772 ( .A1(DATA_IN_5_), .A2(REG4_REG_5__SCAN_IN), .ZN(n2134) );
NAND2_X1 U1773 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2127) );
XOR2_X1 U1774 ( .A(n2152), .B(KEYINPUT33), .Z(n2121) );
NAND2_X1 U1775 ( .A1(DATA_IN_7_), .A2(n2153), .ZN(n2152) );
XOR2_X1 U1776 ( .A(REG4_REG_7__SCAN_IN), .B(KEYINPUT10), .Z(n2153) );
NAND2_X1 U1777 ( .A1(n2154), .A2(n2155), .ZN(n2047) );
NAND2_X1 U1778 ( .A1(n2156), .A2(n2157), .ZN(n2155) );
NAND2_X1 U1779 ( .A1(n2114), .A2(n2158), .ZN(n2157) );
NAND2_X1 U1780 ( .A1(n2089), .A2(n2158), .ZN(n2154) );
INV_X1 U1781 ( .A(KEYINPUT0), .ZN(n2158) );
NAND2_X1 U1782 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1657), .ZN(n2108) );
NAND2_X1 U1783 ( .A1(n2051), .A2(n1915), .ZN(n2107) );
INV_X1 U1784 ( .A(n1890), .ZN(n1915) );
NAND3_X1 U1785 ( .A1(n2117), .A2(RESTART), .A3(n2159), .ZN(n1890) );
XOR2_X1 U1786 ( .A(n2119), .B(KEYINPUT13), .Z(n2159) );
NAND2_X1 U1787 ( .A1(n2160), .A2(n2161), .ZN(n2119) );
NAND2_X1 U1788 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n2162), .ZN(n2161) );
OR2_X1 U1789 ( .A1(n2163), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2162) );
NAND2_X1 U1790 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n2163), .ZN(n2160) );
NAND2_X1 U1791 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
NAND3_X1 U1792 ( .A1(n2166), .A2(n2167), .A3(n2168), .ZN(n2165) );
NAND2_X1 U1793 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2168) );
NAND2_X1 U1794 ( .A1(n2169), .A2(n2170), .ZN(n2167) );
NAND2_X1 U1795 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
NAND3_X1 U1796 ( .A1(n2173), .A2(n2174), .A3(n2175), .ZN(n2172) );
OR2_X1 U1797 ( .A1(RMAX_REG_4__SCAN_IN), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2175) );
NAND3_X1 U1798 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(n2174) );
NAND2_X1 U1799 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2178) );
NAND3_X1 U1800 ( .A1(n2179), .A2(n2180), .A3(n2181), .ZN(n2177) );
NAND2_X1 U1801 ( .A1(n1764), .A2(n1731), .ZN(n2181) );
INV_X1 U1802 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1731) );
INV_X1 U1803 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1764) );
NAND2_X1 U1804 ( .A1(n2182), .A2(n1737), .ZN(n2180) );
INV_X1 U1805 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1737) );
OR2_X1 U1806 ( .A1(n2183), .A2(n1772), .ZN(n2182) );
NAND2_X1 U1807 ( .A1(n2183), .A2(n1772), .ZN(n2179) );
INV_X1 U1808 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1772) );
NAND2_X1 U1809 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2183) );
NAND2_X1 U1810 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2176) );
OR2_X1 U1811 ( .A1(RMAX_REG_3__SCAN_IN), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2173) );
NAND2_X1 U1812 ( .A1(n2184), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2171) );
XNOR2_X1 U1813 ( .A(RMAX_REG_4__SCAN_IN), .B(KEYINPUT14), .ZN(n2184) );
OR2_X1 U1814 ( .A1(RMAX_REG_5__SCAN_IN), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2169) );
NAND2_X1 U1815 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2166) );
NAND2_X1 U1816 ( .A1(n1753), .A2(n1744), .ZN(n2164) );
INV_X1 U1817 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1744) );
INV_X1 U1818 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1753) );
AND2_X1 U1819 ( .A1(STATO_REG_1__SCAN_IN), .A2(U280), .ZN(n2117) );
INV_X1 U1820 ( .A(n2054), .ZN(n2051) );
NAND2_X1 U1821 ( .A1(n2085), .A2(n2185), .ZN(n2054) );
NAND2_X1 U1822 ( .A1(n2186), .A2(n2156), .ZN(n2185) );
INV_X1 U1823 ( .A(n2089), .ZN(n2085) );
NOR2_X1 U1824 ( .A1(n2156), .A2(n2186), .ZN(n2089) );
INV_X1 U1825 ( .A(n2114), .ZN(n2186) );
XNOR2_X1 U1826 ( .A(n2187), .B(n2099), .ZN(n2114) );
NAND2_X1 U1827 ( .A1(n2188), .A2(n2189), .ZN(n2099) );
NAND2_X1 U1828 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1942), .ZN(n2189) );
NAND2_X1 U1829 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2188) );
NAND2_X1 U1830 ( .A1(n2190), .A2(n2191), .ZN(n2187) );
NAND2_X1 U1831 ( .A1(n2096), .A2(n2098), .ZN(n2191) );
INV_X1 U1832 ( .A(n2192), .ZN(n2096) );
NAND2_X1 U1833 ( .A1(n2193), .A2(n2192), .ZN(n2190) );
NAND2_X1 U1834 ( .A1(n2194), .A2(n2195), .ZN(n2192) );
NAND2_X1 U1835 ( .A1(DATA_IN_1_), .A2(n1942), .ZN(n2195) );
NAND2_X1 U1836 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2194) );
NAND2_X1 U1837 ( .A1(KEYINPUT7), .A2(n2098), .ZN(n2193) );
AND2_X1 U1838 ( .A1(n2196), .A2(n2197), .ZN(n2098) );
XOR2_X1 U1839 ( .A(KEYINPUT17), .B(n2198), .Z(n2196) );
XOR2_X1 U1840 ( .A(n2197), .B(n2199), .Z(n2156) );
NOR2_X1 U1841 ( .A1(n2198), .A2(KEYINPUT32), .ZN(n2199) );
AND2_X1 U1842 ( .A1(n2200), .A2(n2201), .ZN(n2198) );
NAND2_X1 U1843 ( .A1(DATA_IN_0_), .A2(n1942), .ZN(n2201) );
NAND2_X1 U1844 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2200) );
NAND2_X1 U1845 ( .A1(n2202), .A2(n2203), .ZN(n2197) );
NAND2_X1 U1846 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1942), .ZN(n2203) );
NAND2_X1 U1847 ( .A1(RESTART), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2202) );
NAND2_X1 U1848 ( .A1(n1814), .A2(n2204), .ZN(U280) );
NAND2_X1 U1849 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1799), .ZN(n2204) );
INV_X1 U1850 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1799) );
NAND2_X1 U1851 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1685), .ZN(n1814) );
INV_X1 U1852 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1685) );
endmodule


