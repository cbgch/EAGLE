//Key = 0011010010101110111001011111010010011011011011000000111010001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304;

XOR2_X1 U712 ( .A(n993), .B(n994), .Z(G9) );
XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT34), .ZN(n994) );
NOR2_X1 U714 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR3_X1 U715 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NOR2_X1 U716 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U717 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
XOR2_X1 U718 ( .A(KEYINPUT6), .B(n1004), .Z(n1003) );
AND3_X1 U719 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NOR3_X1 U720 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1002) );
NOR2_X1 U721 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U722 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U723 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
XNOR2_X1 U724 ( .A(n1017), .B(KEYINPUT44), .ZN(n1016) );
NOR2_X1 U725 ( .A1(n1018), .A2(n1019), .ZN(n1011) );
NOR2_X1 U726 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NAND3_X1 U727 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n997) );
NAND2_X1 U728 ( .A1(n1006), .A2(n1025), .ZN(n1024) );
NAND2_X1 U729 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U730 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U731 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U732 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR3_X1 U733 ( .A1(n1019), .A2(n1014), .A3(n1008), .ZN(n1006) );
INV_X1 U734 ( .A(n1034), .ZN(n1014) );
NOR3_X1 U735 ( .A1(n1035), .A2(G953), .A3(G952), .ZN(n995) );
INV_X1 U736 ( .A(n1022), .ZN(n1035) );
NAND4_X1 U737 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1022) );
NOR4_X1 U738 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
XOR2_X1 U739 ( .A(n1044), .B(n1045), .Z(n1043) );
XOR2_X1 U740 ( .A(KEYINPUT63), .B(n1046), .Z(n1042) );
NOR2_X1 U741 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U742 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U743 ( .A(G475), .ZN(n1050) );
NOR2_X1 U744 ( .A1(G902), .A2(n1051), .ZN(n1049) );
XOR2_X1 U745 ( .A(n1052), .B(n1053), .Z(n1041) );
NAND2_X1 U746 ( .A1(KEYINPUT60), .A2(n1054), .ZN(n1053) );
NOR3_X1 U747 ( .A1(n1005), .A2(n1055), .A3(n1032), .ZN(n1038) );
XOR2_X1 U748 ( .A(KEYINPUT61), .B(n1056), .Z(n1036) );
XOR2_X1 U749 ( .A(n1057), .B(n1058), .Z(G72) );
NOR2_X1 U750 ( .A1(n1059), .A2(n1023), .ZN(n1058) );
NOR2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1062), .A2(n1063), .ZN(n1057) );
NAND2_X1 U753 ( .A1(n1064), .A2(n1023), .ZN(n1063) );
XNOR2_X1 U754 ( .A(n1065), .B(n1066), .ZN(n1064) );
NAND3_X1 U755 ( .A1(n1065), .A2(G900), .A3(G953), .ZN(n1062) );
XNOR2_X1 U756 ( .A(n1067), .B(n1068), .ZN(n1065) );
XOR2_X1 U757 ( .A(n1069), .B(n1070), .Z(n1068) );
INV_X1 U758 ( .A(n1071), .ZN(n1069) );
NAND2_X1 U759 ( .A1(n1072), .A2(n1073), .ZN(G69) );
NAND2_X1 U760 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U761 ( .A(n1076), .B(KEYINPUT33), .Z(n1074) );
XOR2_X1 U762 ( .A(n1077), .B(n1078), .Z(n1072) );
XOR2_X1 U763 ( .A(KEYINPUT18), .B(n1079), .Z(n1078) );
NOR2_X1 U764 ( .A1(n1076), .A2(n1080), .ZN(n1079) );
XOR2_X1 U765 ( .A(KEYINPUT55), .B(n1075), .Z(n1080) );
AND2_X1 U766 ( .A1(n1081), .A2(n1023), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1076) );
NAND2_X1 U769 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NOR2_X1 U770 ( .A1(n1087), .A2(n1023), .ZN(n1077) );
AND2_X1 U771 ( .A1(G224), .A2(G898), .ZN(n1087) );
NOR2_X1 U772 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U773 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U774 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR3_X1 U775 ( .A1(n1088), .A2(n1094), .A3(n1095), .ZN(G63) );
NOR3_X1 U776 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
NOR2_X1 U777 ( .A1(KEYINPUT45), .A2(n1099), .ZN(n1098) );
NOR2_X1 U778 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
INV_X1 U779 ( .A(n1096), .ZN(n1101) );
NOR2_X1 U780 ( .A1(n1099), .A2(n1102), .ZN(n1100) );
INV_X1 U781 ( .A(KEYINPUT45), .ZN(n1102) );
XNOR2_X1 U782 ( .A(n1097), .B(KEYINPUT8), .ZN(n1099) );
AND2_X1 U783 ( .A1(n1092), .A2(G478), .ZN(n1097) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1103), .ZN(G60) );
XNOR2_X1 U785 ( .A(n1104), .B(n1051), .ZN(n1103) );
NAND2_X1 U786 ( .A1(n1092), .A2(G475), .ZN(n1104) );
NAND2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(G6) );
OR2_X1 U788 ( .A1(n1107), .A2(G104), .ZN(n1106) );
NAND2_X1 U789 ( .A1(G104), .A2(n1108), .ZN(n1105) );
NAND2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
OR2_X1 U791 ( .A1(n1111), .A2(KEYINPUT56), .ZN(n1110) );
NAND2_X1 U792 ( .A1(KEYINPUT56), .A2(n1107), .ZN(n1109) );
NAND2_X1 U793 ( .A1(KEYINPUT41), .A2(n1112), .ZN(n1107) );
INV_X1 U794 ( .A(n1111), .ZN(n1112) );
NOR2_X1 U795 ( .A1(n1088), .A2(n1113), .ZN(G57) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U797 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U798 ( .A1(n1092), .A2(G472), .ZN(n1116) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1114) );
NAND2_X1 U800 ( .A1(KEYINPUT35), .A2(n1071), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1088), .A2(n1120), .ZN(G54) );
NOR2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U805 ( .A1(n1092), .A2(G469), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
INV_X1 U807 ( .A(KEYINPUT50), .ZN(n1126) );
XOR2_X1 U808 ( .A(n1071), .B(n1127), .Z(n1125) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U810 ( .A1(n1130), .A2(KEYINPUT14), .ZN(n1129) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U812 ( .A(n1133), .B(KEYINPUT0), .ZN(n1132) );
NAND2_X1 U813 ( .A1(KEYINPUT26), .A2(n1134), .ZN(n1133) );
NAND2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U816 ( .A(n1139), .B(KEYINPUT37), .Z(n1135) );
OR2_X1 U817 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
XNOR2_X1 U818 ( .A(n1067), .B(KEYINPUT15), .ZN(n1137) );
NOR2_X1 U819 ( .A1(n1088), .A2(n1140), .ZN(G51) );
XOR2_X1 U820 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND3_X1 U822 ( .A1(n1092), .A2(n1145), .A3(KEYINPUT36), .ZN(n1144) );
AND2_X1 U823 ( .A1(G902), .A2(n999), .ZN(n1092) );
NAND3_X1 U824 ( .A1(n1066), .A2(n1082), .A3(n1146), .ZN(n999) );
XOR2_X1 U825 ( .A(n1083), .B(KEYINPUT22), .Z(n1146) );
AND4_X1 U826 ( .A1(n1111), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1082) );
AND4_X1 U827 ( .A1(n993), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1149) );
NAND3_X1 U828 ( .A1(n1021), .A2(n1153), .A3(n1154), .ZN(n993) );
NAND2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
XOR2_X1 U830 ( .A(n1157), .B(KEYINPUT21), .Z(n1155) );
NAND3_X1 U831 ( .A1(n1154), .A2(n1153), .A3(n1020), .ZN(n1111) );
AND4_X1 U832 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1066) );
AND4_X1 U833 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1166), .A2(n1167), .ZN(n1160) );
INV_X1 U835 ( .A(n1168), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1143) );
XOR2_X1 U837 ( .A(n1171), .B(KEYINPUT49), .Z(n1169) );
AND2_X1 U838 ( .A1(G953), .A2(n1172), .ZN(n1088) );
XOR2_X1 U839 ( .A(KEYINPUT42), .B(G952), .Z(n1172) );
XOR2_X1 U840 ( .A(n1173), .B(n1165), .Z(G48) );
NAND4_X1 U841 ( .A1(n1174), .A2(n1020), .A3(n1175), .A4(n1156), .ZN(n1165) );
XNOR2_X1 U842 ( .A(G143), .B(n1158), .ZN(G45) );
NAND4_X1 U843 ( .A1(n1176), .A2(n1156), .A3(n1177), .A4(n1178), .ZN(n1158) );
XOR2_X1 U844 ( .A(n1179), .B(n1164), .Z(G42) );
NAND4_X1 U845 ( .A1(n1017), .A2(n1020), .A3(n1180), .A4(n1181), .ZN(n1164) );
XNOR2_X1 U846 ( .A(G137), .B(n1163), .ZN(G39) );
NAND3_X1 U847 ( .A1(n1175), .A2(n1034), .A3(n1180), .ZN(n1163) );
INV_X1 U848 ( .A(n1026), .ZN(n1180) );
NAND2_X1 U849 ( .A1(n1182), .A2(n1174), .ZN(n1026) );
XOR2_X1 U850 ( .A(n1183), .B(G134), .Z(G36) );
NAND2_X1 U851 ( .A1(KEYINPUT62), .A2(n1159), .ZN(n1183) );
NAND3_X1 U852 ( .A1(n1182), .A2(n1021), .A3(n1176), .ZN(n1159) );
XNOR2_X1 U853 ( .A(G131), .B(n1184), .ZN(G33) );
NOR2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR3_X1 U855 ( .A1(n1187), .A2(n1188), .A3(n1001), .ZN(n1186) );
INV_X1 U856 ( .A(KEYINPUT43), .ZN(n1187) );
NOR2_X1 U857 ( .A1(KEYINPUT43), .A2(n1168), .ZN(n1185) );
NAND2_X1 U858 ( .A1(n1188), .A2(n1182), .ZN(n1168) );
INV_X1 U859 ( .A(n1001), .ZN(n1182) );
NAND2_X1 U860 ( .A1(n1033), .A2(n1189), .ZN(n1001) );
AND2_X1 U861 ( .A1(n1176), .A2(n1020), .ZN(n1188) );
AND3_X1 U862 ( .A1(n1174), .A2(n1181), .A3(n1015), .ZN(n1176) );
XOR2_X1 U863 ( .A(n1190), .B(KEYINPUT39), .Z(n1174) );
XOR2_X1 U864 ( .A(n1162), .B(n1191), .Z(G30) );
XNOR2_X1 U865 ( .A(G128), .B(KEYINPUT59), .ZN(n1191) );
NAND4_X1 U866 ( .A1(n1175), .A2(n1021), .A3(n1192), .A4(n1156), .ZN(n1162) );
AND3_X1 U867 ( .A1(n1040), .A2(n1181), .A3(n1056), .ZN(n1175) );
INV_X1 U868 ( .A(n1193), .ZN(n1040) );
XOR2_X1 U869 ( .A(n1194), .B(n1195), .Z(G3) );
XNOR2_X1 U870 ( .A(G101), .B(KEYINPUT29), .ZN(n1195) );
NAND2_X1 U871 ( .A1(KEYINPUT2), .A2(n1083), .ZN(n1194) );
NAND3_X1 U872 ( .A1(n1154), .A2(n1034), .A3(n1015), .ZN(n1083) );
XOR2_X1 U873 ( .A(n1196), .B(G125), .Z(G27) );
NAND2_X1 U874 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U875 ( .A1(n1167), .A2(n1199), .ZN(n1198) );
INV_X1 U876 ( .A(KEYINPUT1), .ZN(n1199) );
NOR2_X1 U877 ( .A1(n1200), .A2(n1030), .ZN(n1167) );
NAND3_X1 U878 ( .A1(n1156), .A2(n1200), .A3(KEYINPUT1), .ZN(n1197) );
NAND4_X1 U879 ( .A1(n1028), .A2(n1017), .A3(n1020), .A4(n1181), .ZN(n1200) );
NAND2_X1 U880 ( .A1(n1008), .A2(n1201), .ZN(n1181) );
NAND4_X1 U881 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1061), .ZN(n1201) );
INV_X1 U882 ( .A(G900), .ZN(n1061) );
XOR2_X1 U883 ( .A(n1203), .B(n1147), .Z(G24) );
NAND4_X1 U884 ( .A1(n1204), .A2(n1153), .A3(n1177), .A4(n1178), .ZN(n1147) );
INV_X1 U885 ( .A(n1019), .ZN(n1153) );
NAND2_X1 U886 ( .A1(n1205), .A2(n1206), .ZN(n1019) );
INV_X1 U887 ( .A(n1207), .ZN(n1206) );
XOR2_X1 U888 ( .A(G119), .B(n1208), .Z(G21) );
NOR2_X1 U889 ( .A1(n1030), .A2(n1157), .ZN(n1208) );
NAND3_X1 U890 ( .A1(n1028), .A2(n1034), .A3(n1209), .ZN(n1157) );
NOR3_X1 U891 ( .A1(n1205), .A2(n1210), .A3(n1193), .ZN(n1209) );
INV_X1 U892 ( .A(n1010), .ZN(n1028) );
XNOR2_X1 U893 ( .A(G116), .B(n1152), .ZN(G18) );
NAND3_X1 U894 ( .A1(n1015), .A2(n1021), .A3(n1204), .ZN(n1152) );
XNOR2_X1 U895 ( .A(G113), .B(n1151), .ZN(G15) );
NAND3_X1 U896 ( .A1(n1015), .A2(n1020), .A3(n1204), .ZN(n1151) );
NOR3_X1 U897 ( .A1(n1030), .A2(n1210), .A3(n1010), .ZN(n1204) );
NAND2_X1 U898 ( .A1(n1007), .A2(n1211), .ZN(n1010) );
AND2_X1 U899 ( .A1(n1212), .A2(n1178), .ZN(n1020) );
XOR2_X1 U900 ( .A(KEYINPUT46), .B(n1213), .Z(n1212) );
NOR2_X1 U901 ( .A1(n1056), .A2(n1193), .ZN(n1015) );
XNOR2_X1 U902 ( .A(G110), .B(n1150), .ZN(G12) );
NAND3_X1 U903 ( .A1(n1154), .A2(n1034), .A3(n1017), .ZN(n1150) );
AND2_X1 U904 ( .A1(n1214), .A2(n1056), .ZN(n1017) );
INV_X1 U905 ( .A(n1205), .ZN(n1056) );
XOR2_X1 U906 ( .A(n1215), .B(n1093), .Z(n1205) );
AND2_X1 U907 ( .A1(G217), .A2(n1216), .ZN(n1093) );
NAND2_X1 U908 ( .A1(n1091), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U909 ( .A(n1218), .B(n1219), .ZN(n1091) );
XOR2_X1 U910 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U911 ( .A(n1222), .B(G110), .Z(n1221) );
NAND2_X1 U912 ( .A1(KEYINPUT32), .A2(n1223), .ZN(n1222) );
XOR2_X1 U913 ( .A(G146), .B(n1070), .Z(n1223) );
XNOR2_X1 U914 ( .A(G125), .B(n1179), .ZN(n1070) );
NAND2_X1 U915 ( .A1(n1224), .A2(G221), .ZN(n1220) );
XNOR2_X1 U916 ( .A(G119), .B(n1225), .ZN(n1218) );
XOR2_X1 U917 ( .A(G137), .B(G128), .Z(n1225) );
XOR2_X1 U918 ( .A(n1207), .B(KEYINPUT27), .Z(n1214) );
XOR2_X1 U919 ( .A(n1193), .B(KEYINPUT16), .Z(n1207) );
XOR2_X1 U920 ( .A(n1226), .B(n1227), .Z(n1193) );
XOR2_X1 U921 ( .A(KEYINPUT30), .B(G472), .Z(n1227) );
NAND2_X1 U922 ( .A1(n1228), .A2(n1217), .ZN(n1226) );
XOR2_X1 U923 ( .A(n1117), .B(n1229), .Z(n1228) );
XNOR2_X1 U924 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U925 ( .A1(KEYINPUT4), .A2(n1118), .ZN(n1231) );
NAND3_X1 U926 ( .A1(n1232), .A2(n1023), .A3(G210), .ZN(n1118) );
NAND2_X1 U927 ( .A1(KEYINPUT17), .A2(n1071), .ZN(n1230) );
XOR2_X1 U928 ( .A(n1233), .B(n1234), .Z(n1117) );
XOR2_X1 U929 ( .A(n1235), .B(KEYINPUT28), .Z(n1233) );
NAND2_X1 U930 ( .A1(n1236), .A2(n1237), .ZN(n1034) );
OR3_X1 U931 ( .A1(n1177), .A2(n1178), .A3(KEYINPUT46), .ZN(n1237) );
NAND2_X1 U932 ( .A1(KEYINPUT46), .A2(n1021), .ZN(n1236) );
NOR2_X1 U933 ( .A1(n1178), .A2(n1213), .ZN(n1021) );
INV_X1 U934 ( .A(n1177), .ZN(n1213) );
NAND2_X1 U935 ( .A1(n1238), .A2(n1037), .ZN(n1177) );
NAND2_X1 U936 ( .A1(n1239), .A2(n1240), .ZN(n1037) );
XNOR2_X1 U937 ( .A(n1055), .B(KEYINPUT57), .ZN(n1238) );
NOR2_X1 U938 ( .A1(n1240), .A2(n1239), .ZN(n1055) );
XNOR2_X1 U939 ( .A(G478), .B(KEYINPUT24), .ZN(n1239) );
NAND2_X1 U940 ( .A1(n1241), .A2(n1217), .ZN(n1240) );
XOR2_X1 U941 ( .A(n1096), .B(KEYINPUT31), .Z(n1241) );
XOR2_X1 U942 ( .A(n1242), .B(n1243), .Z(n1096) );
XOR2_X1 U943 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U944 ( .A1(G217), .A2(n1224), .ZN(n1245) );
AND2_X1 U945 ( .A1(G234), .A2(n1023), .ZN(n1224) );
NAND2_X1 U946 ( .A1(KEYINPUT3), .A2(n1246), .ZN(n1244) );
XOR2_X1 U947 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U948 ( .A(G122), .B(G116), .Z(n1248) );
NOR2_X1 U949 ( .A1(G107), .A2(KEYINPUT11), .ZN(n1247) );
XNOR2_X1 U950 ( .A(n1249), .B(n1250), .ZN(n1242) );
NAND2_X1 U951 ( .A1(n1251), .A2(n1252), .ZN(n1178) );
NAND2_X1 U952 ( .A1(G475), .A2(n1253), .ZN(n1252) );
OR2_X1 U953 ( .A1(n1051), .A2(G902), .ZN(n1253) );
XNOR2_X1 U954 ( .A(n1047), .B(KEYINPUT9), .ZN(n1251) );
NOR3_X1 U955 ( .A1(G475), .A2(G902), .A3(n1051), .ZN(n1047) );
XOR2_X1 U956 ( .A(n1254), .B(n1255), .Z(n1051) );
XOR2_X1 U957 ( .A(n1256), .B(n1257), .Z(n1255) );
XNOR2_X1 U958 ( .A(n1258), .B(n1259), .ZN(n1257) );
NAND2_X1 U959 ( .A1(KEYINPUT38), .A2(n1179), .ZN(n1259) );
NAND2_X1 U960 ( .A1(KEYINPUT13), .A2(n1260), .ZN(n1258) );
XOR2_X1 U961 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U962 ( .A(G131), .B(G143), .ZN(n1262) );
NAND3_X1 U963 ( .A1(G214), .A2(n1023), .A3(n1263), .ZN(n1261) );
XOR2_X1 U964 ( .A(n1232), .B(KEYINPUT51), .Z(n1263) );
NAND2_X1 U965 ( .A1(KEYINPUT53), .A2(n1264), .ZN(n1256) );
INV_X1 U966 ( .A(G104), .ZN(n1264) );
XOR2_X1 U967 ( .A(n1265), .B(n1266), .Z(n1254) );
NOR2_X1 U968 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U969 ( .A(KEYINPUT20), .B(n1269), .Z(n1268) );
AND2_X1 U970 ( .A1(n1203), .A2(G113), .ZN(n1269) );
NOR2_X1 U971 ( .A1(G113), .A2(n1203), .ZN(n1267) );
XNOR2_X1 U972 ( .A(G125), .B(n1270), .ZN(n1265) );
NOR2_X1 U973 ( .A1(KEYINPUT48), .A2(n1271), .ZN(n1270) );
XOR2_X1 U974 ( .A(n1173), .B(KEYINPUT12), .Z(n1271) );
NOR3_X1 U975 ( .A1(n1030), .A2(n1210), .A3(n1190), .ZN(n1154) );
INV_X1 U976 ( .A(n1192), .ZN(n1190) );
NOR2_X1 U977 ( .A1(n1007), .A2(n1005), .ZN(n1192) );
INV_X1 U978 ( .A(n1211), .ZN(n1005) );
NAND2_X1 U979 ( .A1(G221), .A2(n1216), .ZN(n1211) );
NAND2_X1 U980 ( .A1(G234), .A2(n1217), .ZN(n1216) );
XOR2_X1 U981 ( .A(n1045), .B(n1272), .Z(n1007) );
NOR2_X1 U982 ( .A1(KEYINPUT40), .A2(n1044), .ZN(n1272) );
INV_X1 U983 ( .A(G469), .ZN(n1044) );
NAND2_X1 U984 ( .A1(n1273), .A2(n1217), .ZN(n1045) );
XOR2_X1 U985 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U986 ( .A(n1276), .B(n1131), .Z(n1275) );
XOR2_X1 U987 ( .A(G110), .B(n1179), .Z(n1131) );
INV_X1 U988 ( .A(G140), .ZN(n1179) );
NAND3_X1 U989 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1276) );
NAND2_X1 U990 ( .A1(n1067), .A2(n1280), .ZN(n1279) );
NAND2_X1 U991 ( .A1(n1281), .A2(KEYINPUT52), .ZN(n1280) );
XNOR2_X1 U992 ( .A(n1138), .B(KEYINPUT54), .ZN(n1281) );
NAND3_X1 U993 ( .A1(KEYINPUT52), .A2(n1282), .A3(n1138), .ZN(n1278) );
INV_X1 U994 ( .A(n1067), .ZN(n1282) );
NAND2_X1 U995 ( .A1(n1283), .A2(n1284), .ZN(n1067) );
NAND2_X1 U996 ( .A1(n1250), .A2(n1173), .ZN(n1284) );
NAND2_X1 U997 ( .A1(n1285), .A2(G146), .ZN(n1283) );
XOR2_X1 U998 ( .A(KEYINPUT25), .B(n1250), .Z(n1285) );
OR2_X1 U999 ( .A1(n1138), .A2(KEYINPUT52), .ZN(n1277) );
XOR2_X1 U1000 ( .A(n1286), .B(n1287), .Z(n1138) );
NOR2_X1 U1001 ( .A1(G101), .A2(KEYINPUT58), .ZN(n1287) );
XOR2_X1 U1002 ( .A(n1134), .B(n1288), .Z(n1274) );
NOR2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1071), .ZN(n1288) );
XOR2_X1 U1004 ( .A(n1289), .B(n1249), .Z(n1071) );
XOR2_X1 U1005 ( .A(G134), .B(KEYINPUT7), .Z(n1249) );
XNOR2_X1 U1006 ( .A(G131), .B(G137), .ZN(n1289) );
NOR2_X1 U1007 ( .A1(n1060), .A2(G953), .ZN(n1134) );
INV_X1 U1008 ( .A(G227), .ZN(n1060) );
AND2_X1 U1009 ( .A1(n1008), .A2(n1290), .ZN(n1210) );
NAND4_X1 U1010 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1086), .ZN(n1290) );
INV_X1 U1011 ( .A(G898), .ZN(n1086) );
NAND3_X1 U1012 ( .A1(n1202), .A2(n1023), .A3(G952), .ZN(n1008) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1202) );
INV_X1 U1014 ( .A(n1156), .ZN(n1030) );
NOR2_X1 U1015 ( .A1(n1033), .A2(n1032), .ZN(n1156) );
INV_X1 U1016 ( .A(n1189), .ZN(n1032) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1291), .ZN(n1189) );
XNOR2_X1 U1018 ( .A(n1054), .B(n1145), .ZN(n1033) );
INV_X1 U1019 ( .A(n1052), .ZN(n1145) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1291), .ZN(n1052) );
NAND2_X1 U1021 ( .A1(n1232), .A2(n1217), .ZN(n1291) );
INV_X1 U1022 ( .A(G237), .ZN(n1232) );
AND2_X1 U1023 ( .A1(n1292), .A2(n1217), .ZN(n1054) );
INV_X1 U1024 ( .A(G902), .ZN(n1217) );
XNOR2_X1 U1025 ( .A(n1141), .B(n1293), .ZN(n1292) );
XOR2_X1 U1026 ( .A(n1294), .B(KEYINPUT5), .Z(n1293) );
NAND2_X1 U1027 ( .A1(n1171), .A2(n1170), .ZN(n1294) );
NAND3_X1 U1028 ( .A1(G224), .A2(n1023), .A3(n1295), .ZN(n1170) );
XOR2_X1 U1029 ( .A(n1235), .B(G125), .Z(n1295) );
NAND2_X1 U1030 ( .A1(n1296), .A2(n1297), .ZN(n1171) );
NAND2_X1 U1031 ( .A1(G224), .A2(n1023), .ZN(n1297) );
INV_X1 U1032 ( .A(G953), .ZN(n1023) );
XOR2_X1 U1033 ( .A(G125), .B(n1298), .Z(n1296) );
INV_X1 U1034 ( .A(n1235), .ZN(n1298) );
XOR2_X1 U1035 ( .A(n1173), .B(n1250), .Z(n1235) );
XOR2_X1 U1036 ( .A(G128), .B(G143), .Z(n1250) );
INV_X1 U1037 ( .A(G146), .ZN(n1173) );
XNOR2_X1 U1038 ( .A(n1084), .B(KEYINPUT47), .ZN(n1141) );
XOR2_X1 U1039 ( .A(n1299), .B(n1300), .Z(n1084) );
XOR2_X1 U1040 ( .A(n1203), .B(n1301), .Z(n1300) );
XNOR2_X1 U1041 ( .A(KEYINPUT23), .B(KEYINPUT10), .ZN(n1301) );
INV_X1 U1042 ( .A(G122), .ZN(n1203) );
XOR2_X1 U1043 ( .A(n1302), .B(n1286), .Z(n1299) );
XOR2_X1 U1044 ( .A(G107), .B(G104), .Z(n1286) );
XNOR2_X1 U1045 ( .A(G110), .B(n1234), .ZN(n1302) );
XNOR2_X1 U1046 ( .A(n1303), .B(n1304), .ZN(n1234) );
XOR2_X1 U1047 ( .A(G119), .B(G116), .Z(n1304) );
XNOR2_X1 U1048 ( .A(G101), .B(G113), .ZN(n1303) );
endmodule


