//Key = 0010111010010100000101011110100101011000100110110001000010100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393;

XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(G9) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(G75) );
NOR4_X1 U773 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
XOR2_X1 U774 ( .A(n1080), .B(KEYINPUT37), .Z(n1079) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND4_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
OR2_X1 U778 ( .A1(n1087), .A2(n1089), .ZN(n1085) );
NAND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND3_X1 U781 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NAND3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1092) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1078) );
INV_X1 U784 ( .A(n1090), .ZN(n1101) );
NOR3_X1 U785 ( .A1(n1102), .A2(n1088), .A3(n1103), .ZN(n1090) );
INV_X1 U786 ( .A(n1104), .ZN(n1088) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
AND2_X1 U789 ( .A1(n1096), .A2(n1109), .ZN(n1105) );
NAND3_X1 U790 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1076) );
NAND2_X1 U791 ( .A1(n1084), .A2(n1113), .ZN(n1112) );
NAND2_X1 U792 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1118), .ZN(n1114) );
NOR3_X1 U795 ( .A1(n1119), .A2(n1108), .A3(n1103), .ZN(n1084) );
INV_X1 U796 ( .A(n1098), .ZN(n1108) );
AND3_X1 U797 ( .A1(n1110), .A2(n1111), .A3(n1120), .ZN(n1074) );
NAND4_X1 U798 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1110) );
NOR4_X1 U799 ( .A1(n1087), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1124) );
XNOR2_X1 U800 ( .A(n1128), .B(n1129), .ZN(n1126) );
NAND2_X1 U801 ( .A1(KEYINPUT28), .A2(n1130), .ZN(n1128) );
INV_X1 U802 ( .A(n1131), .ZN(n1125) );
NOR2_X1 U803 ( .A1(n1119), .A2(n1132), .ZN(n1123) );
XNOR2_X1 U804 ( .A(KEYINPUT20), .B(n1133), .ZN(n1132) );
XOR2_X1 U805 ( .A(n1134), .B(G469), .Z(n1122) );
XOR2_X1 U806 ( .A(n1135), .B(n1136), .Z(n1121) );
XOR2_X1 U807 ( .A(n1137), .B(n1138), .Z(G72) );
NAND2_X1 U808 ( .A1(G953), .A2(n1139), .ZN(n1138) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1139) );
NAND2_X1 U810 ( .A1(n1140), .A2(KEYINPUT5), .ZN(n1137) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U812 ( .A1(KEYINPUT22), .A2(n1143), .ZN(n1142) );
NOR2_X1 U813 ( .A1(n1144), .A2(G953), .ZN(n1143) );
NAND2_X1 U814 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
NAND2_X1 U815 ( .A1(G953), .A2(n1147), .ZN(n1146) );
XOR2_X1 U816 ( .A(n1148), .B(n1149), .Z(n1145) );
XOR2_X1 U817 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR3_X1 U818 ( .A1(KEYINPUT48), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR3_X1 U819 ( .A1(G131), .A2(n1154), .A3(n1155), .ZN(n1153) );
NOR2_X1 U820 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1156) );
XOR2_X1 U822 ( .A(n1158), .B(KEYINPUT2), .Z(n1155) );
NAND2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U824 ( .A1(n1159), .A2(n1160), .ZN(n1154) );
INV_X1 U825 ( .A(G134), .ZN(n1160) );
XOR2_X1 U826 ( .A(n1161), .B(n1162), .Z(G69) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U828 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U829 ( .A(KEYINPUT59), .B(G953), .Z(n1166) );
NAND2_X1 U830 ( .A1(n1167), .A2(n1168), .ZN(n1163) );
NAND2_X1 U831 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U832 ( .A(KEYINPUT52), .B(G953), .Z(n1169) );
XOR2_X1 U833 ( .A(KEYINPUT35), .B(n1171), .Z(n1167) );
NAND2_X1 U834 ( .A1(G953), .A2(n1172), .ZN(n1161) );
NAND2_X1 U835 ( .A1(G898), .A2(G224), .ZN(n1172) );
NOR2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND4_X1 U838 ( .A1(n1177), .A2(G217), .A3(n1077), .A4(n1178), .ZN(n1175) );
XOR2_X1 U839 ( .A(n1179), .B(KEYINPUT26), .Z(n1177) );
NOR3_X1 U840 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G63) );
AND2_X1 U841 ( .A1(KEYINPUT51), .A2(n1173), .ZN(n1182) );
NOR3_X1 U842 ( .A1(KEYINPUT51), .A2(n1111), .A3(n1120), .ZN(n1181) );
INV_X1 U843 ( .A(G952), .ZN(n1120) );
NOR3_X1 U844 ( .A1(n1135), .A2(n1183), .A3(n1184), .ZN(n1180) );
AND3_X1 U845 ( .A1(n1185), .A2(G478), .A3(n1186), .ZN(n1184) );
NOR2_X1 U846 ( .A1(n1185), .A2(n1187), .ZN(n1183) );
AND2_X1 U847 ( .A1(n1077), .A2(G478), .ZN(n1187) );
NOR2_X1 U848 ( .A1(n1173), .A2(n1188), .ZN(G60) );
XOR2_X1 U849 ( .A(n1189), .B(n1190), .Z(n1188) );
AND2_X1 U850 ( .A1(G475), .A2(n1186), .ZN(n1190) );
XNOR2_X1 U851 ( .A(G104), .B(n1191), .ZN(G6) );
NOR3_X1 U852 ( .A1(n1173), .A2(n1192), .A3(n1193), .ZN(G57) );
NOR2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U854 ( .A(KEYINPUT54), .B(n1196), .ZN(n1194) );
NOR2_X1 U855 ( .A1(n1197), .A2(n1196), .ZN(n1192) );
NAND2_X1 U856 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
OR2_X1 U857 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U858 ( .A(n1202), .B(KEYINPUT15), .Z(n1198) );
NAND2_X1 U859 ( .A1(n1201), .A2(n1200), .ZN(n1202) );
XNOR2_X1 U860 ( .A(n1203), .B(n1204), .ZN(n1200) );
XOR2_X1 U861 ( .A(n1205), .B(n1206), .Z(n1203) );
NAND2_X1 U862 ( .A1(KEYINPUT44), .A2(n1207), .ZN(n1205) );
NOR2_X1 U863 ( .A1(n1208), .A2(n1130), .ZN(n1201) );
INV_X1 U864 ( .A(G472), .ZN(n1130) );
INV_X1 U865 ( .A(n1195), .ZN(n1197) );
XOR2_X1 U866 ( .A(n1209), .B(n1210), .Z(n1195) );
NAND2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
XNOR2_X1 U868 ( .A(KEYINPUT39), .B(KEYINPUT17), .ZN(n1211) );
NOR3_X1 U869 ( .A1(n1173), .A2(n1213), .A3(n1214), .ZN(G54) );
NOR2_X1 U870 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U871 ( .A(n1217), .B(n1218), .Z(n1215) );
NOR2_X1 U872 ( .A1(KEYINPUT45), .A2(n1219), .ZN(n1218) );
INV_X1 U873 ( .A(n1220), .ZN(n1219) );
NOR2_X1 U874 ( .A1(n1221), .A2(n1222), .ZN(n1213) );
XOR2_X1 U875 ( .A(n1217), .B(n1223), .Z(n1222) );
NOR2_X1 U876 ( .A1(KEYINPUT45), .A2(n1220), .ZN(n1223) );
XOR2_X1 U877 ( .A(n1224), .B(n1225), .Z(n1220) );
NOR2_X1 U878 ( .A1(KEYINPUT50), .A2(n1226), .ZN(n1225) );
XOR2_X1 U879 ( .A(n1227), .B(KEYINPUT49), .Z(n1226) );
AND2_X1 U880 ( .A1(n1186), .A2(G469), .ZN(n1217) );
INV_X1 U881 ( .A(n1216), .ZN(n1221) );
NAND3_X1 U882 ( .A1(n1228), .A2(n1229), .A3(KEYINPUT56), .ZN(n1216) );
NAND2_X1 U883 ( .A1(G110), .A2(n1230), .ZN(n1229) );
NAND2_X1 U884 ( .A1(n1231), .A2(n1232), .ZN(n1228) );
XOR2_X1 U885 ( .A(n1230), .B(KEYINPUT19), .Z(n1231) );
NOR2_X1 U886 ( .A1(n1173), .A2(n1233), .ZN(G51) );
NOR3_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NOR2_X1 U888 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U889 ( .A(n1239), .B(n1240), .ZN(n1237) );
NOR3_X1 U890 ( .A1(G125), .A2(n1239), .A3(n1240), .ZN(n1235) );
AND2_X1 U891 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
XOR2_X1 U892 ( .A(n1242), .B(n1243), .Z(n1240) );
NAND3_X1 U893 ( .A1(n1186), .A2(n1244), .A3(KEYINPUT6), .ZN(n1242) );
INV_X1 U894 ( .A(n1208), .ZN(n1186) );
NAND2_X1 U895 ( .A1(G902), .A2(n1077), .ZN(n1208) );
NAND2_X1 U896 ( .A1(n1165), .A2(n1144), .ZN(n1077) );
AND2_X1 U897 ( .A1(n1245), .A2(n1246), .ZN(n1144) );
NOR4_X1 U898 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
INV_X1 U899 ( .A(n1251), .ZN(n1250) );
INV_X1 U900 ( .A(n1252), .ZN(n1249) );
NOR4_X1 U901 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1245) );
NOR2_X1 U902 ( .A1(n1107), .A2(n1257), .ZN(n1256) );
INV_X1 U903 ( .A(n1258), .ZN(n1255) );
NOR2_X1 U904 ( .A1(n1119), .A2(n1259), .ZN(n1253) );
AND2_X1 U905 ( .A1(n1260), .A2(n1261), .ZN(n1165) );
AND4_X1 U906 ( .A1(n1262), .A2(n1191), .A3(n1073), .A4(n1263), .ZN(n1261) );
NAND3_X1 U907 ( .A1(n1089), .A2(n1098), .A3(n1264), .ZN(n1073) );
NAND3_X1 U908 ( .A1(n1264), .A2(n1098), .A3(n1117), .ZN(n1191) );
AND4_X1 U909 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1260) );
OR2_X1 U910 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U911 ( .A(n1107), .B(KEYINPUT3), .Z(n1269) );
NOR2_X1 U912 ( .A1(n1111), .A2(G952), .ZN(n1173) );
XOR2_X1 U913 ( .A(n1271), .B(n1272), .Z(G48) );
NAND2_X1 U914 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U915 ( .A(KEYINPUT27), .B(n1257), .ZN(n1274) );
NAND2_X1 U916 ( .A1(n1275), .A2(n1117), .ZN(n1257) );
XOR2_X1 U917 ( .A(n1276), .B(n1252), .Z(G45) );
NAND4_X1 U918 ( .A1(n1277), .A2(n1278), .A3(n1273), .A4(n1127), .ZN(n1252) );
XOR2_X1 U919 ( .A(n1279), .B(n1258), .Z(G42) );
NAND3_X1 U920 ( .A1(n1096), .A2(n1118), .A3(n1280), .ZN(n1258) );
XOR2_X1 U921 ( .A(G137), .B(n1248), .Z(G39) );
AND3_X1 U922 ( .A1(n1104), .A2(n1096), .A3(n1275), .ZN(n1248) );
XOR2_X1 U923 ( .A(G134), .B(n1281), .Z(G36) );
NOR3_X1 U924 ( .A1(n1119), .A2(KEYINPUT7), .A3(n1282), .ZN(n1281) );
XOR2_X1 U925 ( .A(n1259), .B(KEYINPUT55), .Z(n1282) );
NAND2_X1 U926 ( .A1(n1278), .A2(n1089), .ZN(n1259) );
XOR2_X1 U927 ( .A(G131), .B(n1254), .Z(G33) );
AND3_X1 U928 ( .A1(n1117), .A2(n1096), .A3(n1278), .ZN(n1254) );
AND3_X1 U929 ( .A1(n1118), .A2(n1283), .A3(n1109), .ZN(n1278) );
INV_X1 U930 ( .A(n1119), .ZN(n1096) );
NAND2_X1 U931 ( .A1(n1097), .A2(n1284), .ZN(n1119) );
XOR2_X1 U932 ( .A(G128), .B(n1247), .Z(G30) );
AND3_X1 U933 ( .A1(n1089), .A2(n1273), .A3(n1275), .ZN(n1247) );
AND4_X1 U934 ( .A1(n1118), .A2(n1285), .A3(n1283), .A4(n1095), .ZN(n1275) );
XNOR2_X1 U935 ( .A(n1262), .B(n1286), .ZN(G3) );
NOR2_X1 U936 ( .A1(KEYINPUT1), .A2(n1212), .ZN(n1286) );
NAND3_X1 U937 ( .A1(n1109), .A2(n1264), .A3(n1104), .ZN(n1262) );
XOR2_X1 U938 ( .A(n1238), .B(n1251), .Z(G27) );
NAND3_X1 U939 ( .A1(n1116), .A2(n1273), .A3(n1280), .ZN(n1251) );
AND4_X1 U940 ( .A1(n1094), .A2(n1117), .A3(n1283), .A4(n1095), .ZN(n1280) );
NAND2_X1 U941 ( .A1(n1103), .A2(n1287), .ZN(n1283) );
NAND4_X1 U942 ( .A1(G953), .A2(G902), .A3(n1288), .A4(n1147), .ZN(n1287) );
INV_X1 U943 ( .A(G900), .ZN(n1147) );
NAND2_X1 U944 ( .A1(n1289), .A2(n1290), .ZN(G24) );
NAND2_X1 U945 ( .A1(G122), .A2(n1267), .ZN(n1290) );
XOR2_X1 U946 ( .A(n1291), .B(KEYINPUT61), .Z(n1289) );
OR2_X1 U947 ( .A1(n1267), .A2(G122), .ZN(n1291) );
NAND4_X1 U948 ( .A1(n1292), .A2(n1098), .A3(n1277), .A4(n1127), .ZN(n1267) );
NOR2_X1 U949 ( .A1(n1095), .A2(n1285), .ZN(n1098) );
XNOR2_X1 U950 ( .A(G119), .B(n1266), .ZN(G21) );
NAND4_X1 U951 ( .A1(n1292), .A2(n1104), .A3(n1285), .A4(n1095), .ZN(n1266) );
INV_X1 U952 ( .A(n1094), .ZN(n1285) );
XNOR2_X1 U953 ( .A(G116), .B(n1265), .ZN(G18) );
NAND3_X1 U954 ( .A1(n1109), .A2(n1089), .A3(n1292), .ZN(n1265) );
AND3_X1 U955 ( .A1(n1273), .A2(n1293), .A3(n1116), .ZN(n1292) );
NOR2_X1 U956 ( .A1(n1127), .A2(n1294), .ZN(n1089) );
XOR2_X1 U957 ( .A(G113), .B(n1295), .Z(G15) );
NOR2_X1 U958 ( .A1(n1107), .A2(n1270), .ZN(n1295) );
NAND4_X1 U959 ( .A1(n1116), .A2(n1117), .A3(n1109), .A4(n1293), .ZN(n1270) );
NOR2_X1 U960 ( .A1(n1095), .A2(n1094), .ZN(n1109) );
AND2_X1 U961 ( .A1(n1294), .A2(n1127), .ZN(n1117) );
INV_X1 U962 ( .A(n1277), .ZN(n1294) );
INV_X1 U963 ( .A(n1102), .ZN(n1116) );
NAND2_X1 U964 ( .A1(n1083), .A2(n1296), .ZN(n1102) );
INV_X1 U965 ( .A(n1273), .ZN(n1107) );
XOR2_X1 U966 ( .A(n1232), .B(n1263), .Z(G12) );
NAND4_X1 U967 ( .A1(n1104), .A2(n1264), .A3(n1094), .A4(n1095), .ZN(n1263) );
NAND2_X1 U968 ( .A1(n1131), .A2(n1133), .ZN(n1095) );
NAND3_X1 U969 ( .A1(n1297), .A2(n1179), .A3(n1176), .ZN(n1133) );
NAND2_X1 U970 ( .A1(G217), .A2(n1178), .ZN(n1297) );
NAND3_X1 U971 ( .A1(n1298), .A2(n1178), .A3(G217), .ZN(n1131) );
NAND2_X1 U972 ( .A1(n1176), .A2(n1179), .ZN(n1298) );
XNOR2_X1 U973 ( .A(n1299), .B(n1300), .ZN(n1176) );
XNOR2_X1 U974 ( .A(n1159), .B(n1301), .ZN(n1300) );
XOR2_X1 U975 ( .A(n1302), .B(n1303), .Z(n1301) );
AND3_X1 U976 ( .A1(n1304), .A2(n1111), .A3(G221), .ZN(n1303) );
NAND2_X1 U977 ( .A1(KEYINPUT8), .A2(G128), .ZN(n1302) );
XOR2_X1 U978 ( .A(n1305), .B(n1306), .Z(n1299) );
XOR2_X1 U979 ( .A(G119), .B(G110), .Z(n1306) );
NAND3_X1 U980 ( .A1(n1307), .A2(n1308), .A3(KEYINPUT40), .ZN(n1305) );
NAND2_X1 U981 ( .A1(n1309), .A2(n1271), .ZN(n1308) );
XOR2_X1 U982 ( .A(KEYINPUT47), .B(n1310), .Z(n1307) );
NOR2_X1 U983 ( .A1(n1309), .A2(n1271), .ZN(n1310) );
INV_X1 U984 ( .A(n1151), .ZN(n1309) );
XOR2_X1 U985 ( .A(n1129), .B(G472), .Z(n1094) );
NAND2_X1 U986 ( .A1(n1311), .A2(n1179), .ZN(n1129) );
XOR2_X1 U987 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U988 ( .A(n1212), .B(n1210), .Z(n1313) );
AND3_X1 U989 ( .A1(n1314), .A2(n1111), .A3(G210), .ZN(n1210) );
NAND2_X1 U990 ( .A1(n1315), .A2(n1316), .ZN(n1312) );
NAND2_X1 U991 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U992 ( .A(KEYINPUT24), .B(n1206), .Z(n1318) );
XOR2_X1 U993 ( .A(n1224), .B(n1204), .Z(n1317) );
XOR2_X1 U994 ( .A(n1319), .B(KEYINPUT10), .Z(n1315) );
NAND2_X1 U995 ( .A1(n1320), .A2(n1206), .ZN(n1319) );
XNOR2_X1 U996 ( .A(n1321), .B(n1322), .ZN(n1206) );
XOR2_X1 U997 ( .A(KEYINPUT23), .B(n1323), .Z(n1322) );
XOR2_X1 U998 ( .A(n1204), .B(n1207), .Z(n1320) );
XOR2_X1 U999 ( .A(n1239), .B(KEYINPUT9), .Z(n1204) );
AND3_X1 U1000 ( .A1(n1118), .A2(n1293), .A3(n1273), .ZN(n1264) );
NOR2_X1 U1001 ( .A1(n1097), .A2(n1099), .ZN(n1273) );
INV_X1 U1002 ( .A(n1284), .ZN(n1099) );
NAND2_X1 U1003 ( .A1(n1324), .A2(n1325), .ZN(n1284) );
XNOR2_X1 U1004 ( .A(G214), .B(KEYINPUT11), .ZN(n1324) );
XOR2_X1 U1005 ( .A(n1326), .B(n1244), .Z(n1097) );
AND2_X1 U1006 ( .A1(G210), .A2(n1325), .ZN(n1244) );
NAND2_X1 U1007 ( .A1(n1327), .A2(n1314), .ZN(n1325) );
NAND2_X1 U1008 ( .A1(n1328), .A2(n1179), .ZN(n1326) );
XNOR2_X1 U1009 ( .A(n1243), .B(n1329), .ZN(n1328) );
NOR3_X1 U1010 ( .A1(n1330), .A2(KEYINPUT12), .A3(n1241), .ZN(n1329) );
AND2_X1 U1011 ( .A1(n1239), .A2(n1238), .ZN(n1241) );
XOR2_X1 U1012 ( .A(KEYINPUT32), .B(n1331), .Z(n1330) );
NOR2_X1 U1013 ( .A1(n1332), .A2(n1239), .ZN(n1331) );
XOR2_X1 U1014 ( .A(G146), .B(n1333), .Z(n1239) );
XOR2_X1 U1015 ( .A(n1238), .B(KEYINPUT30), .Z(n1332) );
INV_X1 U1016 ( .A(G125), .ZN(n1238) );
XNOR2_X1 U1017 ( .A(n1334), .B(n1171), .ZN(n1243) );
XNOR2_X1 U1018 ( .A(n1335), .B(n1336), .ZN(n1171) );
XOR2_X1 U1019 ( .A(G107), .B(n1337), .Z(n1336) );
XOR2_X1 U1020 ( .A(KEYINPUT38), .B(G110), .Z(n1337) );
XNOR2_X1 U1021 ( .A(n1338), .B(n1339), .ZN(n1335) );
XOR2_X1 U1022 ( .A(n1212), .B(n1340), .Z(n1339) );
NAND2_X1 U1023 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1024 ( .A1(n1321), .A2(n1323), .ZN(n1342) );
XOR2_X1 U1025 ( .A(n1343), .B(KEYINPUT14), .Z(n1341) );
OR2_X1 U1026 ( .A1(n1323), .A2(n1321), .ZN(n1343) );
XOR2_X1 U1027 ( .A(G116), .B(G119), .Z(n1323) );
NAND2_X1 U1028 ( .A1(G224), .A2(n1111), .ZN(n1334) );
NAND2_X1 U1029 ( .A1(n1103), .A2(n1344), .ZN(n1293) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1288), .A4(n1170), .ZN(n1344) );
INV_X1 U1031 ( .A(G898), .ZN(n1170) );
NAND3_X1 U1032 ( .A1(n1288), .A2(n1111), .A3(G952), .ZN(n1103) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1288) );
NOR2_X1 U1034 ( .A1(n1083), .A2(n1087), .ZN(n1118) );
INV_X1 U1035 ( .A(n1296), .ZN(n1087) );
NAND2_X1 U1036 ( .A1(G221), .A2(n1178), .ZN(n1296) );
NAND2_X1 U1037 ( .A1(G234), .A2(n1327), .ZN(n1178) );
XOR2_X1 U1038 ( .A(n1179), .B(KEYINPUT62), .Z(n1327) );
XNOR2_X1 U1039 ( .A(n1345), .B(G469), .ZN(n1083) );
NAND2_X1 U1040 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND2_X1 U1041 ( .A1(KEYINPUT41), .A2(n1134), .ZN(n1347) );
NAND2_X1 U1042 ( .A1(KEYINPUT31), .A2(n1348), .ZN(n1346) );
INV_X1 U1043 ( .A(n1134), .ZN(n1348) );
NAND2_X1 U1044 ( .A1(n1349), .A2(n1179), .ZN(n1134) );
INV_X1 U1045 ( .A(G902), .ZN(n1179) );
XOR2_X1 U1046 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1047 ( .A(n1230), .B(n1227), .Z(n1351) );
XOR2_X1 U1048 ( .A(n1148), .B(n1352), .Z(n1227) );
XOR2_X1 U1049 ( .A(n1212), .B(n1353), .Z(n1352) );
NAND2_X1 U1050 ( .A1(n1354), .A2(KEYINPUT46), .ZN(n1353) );
XOR2_X1 U1051 ( .A(G104), .B(n1072), .Z(n1354) );
INV_X1 U1052 ( .A(G107), .ZN(n1072) );
INV_X1 U1053 ( .A(G101), .ZN(n1212) );
NAND2_X1 U1054 ( .A1(n1355), .A2(n1356), .ZN(n1148) );
NAND2_X1 U1055 ( .A1(n1333), .A2(G146), .ZN(n1356) );
NAND2_X1 U1056 ( .A1(n1357), .A2(n1271), .ZN(n1355) );
INV_X1 U1057 ( .A(G146), .ZN(n1271) );
XNOR2_X1 U1058 ( .A(n1333), .B(KEYINPUT42), .ZN(n1357) );
XOR2_X1 U1059 ( .A(n1358), .B(G140), .Z(n1230) );
NAND2_X1 U1060 ( .A1(n1359), .A2(n1111), .ZN(n1358) );
XNOR2_X1 U1061 ( .A(G227), .B(KEYINPUT36), .ZN(n1359) );
XOR2_X1 U1062 ( .A(n1207), .B(n1360), .Z(n1350) );
XOR2_X1 U1063 ( .A(KEYINPUT58), .B(G110), .Z(n1360) );
INV_X1 U1064 ( .A(n1224), .ZN(n1207) );
XOR2_X1 U1065 ( .A(n1361), .B(n1362), .Z(n1224) );
XOR2_X1 U1066 ( .A(G131), .B(n1159), .Z(n1362) );
XOR2_X1 U1067 ( .A(G137), .B(KEYINPUT16), .Z(n1159) );
XOR2_X1 U1068 ( .A(n1363), .B(G134), .Z(n1361) );
XNOR2_X1 U1069 ( .A(KEYINPUT60), .B(KEYINPUT18), .ZN(n1363) );
NOR2_X1 U1070 ( .A1(n1127), .A2(n1277), .ZN(n1104) );
XOR2_X1 U1071 ( .A(n1364), .B(n1135), .Z(n1277) );
NOR2_X1 U1072 ( .A1(n1185), .A2(G902), .ZN(n1135) );
AND2_X1 U1073 ( .A1(n1365), .A2(n1366), .ZN(n1185) );
NAND2_X1 U1074 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND3_X1 U1075 ( .A1(n1304), .A2(n1111), .A3(G217), .ZN(n1368) );
XOR2_X1 U1076 ( .A(n1369), .B(KEYINPUT25), .Z(n1367) );
XOR2_X1 U1077 ( .A(n1370), .B(KEYINPUT0), .Z(n1365) );
NAND4_X1 U1078 ( .A1(n1369), .A2(G217), .A3(n1304), .A4(n1111), .ZN(n1370) );
XNOR2_X1 U1079 ( .A(G234), .B(KEYINPUT4), .ZN(n1304) );
XOR2_X1 U1080 ( .A(n1371), .B(n1372), .Z(n1369) );
NOR2_X1 U1081 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1082 ( .A(KEYINPUT34), .B(n1375), .Z(n1374) );
NOR2_X1 U1083 ( .A1(G107), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1084 ( .A(KEYINPUT53), .B(n1377), .Z(n1376) );
AND2_X1 U1085 ( .A1(n1377), .A2(G107), .ZN(n1373) );
XOR2_X1 U1086 ( .A(G116), .B(G122), .Z(n1377) );
NAND2_X1 U1087 ( .A1(KEYINPUT33), .A2(n1378), .ZN(n1371) );
XOR2_X1 U1088 ( .A(G134), .B(n1333), .Z(n1378) );
XOR2_X1 U1089 ( .A(G128), .B(G143), .Z(n1333) );
NAND2_X1 U1090 ( .A1(KEYINPUT43), .A2(n1136), .ZN(n1364) );
XNOR2_X1 U1091 ( .A(G478), .B(KEYINPUT29), .ZN(n1136) );
XOR2_X1 U1092 ( .A(G475), .B(n1379), .Z(n1127) );
NOR2_X1 U1093 ( .A1(G902), .A2(n1189), .ZN(n1379) );
XOR2_X1 U1094 ( .A(n1380), .B(n1381), .Z(n1189) );
XNOR2_X1 U1095 ( .A(n1321), .B(n1338), .ZN(n1381) );
XOR2_X1 U1096 ( .A(G104), .B(G122), .Z(n1338) );
XNOR2_X1 U1097 ( .A(G113), .B(KEYINPUT63), .ZN(n1321) );
XOR2_X1 U1098 ( .A(n1382), .B(n1383), .Z(n1380) );
NOR2_X1 U1099 ( .A1(KEYINPUT57), .A2(n1384), .ZN(n1383) );
XOR2_X1 U1100 ( .A(G146), .B(n1151), .Z(n1384) );
XNOR2_X1 U1101 ( .A(n1279), .B(G125), .ZN(n1151) );
INV_X1 U1102 ( .A(G140), .ZN(n1279) );
NAND2_X1 U1103 ( .A1(n1385), .A2(n1386), .ZN(n1382) );
NAND2_X1 U1104 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
NAND2_X1 U1105 ( .A1(KEYINPUT21), .A2(n1389), .ZN(n1388) );
NAND2_X1 U1106 ( .A1(KEYINPUT13), .A2(n1157), .ZN(n1389) );
INV_X1 U1107 ( .A(G131), .ZN(n1157) );
NAND2_X1 U1108 ( .A1(G131), .A2(n1390), .ZN(n1385) );
NAND2_X1 U1109 ( .A1(KEYINPUT13), .A2(n1391), .ZN(n1390) );
NAND2_X1 U1110 ( .A1(KEYINPUT21), .A2(n1392), .ZN(n1391) );
INV_X1 U1111 ( .A(n1387), .ZN(n1392) );
XOR2_X1 U1112 ( .A(n1276), .B(n1393), .Z(n1387) );
AND3_X1 U1113 ( .A1(G214), .A2(n1111), .A3(n1314), .ZN(n1393) );
INV_X1 U1114 ( .A(G237), .ZN(n1314) );
INV_X1 U1115 ( .A(G953), .ZN(n1111) );
INV_X1 U1116 ( .A(G143), .ZN(n1276) );
INV_X1 U1117 ( .A(G110), .ZN(n1232) );
endmodule


