//Key = 0000000100011010011101101001101000010000010100110101110001001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400;

XOR2_X1 U769 ( .A(n1066), .B(n1067), .Z(G9) );
NOR2_X1 U770 ( .A1(KEYINPUT15), .A2(n1068), .ZN(n1067) );
NOR2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(G75) );
NOR4_X1 U772 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
XNOR2_X1 U773 ( .A(n1075), .B(KEYINPUT16), .ZN(n1073) );
NAND3_X1 U774 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND4_X1 U777 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND3_X1 U781 ( .A1(n1084), .A2(n1093), .A3(n1083), .ZN(n1092) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1096), .ZN(n1091) );
NAND3_X1 U784 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NAND2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U786 ( .A(KEYINPUT13), .B(n1083), .Z(n1101) );
NAND3_X1 U787 ( .A1(n1102), .A2(n1083), .A3(n1103), .ZN(n1098) );
NAND2_X1 U788 ( .A1(n1084), .A2(n1104), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U791 ( .A(n1109), .ZN(n1079) );
NOR3_X1 U792 ( .A1(n1110), .A2(G953), .A3(n1111), .ZN(n1069) );
INV_X1 U793 ( .A(n1076), .ZN(n1111) );
NAND4_X1 U794 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1076) );
NOR4_X1 U795 ( .A1(n1107), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1115) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1116) );
NOR2_X1 U797 ( .A1(n1121), .A2(KEYINPUT48), .ZN(n1120) );
XNOR2_X1 U798 ( .A(G475), .B(KEYINPUT50), .ZN(n1119) );
XNOR2_X1 U799 ( .A(n1122), .B(n1123), .ZN(n1114) );
XOR2_X1 U800 ( .A(KEYINPUT3), .B(KEYINPUT1), .Z(n1123) );
XNOR2_X1 U801 ( .A(n1124), .B(n1125), .ZN(n1113) );
XNOR2_X1 U802 ( .A(n1126), .B(n1127), .ZN(n1112) );
NAND2_X1 U803 ( .A1(KEYINPUT53), .A2(G472), .ZN(n1126) );
XNOR2_X1 U804 ( .A(KEYINPUT45), .B(n1074), .ZN(n1110) );
INV_X1 U805 ( .A(G952), .ZN(n1074) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(G72) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1077), .ZN(n1129) );
AND2_X1 U808 ( .A1(G227), .A2(G900), .ZN(n1130) );
NAND2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
NAND3_X1 U810 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U811 ( .A1(G953), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U812 ( .A(n1075), .B(KEYINPUT46), .ZN(n1133) );
OR3_X1 U813 ( .A1(n1075), .A2(G953), .A3(n1135), .ZN(n1131) );
XOR2_X1 U814 ( .A(n1137), .B(n1138), .Z(n1135) );
XOR2_X1 U815 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U816 ( .A(KEYINPUT6), .B(n1141), .ZN(n1140) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1137) );
NAND2_X1 U818 ( .A1(n1144), .A2(n1145), .ZN(G69) );
NAND2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
OR2_X1 U820 ( .A1(n1077), .A2(G224), .ZN(n1147) );
NAND3_X1 U821 ( .A1(G953), .A2(n1148), .A3(n1149), .ZN(n1144) );
XNOR2_X1 U822 ( .A(n1146), .B(KEYINPUT38), .ZN(n1149) );
XNOR2_X1 U823 ( .A(n1150), .B(n1151), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1152), .A2(G953), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(n1150) );
INV_X1 U827 ( .A(n1157), .ZN(n1156) );
XNOR2_X1 U828 ( .A(n1158), .B(n1159), .ZN(n1155) );
NAND2_X1 U829 ( .A1(KEYINPUT62), .A2(n1160), .ZN(n1158) );
XOR2_X1 U830 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U831 ( .A1(G898), .A2(G224), .ZN(n1148) );
NOR2_X1 U832 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U834 ( .A1(n1125), .A2(n1167), .ZN(n1166) );
NAND2_X1 U835 ( .A1(KEYINPUT14), .A2(n1168), .ZN(n1165) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1169), .ZN(G63) );
NOR2_X1 U837 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U838 ( .A(n1172), .B(KEYINPUT60), .Z(n1171) );
NAND2_X1 U839 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1174), .ZN(n1170) );
AND2_X1 U841 ( .A1(n1175), .A2(G478), .ZN(n1173) );
NOR2_X1 U842 ( .A1(n1163), .A2(n1176), .ZN(G60) );
NOR3_X1 U843 ( .A1(n1121), .A2(n1177), .A3(n1178), .ZN(n1176) );
AND3_X1 U844 ( .A1(n1179), .A2(G475), .A3(n1175), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1180), .A2(n1179), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1183), .A2(n1072), .ZN(n1181) );
INV_X1 U848 ( .A(n1184), .ZN(n1072) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(G6) );
NAND2_X1 U850 ( .A1(KEYINPUT7), .A2(G104), .ZN(n1186) );
NOR4_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1163), .A4(n1189), .ZN(G57) );
NOR2_X1 U852 ( .A1(G101), .A2(n1190), .ZN(n1189) );
XOR2_X1 U853 ( .A(n1191), .B(n1192), .Z(n1190) );
AND2_X1 U854 ( .A1(n1193), .A2(KEYINPUT43), .ZN(n1191) );
AND3_X1 U855 ( .A1(n1192), .A2(n1194), .A3(KEYINPUT43), .ZN(n1188) );
NOR3_X1 U856 ( .A1(n1192), .A2(n1195), .A3(n1196), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1193), .A2(n1197), .ZN(n1195) );
INV_X1 U858 ( .A(KEYINPUT43), .ZN(n1197) );
XNOR2_X1 U859 ( .A(n1198), .B(n1199), .ZN(n1192) );
XOR2_X1 U860 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U861 ( .A1(KEYINPUT11), .A2(n1202), .ZN(n1201) );
NAND2_X1 U862 ( .A1(n1175), .A2(G472), .ZN(n1200) );
NOR2_X1 U863 ( .A1(n1163), .A2(n1203), .ZN(G54) );
XOR2_X1 U864 ( .A(n1204), .B(n1205), .Z(n1203) );
XNOR2_X1 U865 ( .A(n1206), .B(n1207), .ZN(n1205) );
XNOR2_X1 U866 ( .A(n1208), .B(n1209), .ZN(n1204) );
NAND2_X1 U867 ( .A1(n1175), .A2(G469), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1163), .A2(n1210), .ZN(G51) );
XOR2_X1 U869 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U870 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U871 ( .A(KEYINPUT56), .B(KEYINPUT21), .Z(n1214) );
XOR2_X1 U872 ( .A(n1215), .B(n1216), .Z(n1211) );
XNOR2_X1 U873 ( .A(n1217), .B(n1218), .ZN(n1215) );
NAND2_X1 U874 ( .A1(n1175), .A2(n1219), .ZN(n1217) );
INV_X1 U875 ( .A(n1167), .ZN(n1175) );
NAND2_X1 U876 ( .A1(G902), .A2(n1220), .ZN(n1167) );
NAND2_X1 U877 ( .A1(n1184), .A2(n1075), .ZN(n1220) );
INV_X1 U878 ( .A(n1183), .ZN(n1075) );
NAND4_X1 U879 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1183) );
NOR4_X1 U880 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
INV_X1 U881 ( .A(n1229), .ZN(n1225) );
NOR2_X1 U882 ( .A1(n1230), .A2(n1231), .ZN(n1223) );
NOR2_X1 U883 ( .A1(KEYINPUT32), .A2(n1232), .ZN(n1231) );
NOR3_X1 U884 ( .A1(n1087), .A2(n1233), .A3(n1234), .ZN(n1230) );
NOR3_X1 U885 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1234) );
AND2_X1 U886 ( .A1(n1238), .A2(KEYINPUT58), .ZN(n1237) );
AND3_X1 U887 ( .A1(KEYINPUT32), .A2(n1084), .A3(n1239), .ZN(n1236) );
NOR2_X1 U888 ( .A1(n1240), .A2(n1094), .ZN(n1233) );
NOR2_X1 U889 ( .A1(KEYINPUT58), .A2(n1241), .ZN(n1240) );
NOR2_X1 U890 ( .A1(n1242), .A2(n1154), .ZN(n1184) );
NAND4_X1 U891 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1154) );
AND4_X1 U892 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
NOR2_X1 U893 ( .A1(n1185), .A2(n1251), .ZN(n1245) );
AND3_X1 U894 ( .A1(n1252), .A2(n1253), .A3(n1089), .ZN(n1251) );
NOR3_X1 U895 ( .A1(n1254), .A2(n1255), .A3(n1087), .ZN(n1185) );
NAND4_X1 U896 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1244) );
INV_X1 U897 ( .A(KEYINPUT22), .ZN(n1259) );
NOR3_X1 U898 ( .A1(n1255), .A2(n1260), .A3(n1105), .ZN(n1258) );
NAND2_X1 U899 ( .A1(n1066), .A2(KEYINPUT22), .ZN(n1243) );
NOR3_X1 U900 ( .A1(n1088), .A2(n1255), .A3(n1254), .ZN(n1066) );
INV_X1 U901 ( .A(n1253), .ZN(n1254) );
XOR2_X1 U902 ( .A(n1153), .B(KEYINPUT34), .Z(n1242) );
NOR2_X1 U903 ( .A1(n1077), .A2(G952), .ZN(n1163) );
XNOR2_X1 U904 ( .A(G146), .B(n1221), .ZN(G48) );
NAND2_X1 U905 ( .A1(n1261), .A2(n1262), .ZN(n1221) );
XNOR2_X1 U906 ( .A(G143), .B(n1222), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1239), .A2(n1252), .A3(n1263), .A4(n1100), .ZN(n1222) );
NOR2_X1 U908 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U909 ( .A(G140), .B(n1266), .Z(G42) );
NOR4_X1 U910 ( .A1(KEYINPUT23), .A2(n1267), .A3(n1094), .A4(n1241), .ZN(n1266) );
XNOR2_X1 U911 ( .A(n1262), .B(KEYINPUT59), .ZN(n1267) );
XOR2_X1 U912 ( .A(G137), .B(n1228), .Z(G39) );
AND2_X1 U913 ( .A1(n1238), .A2(n1268), .ZN(n1228) );
INV_X1 U914 ( .A(n1241), .ZN(n1238) );
XNOR2_X1 U915 ( .A(n1141), .B(n1227), .ZN(G36) );
NOR3_X1 U916 ( .A1(n1095), .A2(n1088), .A3(n1241), .ZN(n1227) );
XOR2_X1 U917 ( .A(G131), .B(n1226), .Z(G33) );
NOR3_X1 U918 ( .A1(n1087), .A2(n1095), .A3(n1241), .ZN(n1226) );
NAND3_X1 U919 ( .A1(n1100), .A2(n1269), .A3(n1083), .ZN(n1241) );
NOR2_X1 U920 ( .A1(n1122), .A2(n1107), .ZN(n1083) );
INV_X1 U921 ( .A(n1262), .ZN(n1087) );
XNOR2_X1 U922 ( .A(n1270), .B(n1271), .ZN(G30) );
NOR2_X1 U923 ( .A1(KEYINPUT36), .A2(n1229), .ZN(n1271) );
NAND2_X1 U924 ( .A1(n1261), .A2(n1257), .ZN(n1229) );
AND4_X1 U925 ( .A1(n1272), .A2(n1239), .A3(n1100), .A4(n1273), .ZN(n1261) );
NAND3_X1 U926 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(G3) );
OR2_X1 U927 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND3_X1 U928 ( .A1(n1278), .A2(n1277), .A3(G101), .ZN(n1275) );
NAND2_X1 U929 ( .A1(n1279), .A2(n1196), .ZN(n1274) );
NAND2_X1 U930 ( .A1(n1280), .A2(n1277), .ZN(n1279) );
INV_X1 U931 ( .A(KEYINPUT31), .ZN(n1277) );
XNOR2_X1 U932 ( .A(KEYINPUT30), .B(n1278), .ZN(n1280) );
NAND3_X1 U933 ( .A1(n1253), .A2(n1281), .A3(n1252), .ZN(n1278) );
XOR2_X1 U934 ( .A(KEYINPUT8), .B(n1089), .Z(n1281) );
XOR2_X1 U935 ( .A(n1232), .B(n1282), .Z(G27) );
NAND2_X1 U936 ( .A1(KEYINPUT57), .A2(G125), .ZN(n1282) );
NAND4_X1 U937 ( .A1(n1239), .A2(n1262), .A3(n1235), .A4(n1084), .ZN(n1232) );
INV_X1 U938 ( .A(n1117), .ZN(n1084) );
AND2_X1 U939 ( .A1(n1283), .A2(n1269), .ZN(n1239) );
NAND2_X1 U940 ( .A1(n1109), .A2(n1284), .ZN(n1269) );
NAND4_X1 U941 ( .A1(G902), .A2(G953), .A3(n1285), .A4(n1136), .ZN(n1284) );
INV_X1 U942 ( .A(G900), .ZN(n1136) );
XOR2_X1 U943 ( .A(G122), .B(n1153), .Z(G24) );
AND4_X1 U944 ( .A1(n1286), .A2(n1085), .A3(n1118), .A4(n1287), .ZN(n1153) );
INV_X1 U945 ( .A(n1255), .ZN(n1085) );
NAND2_X1 U946 ( .A1(n1288), .A2(n1289), .ZN(n1255) );
XNOR2_X1 U947 ( .A(G119), .B(n1250), .ZN(G21) );
NAND2_X1 U948 ( .A1(n1268), .A2(n1286), .ZN(n1250) );
AND3_X1 U949 ( .A1(n1272), .A2(n1273), .A3(n1089), .ZN(n1268) );
XOR2_X1 U950 ( .A(G116), .B(n1290), .Z(G18) );
NOR3_X1 U951 ( .A1(KEYINPUT25), .A2(n1291), .A3(n1292), .ZN(n1290) );
NOR2_X1 U952 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NOR2_X1 U953 ( .A1(n1295), .A2(n1105), .ZN(n1293) );
NOR4_X1 U954 ( .A1(n1256), .A2(n1088), .A3(n1117), .A4(n1095), .ZN(n1295) );
INV_X1 U955 ( .A(n1257), .ZN(n1088) );
AND2_X1 U956 ( .A1(n1294), .A2(n1248), .ZN(n1291) );
NAND3_X1 U957 ( .A1(n1286), .A2(n1257), .A3(n1252), .ZN(n1248) );
NOR2_X1 U958 ( .A1(n1287), .A2(n1265), .ZN(n1257) );
INV_X1 U959 ( .A(n1118), .ZN(n1265) );
INV_X1 U960 ( .A(KEYINPUT39), .ZN(n1294) );
XNOR2_X1 U961 ( .A(G113), .B(n1249), .ZN(G15) );
NAND3_X1 U962 ( .A1(n1252), .A2(n1286), .A3(n1262), .ZN(n1249) );
NOR2_X1 U963 ( .A1(n1118), .A2(n1264), .ZN(n1262) );
INV_X1 U964 ( .A(n1287), .ZN(n1264) );
NOR3_X1 U965 ( .A1(n1105), .A2(n1256), .A3(n1117), .ZN(n1286) );
NAND2_X1 U966 ( .A1(n1102), .A2(n1296), .ZN(n1117) );
INV_X1 U967 ( .A(n1095), .ZN(n1252) );
NAND2_X1 U968 ( .A1(n1288), .A2(n1273), .ZN(n1095) );
XOR2_X1 U969 ( .A(n1247), .B(n1297), .Z(G12) );
XNOR2_X1 U970 ( .A(KEYINPUT18), .B(n1298), .ZN(n1297) );
NAND3_X1 U971 ( .A1(n1235), .A2(n1253), .A3(n1089), .ZN(n1247) );
NOR2_X1 U972 ( .A1(n1118), .A2(n1287), .ZN(n1089) );
XOR2_X1 U973 ( .A(n1299), .B(n1182), .Z(n1287) );
INV_X1 U974 ( .A(G475), .ZN(n1182) );
NAND2_X1 U975 ( .A1(KEYINPUT12), .A2(n1121), .ZN(n1299) );
NOR2_X1 U976 ( .A1(n1179), .A2(G902), .ZN(n1121) );
XNOR2_X1 U977 ( .A(n1300), .B(n1301), .ZN(n1179) );
XOR2_X1 U978 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U979 ( .A(G122), .B(n1304), .ZN(n1303) );
XNOR2_X1 U980 ( .A(n1305), .B(G131), .ZN(n1302) );
XOR2_X1 U981 ( .A(n1306), .B(n1307), .Z(n1300) );
XNOR2_X1 U982 ( .A(G104), .B(n1308), .ZN(n1307) );
NAND2_X1 U983 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U984 ( .A(KEYINPUT55), .B(KEYINPUT52), .Z(n1310) );
XOR2_X1 U985 ( .A(n1311), .B(G143), .Z(n1309) );
NAND2_X1 U986 ( .A1(n1312), .A2(G214), .ZN(n1311) );
NAND2_X1 U987 ( .A1(KEYINPUT17), .A2(n1143), .ZN(n1306) );
XNOR2_X1 U988 ( .A(n1313), .B(G478), .ZN(n1118) );
OR2_X1 U989 ( .A1(n1174), .A2(G902), .ZN(n1313) );
XOR2_X1 U990 ( .A(n1314), .B(n1315), .Z(n1174) );
XNOR2_X1 U991 ( .A(n1068), .B(n1316), .ZN(n1315) );
NOR2_X1 U992 ( .A1(KEYINPUT29), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U993 ( .A(n1270), .B(n1318), .ZN(n1317) );
XNOR2_X1 U994 ( .A(G143), .B(n1141), .ZN(n1318) );
XOR2_X1 U995 ( .A(n1319), .B(n1320), .Z(n1314) );
NOR2_X1 U996 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U997 ( .A(n1323), .B(KEYINPUT24), .Z(n1322) );
NAND2_X1 U998 ( .A1(G122), .A2(n1324), .ZN(n1323) );
NOR2_X1 U999 ( .A1(G122), .A2(n1324), .ZN(n1321) );
XOR2_X1 U1000 ( .A(KEYINPUT27), .B(G116), .Z(n1324) );
NAND2_X1 U1001 ( .A1(G217), .A2(n1325), .ZN(n1319) );
NOR3_X1 U1002 ( .A1(n1260), .A2(n1256), .A3(n1105), .ZN(n1253) );
INV_X1 U1003 ( .A(n1283), .ZN(n1105) );
NOR2_X1 U1004 ( .A1(n1108), .A2(n1107), .ZN(n1283) );
AND2_X1 U1005 ( .A1(G214), .A2(n1326), .ZN(n1107) );
INV_X1 U1006 ( .A(n1122), .ZN(n1108) );
XNOR2_X1 U1007 ( .A(n1327), .B(n1219), .ZN(n1122) );
AND2_X1 U1008 ( .A1(G210), .A2(n1326), .ZN(n1219) );
NAND2_X1 U1009 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
NAND2_X1 U1010 ( .A1(n1330), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1011 ( .A(n1331), .B(n1332), .Z(n1330) );
NOR2_X1 U1012 ( .A1(KEYINPUT54), .A2(n1218), .ZN(n1332) );
XNOR2_X1 U1013 ( .A(n1333), .B(n1162), .ZN(n1218) );
XNOR2_X1 U1014 ( .A(n1334), .B(n1335), .ZN(n1162) );
XNOR2_X1 U1015 ( .A(KEYINPUT35), .B(n1196), .ZN(n1335) );
XNOR2_X1 U1016 ( .A(n1336), .B(n1337), .ZN(n1333) );
INV_X1 U1017 ( .A(n1159), .ZN(n1337) );
XOR2_X1 U1018 ( .A(G110), .B(n1338), .Z(n1159) );
XOR2_X1 U1019 ( .A(KEYINPUT2), .B(G122), .Z(n1338) );
NAND2_X1 U1020 ( .A1(n1339), .A2(n1161), .ZN(n1336) );
NAND3_X1 U1021 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1161) );
NAND2_X1 U1022 ( .A1(n1343), .A2(G113), .ZN(n1342) );
NAND3_X1 U1023 ( .A1(G116), .A2(n1304), .A3(G119), .ZN(n1341) );
INV_X1 U1024 ( .A(G113), .ZN(n1304) );
NAND2_X1 U1025 ( .A1(n1344), .A2(n1345), .ZN(n1340) );
XNOR2_X1 U1026 ( .A(G113), .B(G116), .ZN(n1344) );
XOR2_X1 U1027 ( .A(KEYINPUT47), .B(KEYINPUT44), .Z(n1339) );
NAND2_X1 U1028 ( .A1(n1346), .A2(n1347), .ZN(n1331) );
NAND2_X1 U1029 ( .A1(KEYINPUT37), .A2(n1216), .ZN(n1347) );
XOR2_X1 U1030 ( .A(n1348), .B(n1213), .Z(n1346) );
AND2_X1 U1031 ( .A1(G224), .A2(n1349), .ZN(n1213) );
OR2_X1 U1032 ( .A1(n1216), .A2(KEYINPUT37), .ZN(n1348) );
XOR2_X1 U1033 ( .A(G125), .B(n1202), .Z(n1216) );
AND2_X1 U1034 ( .A1(n1350), .A2(n1109), .ZN(n1256) );
NAND3_X1 U1035 ( .A1(n1285), .A2(n1077), .A3(G952), .ZN(n1109) );
NAND3_X1 U1036 ( .A1(n1157), .A2(n1285), .A3(G902), .ZN(n1350) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1285) );
NOR2_X1 U1038 ( .A1(n1077), .A2(G898), .ZN(n1157) );
INV_X1 U1039 ( .A(G953), .ZN(n1077) );
INV_X1 U1040 ( .A(n1100), .ZN(n1260) );
NOR2_X1 U1041 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
INV_X1 U1042 ( .A(n1296), .ZN(n1103) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1351), .ZN(n1296) );
XOR2_X1 U1044 ( .A(n1352), .B(G469), .Z(n1102) );
NAND2_X1 U1045 ( .A1(n1353), .A2(n1329), .ZN(n1352) );
XOR2_X1 U1046 ( .A(n1354), .B(n1206), .Z(n1353) );
XNOR2_X1 U1047 ( .A(G140), .B(n1298), .ZN(n1206) );
XNOR2_X1 U1048 ( .A(n1207), .B(n1355), .ZN(n1354) );
NOR2_X1 U1049 ( .A1(KEYINPUT4), .A2(n1209), .ZN(n1355) );
NAND2_X1 U1050 ( .A1(G227), .A2(n1349), .ZN(n1209) );
XNOR2_X1 U1051 ( .A(n1142), .B(n1356), .ZN(n1207) );
XOR2_X1 U1052 ( .A(n1357), .B(n1358), .Z(n1356) );
NAND2_X1 U1053 ( .A1(n1359), .A2(n1360), .ZN(n1357) );
NAND2_X1 U1054 ( .A1(G101), .A2(n1334), .ZN(n1360) );
XOR2_X1 U1055 ( .A(n1361), .B(KEYINPUT40), .Z(n1359) );
OR2_X1 U1056 ( .A1(n1334), .A2(G101), .ZN(n1361) );
XNOR2_X1 U1057 ( .A(G104), .B(n1068), .ZN(n1334) );
INV_X1 U1058 ( .A(G107), .ZN(n1068) );
XNOR2_X1 U1059 ( .A(G128), .B(n1362), .ZN(n1142) );
INV_X1 U1060 ( .A(n1094), .ZN(n1235) );
NAND2_X1 U1061 ( .A1(n1272), .A2(n1289), .ZN(n1094) );
XOR2_X1 U1062 ( .A(n1273), .B(KEYINPUT41), .Z(n1289) );
XNOR2_X1 U1063 ( .A(n1127), .B(G472), .ZN(n1273) );
NAND2_X1 U1064 ( .A1(n1363), .A2(n1329), .ZN(n1127) );
XOR2_X1 U1065 ( .A(n1198), .B(n1364), .Z(n1363) );
XOR2_X1 U1066 ( .A(n1365), .B(n1202), .Z(n1364) );
XOR2_X1 U1067 ( .A(n1362), .B(n1366), .Z(n1202) );
NOR2_X1 U1068 ( .A1(G128), .A2(KEYINPUT10), .ZN(n1366) );
XNOR2_X1 U1069 ( .A(G143), .B(n1305), .ZN(n1362) );
INV_X1 U1070 ( .A(G146), .ZN(n1305) );
NOR2_X1 U1071 ( .A1(n1194), .A2(n1367), .ZN(n1365) );
XOR2_X1 U1072 ( .A(KEYINPUT9), .B(n1368), .Z(n1367) );
NOR2_X1 U1073 ( .A1(G101), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1074 ( .A(n1193), .B(KEYINPUT49), .Z(n1369) );
NOR2_X1 U1075 ( .A1(n1193), .A2(n1196), .ZN(n1194) );
INV_X1 U1076 ( .A(G101), .ZN(n1196) );
NAND2_X1 U1077 ( .A1(n1312), .A2(G210), .ZN(n1193) );
AND2_X1 U1078 ( .A1(n1349), .A2(n1328), .ZN(n1312) );
INV_X1 U1079 ( .A(G237), .ZN(n1328) );
XOR2_X1 U1080 ( .A(n1358), .B(n1370), .Z(n1198) );
XNOR2_X1 U1081 ( .A(G113), .B(n1371), .ZN(n1370) );
NAND2_X1 U1082 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
NAND2_X1 U1083 ( .A1(G116), .A2(n1345), .ZN(n1373) );
XNOR2_X1 U1084 ( .A(n1343), .B(KEYINPUT0), .ZN(n1372) );
NOR2_X1 U1085 ( .A1(n1345), .A2(G116), .ZN(n1343) );
INV_X1 U1086 ( .A(G119), .ZN(n1345) );
XOR2_X1 U1087 ( .A(n1374), .B(n1139), .Z(n1358) );
XOR2_X1 U1088 ( .A(G131), .B(G137), .Z(n1139) );
NAND2_X1 U1089 ( .A1(n1375), .A2(n1141), .ZN(n1374) );
INV_X1 U1090 ( .A(G134), .ZN(n1141) );
XNOR2_X1 U1091 ( .A(KEYINPUT42), .B(KEYINPUT26), .ZN(n1375) );
INV_X1 U1092 ( .A(n1288), .ZN(n1272) );
XOR2_X1 U1093 ( .A(n1376), .B(n1124), .Z(n1288) );
NAND2_X1 U1094 ( .A1(n1168), .A2(n1329), .ZN(n1124) );
XNOR2_X1 U1095 ( .A(n1377), .B(n1378), .ZN(n1168) );
XOR2_X1 U1096 ( .A(KEYINPUT61), .B(G137), .Z(n1378) );
XOR2_X1 U1097 ( .A(n1379), .B(n1380), .Z(n1377) );
AND2_X1 U1098 ( .A1(G221), .A2(n1325), .ZN(n1380) );
AND2_X1 U1099 ( .A1(G234), .A2(n1349), .ZN(n1325) );
XNOR2_X1 U1100 ( .A(G953), .B(KEYINPUT20), .ZN(n1349) );
NAND3_X1 U1101 ( .A1(n1381), .A2(n1382), .A3(n1383), .ZN(n1379) );
NAND2_X1 U1102 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
NAND3_X1 U1103 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1385) );
NAND2_X1 U1104 ( .A1(KEYINPUT28), .A2(KEYINPUT33), .ZN(n1388) );
NAND2_X1 U1105 ( .A1(KEYINPUT63), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1106 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
NAND2_X1 U1107 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1108 ( .A1(n1390), .A2(n1394), .ZN(n1386) );
INV_X1 U1109 ( .A(KEYINPUT63), .ZN(n1394) );
NAND4_X1 U1110 ( .A1(n1390), .A2(n1395), .A3(KEYINPUT28), .A4(n1393), .ZN(n1382) );
INV_X1 U1111 ( .A(KEYINPUT33), .ZN(n1393) );
NAND2_X1 U1112 ( .A1(KEYINPUT33), .A2(n1396), .ZN(n1381) );
NAND2_X1 U1113 ( .A1(n1390), .A2(n1397), .ZN(n1396) );
NAND2_X1 U1114 ( .A1(n1395), .A2(n1392), .ZN(n1397) );
INV_X1 U1115 ( .A(KEYINPUT28), .ZN(n1392) );
INV_X1 U1116 ( .A(n1384), .ZN(n1395) );
XNOR2_X1 U1117 ( .A(n1398), .B(n1143), .ZN(n1384) );
XOR2_X1 U1118 ( .A(G125), .B(G140), .Z(n1143) );
XNOR2_X1 U1119 ( .A(G146), .B(KEYINPUT5), .ZN(n1398) );
XOR2_X1 U1120 ( .A(n1399), .B(n1400), .Z(n1390) );
XNOR2_X1 U1121 ( .A(n1270), .B(G119), .ZN(n1400) );
INV_X1 U1122 ( .A(G128), .ZN(n1270) );
NAND2_X1 U1123 ( .A1(KEYINPUT51), .A2(n1298), .ZN(n1399) );
INV_X1 U1124 ( .A(G110), .ZN(n1298) );
NAND2_X1 U1125 ( .A1(KEYINPUT19), .A2(n1125), .ZN(n1376) );
NAND2_X1 U1126 ( .A1(G217), .A2(n1351), .ZN(n1125) );
NAND2_X1 U1127 ( .A1(G234), .A2(n1329), .ZN(n1351) );
INV_X1 U1128 ( .A(G902), .ZN(n1329) );
endmodule


