//Key = 0011000101100000001100010011111001001000001110110000101001001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;

XNOR2_X1 U763 ( .A(n1061), .B(n1062), .ZN(G9) );
NAND2_X1 U764 ( .A1(KEYINPUT33), .A2(G107), .ZN(n1062) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(G75) );
NOR4_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
NOR2_X1 U767 ( .A1(KEYINPUT10), .A2(n1069), .ZN(n1068) );
NOR4_X1 U768 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1073), .ZN(n1067) );
NOR2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U772 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1070), .ZN(n1080) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1082) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U781 ( .A1(n1096), .A2(n1072), .ZN(n1079) );
NOR2_X1 U782 ( .A1(n1097), .A2(n1072), .ZN(n1075) );
INV_X1 U783 ( .A(n1098), .ZN(n1072) );
NOR2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1070), .ZN(n1100) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
AND2_X1 U787 ( .A1(n1104), .A2(KEYINPUT10), .ZN(n1102) );
NOR4_X1 U788 ( .A1(n1105), .A2(n1106), .A3(n1078), .A4(n1107), .ZN(n1099) );
NAND3_X1 U789 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1065) );
NAND3_X1 U790 ( .A1(n1111), .A2(n1095), .A3(n1112), .ZN(n1110) );
INV_X1 U791 ( .A(KEYINPUT30), .ZN(n1095) );
OR4_X1 U792 ( .A1(n1073), .A2(n1070), .A3(n1094), .A4(n1078), .ZN(n1111) );
INV_X1 U793 ( .A(n1113), .ZN(n1078) );
AND3_X1 U794 ( .A1(n1108), .A2(n1109), .A3(n1114), .ZN(n1063) );
NAND4_X1 U795 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1108) );
NOR3_X1 U796 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NOR2_X1 U797 ( .A1(G472), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U798 ( .A(n1123), .B(KEYINPUT7), .ZN(n1120) );
NAND3_X1 U799 ( .A1(n1089), .A2(n1124), .A3(n1125), .ZN(n1119) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U801 ( .A(n1128), .B(KEYINPUT57), .Z(n1126) );
NOR3_X1 U802 ( .A1(n1070), .A2(n1129), .A3(n1130), .ZN(n1117) );
NOR2_X1 U803 ( .A1(KEYINPUT18), .A2(G472), .ZN(n1130) );
AND3_X1 U804 ( .A1(G472), .A2(n1122), .A3(KEYINPUT18), .ZN(n1129) );
INV_X1 U805 ( .A(n1131), .ZN(n1070) );
NAND2_X1 U806 ( .A1(n1132), .A2(n1133), .ZN(G72) );
NAND3_X1 U807 ( .A1(n1134), .A2(n1135), .A3(G953), .ZN(n1133) );
XNOR2_X1 U808 ( .A(KEYINPUT49), .B(n1136), .ZN(n1134) );
XOR2_X1 U809 ( .A(n1137), .B(KEYINPUT58), .Z(n1132) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1138), .ZN(n1137) );
NAND2_X1 U811 ( .A1(G953), .A2(n1135), .ZN(n1138) );
NAND2_X1 U812 ( .A1(G900), .A2(G227), .ZN(n1135) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND3_X1 U814 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
XOR2_X1 U815 ( .A(n1144), .B(KEYINPUT55), .Z(n1139) );
NAND2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1142), .ZN(n1146) );
INV_X1 U818 ( .A(n1147), .ZN(n1142) );
XNOR2_X1 U819 ( .A(n1148), .B(n1149), .ZN(n1143) );
XNOR2_X1 U820 ( .A(n1150), .B(n1151), .ZN(n1149) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U823 ( .A(KEYINPUT17), .B(n1156), .Z(n1155) );
AND2_X1 U824 ( .A1(n1157), .A2(G134), .ZN(n1156) );
NOR2_X1 U825 ( .A1(G134), .A2(n1157), .ZN(n1154) );
NAND2_X1 U826 ( .A1(KEYINPUT44), .A2(n1158), .ZN(n1152) );
INV_X1 U827 ( .A(n1141), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1109), .A2(n1159), .ZN(n1141) );
NAND2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U830 ( .A(n1162), .B(KEYINPUT6), .Z(n1160) );
XOR2_X1 U831 ( .A(n1163), .B(n1164), .Z(G69) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U833 ( .A1(n1167), .A2(G953), .ZN(n1166) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
XNOR2_X1 U835 ( .A(n1170), .B(n1171), .ZN(n1169) );
NOR2_X1 U836 ( .A1(n1172), .A2(n1109), .ZN(n1163) );
AND2_X1 U837 ( .A1(G224), .A2(G898), .ZN(n1172) );
NOR2_X1 U838 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U840 ( .A1(n1177), .A2(n1105), .A3(n1178), .ZN(n1175) );
NOR2_X1 U841 ( .A1(n1179), .A2(n1180), .ZN(n1173) );
XNOR2_X1 U842 ( .A(KEYINPUT40), .B(G953), .ZN(n1180) );
XNOR2_X1 U843 ( .A(G952), .B(KEYINPUT23), .ZN(n1179) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(G63) );
XOR2_X1 U845 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U846 ( .A1(n1185), .A2(n1177), .ZN(n1184) );
NOR2_X1 U847 ( .A1(KEYINPUT51), .A2(n1186), .ZN(n1183) );
XNOR2_X1 U848 ( .A(n1187), .B(KEYINPUT43), .ZN(n1186) );
NOR2_X1 U849 ( .A1(n1181), .A2(n1188), .ZN(G60) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U851 ( .A1(n1191), .A2(n1177), .ZN(n1189) );
XOR2_X1 U852 ( .A(G104), .B(n1192), .Z(G6) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U854 ( .A1(n1181), .A2(n1195), .ZN(G57) );
XOR2_X1 U855 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U856 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U857 ( .A1(KEYINPUT12), .A2(n1200), .ZN(n1199) );
NOR2_X1 U858 ( .A1(n1201), .A2(n1177), .ZN(n1198) );
INV_X1 U859 ( .A(G472), .ZN(n1201) );
NOR2_X1 U860 ( .A1(n1181), .A2(n1202), .ZN(G54) );
XOR2_X1 U861 ( .A(n1203), .B(n1204), .Z(n1202) );
XNOR2_X1 U862 ( .A(n1151), .B(n1205), .ZN(n1204) );
XOR2_X1 U863 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U864 ( .A1(n1208), .A2(n1177), .ZN(n1206) );
XOR2_X1 U865 ( .A(n1209), .B(n1210), .Z(n1203) );
XNOR2_X1 U866 ( .A(G140), .B(n1211), .ZN(n1210) );
NOR2_X1 U867 ( .A1(n1181), .A2(n1212), .ZN(G51) );
XOR2_X1 U868 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U869 ( .A(KEYINPUT38), .B(n1215), .Z(n1214) );
NOR2_X1 U870 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U871 ( .A(KEYINPUT63), .B(n1218), .Z(n1217) );
NOR2_X1 U872 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U873 ( .A(n1221), .B(KEYINPUT20), .Z(n1219) );
AND2_X1 U874 ( .A1(n1220), .A2(n1221), .ZN(n1216) );
XOR2_X1 U875 ( .A(n1222), .B(n1223), .Z(n1220) );
NOR2_X1 U876 ( .A1(KEYINPUT53), .A2(n1224), .ZN(n1223) );
NOR2_X1 U877 ( .A1(n1128), .A2(n1177), .ZN(n1213) );
NAND2_X1 U878 ( .A1(G902), .A2(n1066), .ZN(n1177) );
NAND3_X1 U879 ( .A1(n1161), .A2(n1162), .A3(n1167), .ZN(n1066) );
AND2_X1 U880 ( .A1(n1225), .A2(n1226), .ZN(n1167) );
NOR4_X1 U881 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
INV_X1 U882 ( .A(n1231), .ZN(n1227) );
NOR4_X1 U883 ( .A1(n1232), .A2(n1061), .A3(n1233), .A4(n1234), .ZN(n1225) );
NOR2_X1 U884 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U885 ( .A(n1237), .B(KEYINPUT50), .ZN(n1236) );
INV_X1 U886 ( .A(n1087), .ZN(n1235) );
NOR2_X1 U887 ( .A1(n1238), .A2(n1193), .ZN(n1233) );
XOR2_X1 U888 ( .A(n1194), .B(KEYINPUT4), .Z(n1238) );
NAND4_X1 U889 ( .A1(n1093), .A2(n1113), .A3(n1239), .A4(n1240), .ZN(n1194) );
AND3_X1 U890 ( .A1(n1241), .A2(n1113), .A3(n1242), .ZN(n1061) );
INV_X1 U891 ( .A(n1243), .ZN(n1232) );
AND4_X1 U892 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1161) );
AND4_X1 U893 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
NAND2_X1 U894 ( .A1(n1252), .A2(n1112), .ZN(n1246) );
XOR2_X1 U895 ( .A(n1253), .B(KEYINPUT26), .Z(n1252) );
NAND2_X1 U896 ( .A1(n1254), .A2(n1087), .ZN(n1244) );
AND2_X1 U897 ( .A1(n1255), .A2(n1114), .ZN(n1181) );
INV_X1 U898 ( .A(G952), .ZN(n1114) );
XNOR2_X1 U899 ( .A(KEYINPUT40), .B(n1109), .ZN(n1255) );
XNOR2_X1 U900 ( .A(n1245), .B(n1256), .ZN(G48) );
NOR2_X1 U901 ( .A1(KEYINPUT22), .A2(n1257), .ZN(n1256) );
NAND4_X1 U902 ( .A1(n1258), .A2(n1093), .A3(n1259), .A4(n1087), .ZN(n1245) );
XOR2_X1 U903 ( .A(n1251), .B(n1260), .Z(G45) );
XNOR2_X1 U904 ( .A(G143), .B(KEYINPUT32), .ZN(n1260) );
NAND4_X1 U905 ( .A1(n1261), .A2(n1262), .A3(n1087), .A4(n1123), .ZN(n1251) );
XNOR2_X1 U906 ( .A(KEYINPUT62), .B(n1263), .ZN(n1262) );
XOR2_X1 U907 ( .A(G140), .B(n1264), .Z(G42) );
NOR2_X1 U908 ( .A1(KEYINPUT37), .A2(n1250), .ZN(n1264) );
NAND3_X1 U909 ( .A1(n1258), .A2(n1112), .A3(n1265), .ZN(n1250) );
XNOR2_X1 U910 ( .A(G137), .B(n1162), .ZN(G39) );
NAND3_X1 U911 ( .A1(n1098), .A2(n1259), .A3(n1258), .ZN(n1162) );
NOR2_X1 U912 ( .A1(n1091), .A2(n1085), .ZN(n1098) );
INV_X1 U913 ( .A(n1266), .ZN(n1085) );
XNOR2_X1 U914 ( .A(G134), .B(n1267), .ZN(G36) );
NOR2_X1 U915 ( .A1(KEYINPUT16), .A2(n1268), .ZN(n1267) );
NOR2_X1 U916 ( .A1(n1253), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U917 ( .A(KEYINPUT27), .B(n1091), .ZN(n1269) );
INV_X1 U918 ( .A(n1112), .ZN(n1091) );
NAND2_X1 U919 ( .A1(n1261), .A2(n1241), .ZN(n1253) );
XNOR2_X1 U920 ( .A(G131), .B(n1249), .ZN(G33) );
NAND3_X1 U921 ( .A1(n1112), .A2(n1093), .A3(n1261), .ZN(n1249) );
AND2_X1 U922 ( .A1(n1258), .A2(n1104), .ZN(n1261) );
NOR2_X1 U923 ( .A1(n1096), .A2(n1270), .ZN(n1258) );
INV_X1 U924 ( .A(n1271), .ZN(n1270) );
NOR2_X1 U925 ( .A1(n1088), .A2(n1272), .ZN(n1112) );
INV_X1 U926 ( .A(n1089), .ZN(n1272) );
XNOR2_X1 U927 ( .A(G128), .B(n1273), .ZN(G30) );
NAND2_X1 U928 ( .A1(n1274), .A2(n1254), .ZN(n1273) );
AND4_X1 U929 ( .A1(n1239), .A2(n1241), .A3(n1259), .A4(n1271), .ZN(n1254) );
XNOR2_X1 U930 ( .A(n1087), .B(KEYINPUT28), .ZN(n1274) );
XNOR2_X1 U931 ( .A(G101), .B(n1243), .ZN(G3) );
NAND3_X1 U932 ( .A1(n1266), .A2(n1242), .A3(n1104), .ZN(n1243) );
XNOR2_X1 U933 ( .A(G125), .B(n1248), .ZN(G27) );
NAND4_X1 U934 ( .A1(n1265), .A2(n1131), .A3(n1087), .A4(n1271), .ZN(n1248) );
NAND2_X1 U935 ( .A1(n1275), .A2(n1073), .ZN(n1271) );
NAND3_X1 U936 ( .A1(G902), .A2(n1276), .A3(n1147), .ZN(n1275) );
NOR2_X1 U937 ( .A1(n1277), .A2(G900), .ZN(n1147) );
AND2_X1 U938 ( .A1(n1093), .A2(n1103), .ZN(n1265) );
XOR2_X1 U939 ( .A(n1278), .B(n1279), .Z(G24) );
NOR2_X1 U940 ( .A1(KEYINPUT11), .A2(n1280), .ZN(n1279) );
XOR2_X1 U941 ( .A(KEYINPUT8), .B(G122), .Z(n1280) );
NAND2_X1 U942 ( .A1(n1237), .A2(n1087), .ZN(n1278) );
AND4_X1 U943 ( .A1(n1281), .A2(n1113), .A3(n1282), .A4(n1283), .ZN(n1237) );
OR2_X1 U944 ( .A1(n1093), .A2(KEYINPUT62), .ZN(n1283) );
NAND2_X1 U945 ( .A1(KEYINPUT62), .A2(n1284), .ZN(n1282) );
NAND2_X1 U946 ( .A1(n1263), .A2(n1123), .ZN(n1284) );
NOR2_X1 U947 ( .A1(n1285), .A2(n1286), .ZN(n1113) );
XOR2_X1 U948 ( .A(G119), .B(n1230), .Z(G21) );
AND4_X1 U949 ( .A1(n1281), .A2(n1266), .A3(n1259), .A4(n1087), .ZN(n1230) );
NAND2_X1 U950 ( .A1(n1287), .A2(n1288), .ZN(n1259) );
NAND2_X1 U951 ( .A1(n1103), .A2(n1289), .ZN(n1288) );
INV_X1 U952 ( .A(KEYINPUT36), .ZN(n1289) );
NAND3_X1 U953 ( .A1(n1286), .A2(n1285), .A3(KEYINPUT36), .ZN(n1287) );
XOR2_X1 U954 ( .A(G116), .B(n1229), .Z(G18) );
AND4_X1 U955 ( .A1(n1281), .A2(n1104), .A3(n1241), .A4(n1087), .ZN(n1229) );
XOR2_X1 U956 ( .A(n1290), .B(KEYINPUT14), .Z(n1087) );
INV_X1 U957 ( .A(n1094), .ZN(n1241) );
NAND2_X1 U958 ( .A1(n1263), .A2(n1291), .ZN(n1094) );
XOR2_X1 U959 ( .A(G113), .B(n1228), .Z(G15) );
AND4_X1 U960 ( .A1(n1093), .A2(n1281), .A3(n1104), .A4(n1290), .ZN(n1228) );
INV_X1 U961 ( .A(n1071), .ZN(n1104) );
NAND2_X1 U962 ( .A1(n1292), .A2(n1116), .ZN(n1071) );
XNOR2_X1 U963 ( .A(n1286), .B(KEYINPUT36), .ZN(n1292) );
AND2_X1 U964 ( .A1(n1131), .A2(n1240), .ZN(n1281) );
NOR2_X1 U965 ( .A1(n1107), .A2(n1293), .ZN(n1131) );
NOR2_X1 U966 ( .A1(n1106), .A2(n1105), .ZN(n1293) );
NOR2_X1 U967 ( .A1(n1291), .A2(n1263), .ZN(n1093) );
INV_X1 U968 ( .A(n1123), .ZN(n1291) );
XNOR2_X1 U969 ( .A(G110), .B(n1231), .ZN(G12) );
NAND3_X1 U970 ( .A1(n1103), .A2(n1242), .A3(n1266), .ZN(n1231) );
NOR2_X1 U971 ( .A1(n1123), .A2(n1263), .ZN(n1266) );
XOR2_X1 U972 ( .A(n1115), .B(KEYINPUT54), .Z(n1263) );
XNOR2_X1 U973 ( .A(n1294), .B(n1185), .ZN(n1115) );
INV_X1 U974 ( .A(G478), .ZN(n1185) );
NAND2_X1 U975 ( .A1(n1187), .A2(n1295), .ZN(n1294) );
XNOR2_X1 U976 ( .A(n1296), .B(n1297), .ZN(n1187) );
XNOR2_X1 U977 ( .A(n1298), .B(n1299), .ZN(n1297) );
XOR2_X1 U978 ( .A(G134), .B(G122), .Z(n1299) );
XNOR2_X1 U979 ( .A(n1300), .B(n1301), .ZN(n1296) );
XOR2_X1 U980 ( .A(n1302), .B(n1303), .Z(n1300) );
NOR2_X1 U981 ( .A1(n1304), .A2(n1178), .ZN(n1303) );
NAND2_X1 U982 ( .A1(KEYINPUT47), .A2(n1305), .ZN(n1302) );
XOR2_X1 U983 ( .A(n1306), .B(n1191), .Z(n1123) );
INV_X1 U984 ( .A(G475), .ZN(n1191) );
OR2_X1 U985 ( .A1(n1190), .A2(G902), .ZN(n1306) );
XNOR2_X1 U986 ( .A(n1307), .B(n1308), .ZN(n1190) );
XOR2_X1 U987 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U988 ( .A(G113), .B(G104), .Z(n1310) );
XOR2_X1 U989 ( .A(G131), .B(G122), .Z(n1309) );
XOR2_X1 U990 ( .A(n1311), .B(n1312), .Z(n1307) );
XNOR2_X1 U991 ( .A(n1158), .B(n1313), .ZN(n1311) );
AND2_X1 U992 ( .A1(G214), .A2(n1314), .ZN(n1313) );
XOR2_X1 U993 ( .A(G140), .B(n1224), .Z(n1158) );
AND3_X1 U994 ( .A1(n1239), .A2(n1240), .A3(n1290), .ZN(n1242) );
INV_X1 U995 ( .A(n1193), .ZN(n1290) );
NAND2_X1 U996 ( .A1(n1089), .A2(n1088), .ZN(n1193) );
NAND2_X1 U997 ( .A1(n1315), .A2(n1124), .ZN(n1088) );
NAND2_X1 U998 ( .A1(n1316), .A2(n1128), .ZN(n1124) );
INV_X1 U999 ( .A(n1127), .ZN(n1316) );
XOR2_X1 U1000 ( .A(n1317), .B(KEYINPUT15), .Z(n1315) );
NAND2_X1 U1001 ( .A1(n1318), .A2(n1127), .ZN(n1317) );
NAND2_X1 U1002 ( .A1(n1319), .A2(n1295), .ZN(n1127) );
XNOR2_X1 U1003 ( .A(n1320), .B(n1321), .ZN(n1319) );
INV_X1 U1004 ( .A(n1222), .ZN(n1321) );
XNOR2_X1 U1005 ( .A(n1322), .B(n1323), .ZN(n1222) );
NAND2_X1 U1006 ( .A1(G224), .A2(n1109), .ZN(n1322) );
XOR2_X1 U1007 ( .A(n1221), .B(n1224), .Z(n1320) );
XOR2_X1 U1008 ( .A(n1324), .B(n1170), .Z(n1221) );
XOR2_X1 U1009 ( .A(n1325), .B(n1326), .Z(n1170) );
XOR2_X1 U1010 ( .A(G113), .B(n1327), .Z(n1326) );
NOR2_X1 U1011 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1012 ( .A(n1330), .B(KEYINPUT9), .Z(n1329) );
NAND2_X1 U1013 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NOR2_X1 U1014 ( .A1(n1332), .A2(n1331), .ZN(n1328) );
XOR2_X1 U1015 ( .A(n1333), .B(n1334), .Z(n1331) );
XOR2_X1 U1016 ( .A(G104), .B(KEYINPUT52), .Z(n1334) );
NOR2_X1 U1017 ( .A1(KEYINPUT24), .A2(n1298), .ZN(n1333) );
NAND2_X1 U1018 ( .A1(KEYINPUT61), .A2(n1171), .ZN(n1324) );
XNOR2_X1 U1019 ( .A(G122), .B(G110), .ZN(n1171) );
XNOR2_X1 U1020 ( .A(KEYINPUT39), .B(n1128), .ZN(n1318) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1335), .ZN(n1128) );
NAND2_X1 U1022 ( .A1(n1336), .A2(n1335), .ZN(n1089) );
NAND2_X1 U1023 ( .A1(n1337), .A2(n1295), .ZN(n1335) );
INV_X1 U1024 ( .A(G237), .ZN(n1337) );
XOR2_X1 U1025 ( .A(KEYINPUT45), .B(G214), .Z(n1336) );
NAND2_X1 U1026 ( .A1(n1073), .A2(n1338), .ZN(n1240) );
NAND3_X1 U1027 ( .A1(n1168), .A2(n1276), .A3(G902), .ZN(n1338) );
NOR2_X1 U1028 ( .A1(n1277), .A2(G898), .ZN(n1168) );
XNOR2_X1 U1029 ( .A(G953), .B(KEYINPUT13), .ZN(n1277) );
NAND3_X1 U1030 ( .A1(n1276), .A2(n1109), .A3(G952), .ZN(n1073) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1276) );
XOR2_X1 U1032 ( .A(n1096), .B(KEYINPUT3), .Z(n1239) );
NAND2_X1 U1033 ( .A1(n1107), .A2(n1339), .ZN(n1096) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1035 ( .A(n1341), .B(n1208), .Z(n1107) );
INV_X1 U1036 ( .A(G469), .ZN(n1208) );
NAND2_X1 U1037 ( .A1(n1342), .A2(n1295), .ZN(n1341) );
XOR2_X1 U1038 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1039 ( .A(n1345), .B(n1207), .Z(n1344) );
XNOR2_X1 U1040 ( .A(n1346), .B(n1347), .ZN(n1207) );
NAND3_X1 U1041 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1346) );
OR2_X1 U1042 ( .A1(n1332), .A2(KEYINPUT29), .ZN(n1350) );
NAND3_X1 U1043 ( .A1(KEYINPUT29), .A2(n1351), .A3(n1352), .ZN(n1349) );
OR2_X1 U1044 ( .A1(n1352), .A2(n1351), .ZN(n1348) );
NOR2_X1 U1045 ( .A1(G101), .A2(KEYINPUT31), .ZN(n1351) );
XNOR2_X1 U1046 ( .A(G104), .B(n1298), .ZN(n1352) );
INV_X1 U1047 ( .A(G107), .ZN(n1298) );
NOR2_X1 U1048 ( .A1(KEYINPUT59), .A2(n1151), .ZN(n1345) );
XOR2_X1 U1049 ( .A(n1353), .B(n1354), .Z(n1151) );
NAND2_X1 U1050 ( .A1(KEYINPUT60), .A2(n1312), .ZN(n1353) );
XNOR2_X1 U1051 ( .A(n1355), .B(G146), .ZN(n1312) );
INV_X1 U1052 ( .A(G143), .ZN(n1355) );
XNOR2_X1 U1053 ( .A(n1356), .B(n1209), .ZN(n1343) );
NAND2_X1 U1054 ( .A1(G227), .A2(n1109), .ZN(n1209) );
NAND2_X1 U1055 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
NAND2_X1 U1056 ( .A1(G140), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1057 ( .A(n1360), .B(KEYINPUT5), .Z(n1357) );
OR2_X1 U1058 ( .A1(n1359), .A2(G140), .ZN(n1360) );
XOR2_X1 U1059 ( .A(n1211), .B(KEYINPUT41), .Z(n1359) );
INV_X1 U1060 ( .A(G110), .ZN(n1211) );
NOR2_X1 U1061 ( .A1(n1286), .A2(n1116), .ZN(n1103) );
INV_X1 U1062 ( .A(n1285), .ZN(n1116) );
XNOR2_X1 U1063 ( .A(n1361), .B(n1362), .ZN(n1285) );
NOR2_X1 U1064 ( .A1(n1105), .A2(n1363), .ZN(n1362) );
XNOR2_X1 U1065 ( .A(KEYINPUT2), .B(n1178), .ZN(n1363) );
INV_X1 U1066 ( .A(G217), .ZN(n1178) );
INV_X1 U1067 ( .A(n1340), .ZN(n1105) );
NAND2_X1 U1068 ( .A1(n1364), .A2(G234), .ZN(n1340) );
XNOR2_X1 U1069 ( .A(G902), .B(KEYINPUT48), .ZN(n1364) );
OR2_X1 U1070 ( .A1(n1176), .A2(G902), .ZN(n1361) );
XNOR2_X1 U1071 ( .A(n1365), .B(n1366), .ZN(n1176) );
XOR2_X1 U1072 ( .A(n1367), .B(n1368), .Z(n1366) );
OR2_X1 U1073 ( .A1(n1304), .A2(n1106), .ZN(n1368) );
INV_X1 U1074 ( .A(G221), .ZN(n1106) );
NAND2_X1 U1075 ( .A1(G234), .A2(n1109), .ZN(n1304) );
INV_X1 U1076 ( .A(G953), .ZN(n1109) );
NAND2_X1 U1077 ( .A1(n1369), .A2(n1370), .ZN(n1367) );
NAND2_X1 U1078 ( .A1(G110), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1079 ( .A(n1372), .B(KEYINPUT0), .Z(n1369) );
OR2_X1 U1080 ( .A1(n1371), .A2(G110), .ZN(n1372) );
XNOR2_X1 U1081 ( .A(G119), .B(n1354), .ZN(n1371) );
XOR2_X1 U1082 ( .A(n1373), .B(n1374), .Z(n1365) );
XNOR2_X1 U1083 ( .A(n1257), .B(G137), .ZN(n1374) );
INV_X1 U1084 ( .A(G146), .ZN(n1257) );
NAND2_X1 U1085 ( .A1(n1375), .A2(n1376), .ZN(n1373) );
NAND2_X1 U1086 ( .A1(G140), .A2(n1224), .ZN(n1376) );
XOR2_X1 U1087 ( .A(KEYINPUT42), .B(n1377), .Z(n1375) );
NOR2_X1 U1088 ( .A1(G140), .A2(n1224), .ZN(n1377) );
XOR2_X1 U1089 ( .A(G125), .B(KEYINPUT46), .Z(n1224) );
XNOR2_X1 U1090 ( .A(n1122), .B(G472), .ZN(n1286) );
NAND2_X1 U1091 ( .A1(n1378), .A2(n1295), .ZN(n1122) );
INV_X1 U1092 ( .A(G902), .ZN(n1295) );
XOR2_X1 U1093 ( .A(n1196), .B(n1379), .Z(n1378) );
XOR2_X1 U1094 ( .A(KEYINPUT1), .B(n1200), .Z(n1379) );
XOR2_X1 U1095 ( .A(G113), .B(n1380), .Z(n1200) );
NOR3_X1 U1096 ( .A1(KEYINPUT34), .A2(n1381), .A3(n1382), .ZN(n1380) );
NOR3_X1 U1097 ( .A1(n1383), .A2(G119), .A3(n1301), .ZN(n1382) );
INV_X1 U1098 ( .A(KEYINPUT35), .ZN(n1383) );
NOR2_X1 U1099 ( .A1(KEYINPUT35), .A2(n1325), .ZN(n1381) );
XNOR2_X1 U1100 ( .A(G119), .B(n1301), .ZN(n1325) );
XNOR2_X1 U1101 ( .A(G116), .B(KEYINPUT56), .ZN(n1301) );
XOR2_X1 U1102 ( .A(n1384), .B(n1385), .Z(n1196) );
XOR2_X1 U1103 ( .A(n1323), .B(n1347), .Z(n1385) );
XNOR2_X1 U1104 ( .A(n1150), .B(n1386), .ZN(n1347) );
XNOR2_X1 U1105 ( .A(n1157), .B(n1387), .ZN(n1386) );
NOR2_X1 U1106 ( .A1(G134), .A2(KEYINPUT21), .ZN(n1387) );
INV_X1 U1107 ( .A(G137), .ZN(n1157) );
XNOR2_X1 U1108 ( .A(G131), .B(KEYINPUT19), .ZN(n1150) );
XOR2_X1 U1109 ( .A(n1305), .B(n1388), .Z(n1323) );
NOR2_X1 U1110 ( .A1(G146), .A2(KEYINPUT25), .ZN(n1388) );
XNOR2_X1 U1111 ( .A(G143), .B(n1354), .ZN(n1305) );
INV_X1 U1112 ( .A(G128), .ZN(n1354) );
XNOR2_X1 U1113 ( .A(n1389), .B(n1332), .ZN(n1384) );
INV_X1 U1114 ( .A(G101), .ZN(n1332) );
NAND2_X1 U1115 ( .A1(n1314), .A2(G210), .ZN(n1389) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1314) );
endmodule


