//Key = 1111000011010110010010110111101011101110101001010101011110000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338;

XNOR2_X1 U719 ( .A(G107), .B(n1006), .ZN(G9) );
NAND2_X1 U720 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
XOR2_X1 U721 ( .A(n1009), .B(KEYINPUT1), .Z(n1007) );
NOR2_X1 U722 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U723 ( .A1(n1012), .A2(n1013), .A3(G953), .A4(n1014), .ZN(n1011) );
NOR2_X1 U724 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U725 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U726 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
INV_X1 U727 ( .A(n1021), .ZN(n1020) );
NOR2_X1 U728 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NOR2_X1 U729 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U730 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U731 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U732 ( .A1(n1030), .A2(n1008), .ZN(n1028) );
NOR2_X1 U733 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
XNOR2_X1 U734 ( .A(KEYINPUT36), .B(n1033), .ZN(n1031) );
NOR2_X1 U735 ( .A1(n1034), .A2(n1035), .ZN(n1026) );
NOR2_X1 U736 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U737 ( .A1(KEYINPUT7), .A2(n1038), .ZN(n1036) );
NOR3_X1 U738 ( .A1(n1029), .A2(n1039), .A3(n1035), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U740 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U741 ( .A1(n1025), .A2(n1044), .A3(n1035), .ZN(n1017) );
NOR2_X1 U742 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U743 ( .A1(n1047), .A2(n1029), .ZN(n1046) );
NOR2_X1 U744 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR3_X1 U745 ( .A1(n1050), .A2(n1021), .A3(n1038), .ZN(n1045) );
INV_X1 U746 ( .A(KEYINPUT7), .ZN(n1050) );
NOR3_X1 U747 ( .A1(n1014), .A2(G953), .A3(G952), .ZN(n1010) );
AND4_X1 U748 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1014) );
NOR4_X1 U749 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR3_X1 U750 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NOR2_X1 U751 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
AND3_X1 U752 ( .A1(n1063), .A2(n1062), .A3(KEYINPUT61), .ZN(n1060) );
AND2_X1 U753 ( .A1(KEYINPUT14), .A2(n1064), .ZN(n1062) );
NOR2_X1 U754 ( .A1(KEYINPUT61), .A2(n1064), .ZN(n1059) );
NOR2_X1 U755 ( .A1(n1065), .A2(n1066), .ZN(n1055) );
NOR2_X1 U756 ( .A1(G472), .A2(n1067), .ZN(n1066) );
XOR2_X1 U757 ( .A(n1068), .B(KEYINPUT8), .Z(n1067) );
NOR2_X1 U758 ( .A1(n1069), .A2(n1070), .ZN(n1053) );
XNOR2_X1 U759 ( .A(KEYINPUT10), .B(n1071), .ZN(n1070) );
XNOR2_X1 U760 ( .A(KEYINPUT60), .B(n1072), .ZN(n1069) );
XOR2_X1 U761 ( .A(n1073), .B(n1074), .Z(n1052) );
XNOR2_X1 U762 ( .A(n1033), .B(KEYINPUT62), .ZN(n1051) );
XOR2_X1 U763 ( .A(n1075), .B(n1076), .Z(G72) );
XOR2_X1 U764 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1077) );
XOR2_X1 U767 ( .A(KEYINPUT30), .B(n1083), .Z(n1082) );
NOR2_X1 U768 ( .A1(G900), .A2(n1079), .ZN(n1083) );
XOR2_X1 U769 ( .A(n1084), .B(n1085), .Z(n1081) );
XNOR2_X1 U770 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND2_X1 U771 ( .A1(KEYINPUT2), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U772 ( .A(KEYINPUT39), .B(n1089), .ZN(n1088) );
XOR2_X1 U773 ( .A(n1090), .B(n1091), .Z(n1084) );
XOR2_X1 U774 ( .A(G140), .B(G131), .Z(n1091) );
NAND2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
OR2_X1 U776 ( .A1(n1094), .A2(G137), .ZN(n1093) );
XOR2_X1 U777 ( .A(n1095), .B(KEYINPUT15), .Z(n1092) );
NAND2_X1 U778 ( .A1(G137), .A2(n1094), .ZN(n1095) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1079), .ZN(n1075) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1096) );
XOR2_X1 U781 ( .A(n1097), .B(n1098), .Z(G69) );
NAND2_X1 U782 ( .A1(G953), .A2(n1099), .ZN(n1098) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1099) );
NAND2_X1 U784 ( .A1(KEYINPUT49), .A2(n1100), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U787 ( .A1(G898), .A2(n1079), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1105), .A2(G953), .ZN(n1101) );
NOR2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U791 ( .A(n1110), .B(KEYINPUT46), .Z(n1109) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(G63) );
XOR2_X1 U794 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U795 ( .A1(n1111), .A2(G478), .ZN(n1115) );
NOR2_X1 U796 ( .A1(G952), .A2(n1117), .ZN(n1113) );
XNOR2_X1 U797 ( .A(KEYINPUT22), .B(n1118), .ZN(n1117) );
NOR2_X1 U798 ( .A1(n1106), .A2(n1119), .ZN(G60) );
NOR3_X1 U799 ( .A1(n1073), .A2(n1120), .A3(n1121), .ZN(n1119) );
NOR2_X1 U800 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
INV_X1 U802 ( .A(G475), .ZN(n1125) );
NOR2_X1 U803 ( .A1(n1126), .A2(n1080), .ZN(n1124) );
AND3_X1 U804 ( .A1(n1123), .A2(G475), .A3(n1111), .ZN(n1120) );
XNOR2_X1 U805 ( .A(G104), .B(n1127), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1106), .A2(n1128), .ZN(G57) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U808 ( .A(n1131), .B(n1132), .ZN(n1130) );
NAND2_X1 U809 ( .A1(KEYINPUT51), .A2(n1133), .ZN(n1131) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(n1129) );
NAND2_X1 U811 ( .A1(n1111), .A2(G472), .ZN(n1135) );
NOR2_X1 U812 ( .A1(n1106), .A2(n1136), .ZN(G54) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U814 ( .A(n1139), .B(n1087), .ZN(n1138) );
XOR2_X1 U815 ( .A(n1140), .B(n1141), .Z(n1137) );
XOR2_X1 U816 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U817 ( .A1(KEYINPUT5), .A2(n1144), .ZN(n1143) );
NOR2_X1 U818 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
NOR3_X1 U819 ( .A1(KEYINPUT48), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR2_X1 U820 ( .A1(KEYINPUT47), .A2(n1149), .ZN(n1148) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
INV_X1 U822 ( .A(KEYINPUT47), .ZN(n1151) );
NOR2_X1 U823 ( .A1(n1152), .A2(n1149), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1145) );
NOR2_X1 U825 ( .A1(n1155), .A2(n1149), .ZN(n1153) );
AND2_X1 U826 ( .A1(KEYINPUT47), .A2(KEYINPUT48), .ZN(n1155) );
NAND2_X1 U827 ( .A1(KEYINPUT27), .A2(n1156), .ZN(n1140) );
NAND2_X1 U828 ( .A1(n1111), .A2(G469), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1106), .A2(n1157), .ZN(G51) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U832 ( .A(n1162), .B(KEYINPUT24), .Z(n1158) );
NAND2_X1 U833 ( .A1(n1111), .A2(n1163), .ZN(n1162) );
XOR2_X1 U834 ( .A(KEYINPUT4), .B(n1164), .Z(n1163) );
AND2_X1 U835 ( .A1(G902), .A2(n1012), .ZN(n1111) );
NAND2_X1 U836 ( .A1(n1165), .A2(n1105), .ZN(n1012) );
INV_X1 U837 ( .A(n1126), .ZN(n1105) );
NAND4_X1 U838 ( .A1(n1166), .A2(n1127), .A3(n1167), .A4(n1168), .ZN(n1126) );
NOR2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
AND4_X1 U841 ( .A1(n1173), .A2(n1174), .A3(n1009), .A4(n1175), .ZN(n1171) );
NAND3_X1 U842 ( .A1(n1176), .A2(n1177), .A3(n1048), .ZN(n1009) );
NAND4_X1 U843 ( .A1(n1049), .A2(n1008), .A3(n1176), .A4(n1177), .ZN(n1127) );
INV_X1 U844 ( .A(n1029), .ZN(n1177) );
INV_X1 U845 ( .A(n1080), .ZN(n1165) );
NAND4_X1 U846 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1080) );
AND4_X1 U847 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NOR2_X1 U849 ( .A1(KEYINPUT16), .A2(n1188), .ZN(n1187) );
NOR3_X1 U850 ( .A1(n1189), .A2(n1190), .A3(n1035), .ZN(n1186) );
NOR2_X1 U851 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
AND4_X1 U852 ( .A1(n1041), .A2(n1037), .A3(n1193), .A4(KEYINPUT16), .ZN(n1191) );
INV_X1 U853 ( .A(n1049), .ZN(n1189) );
NAND3_X1 U854 ( .A1(n1194), .A2(n1048), .A3(n1192), .ZN(n1178) );
XNOR2_X1 U855 ( .A(n1035), .B(KEYINPUT31), .ZN(n1194) );
NOR2_X1 U856 ( .A1(n1118), .A2(G952), .ZN(n1106) );
XNOR2_X1 U857 ( .A(G953), .B(KEYINPUT43), .ZN(n1118) );
XNOR2_X1 U858 ( .A(G146), .B(n1179), .ZN(G48) );
NAND3_X1 U859 ( .A1(n1049), .A2(n1008), .A3(n1195), .ZN(n1179) );
XNOR2_X1 U860 ( .A(G143), .B(n1184), .ZN(G45) );
NAND4_X1 U861 ( .A1(n1192), .A2(n1008), .A3(n1196), .A4(n1197), .ZN(n1184) );
XNOR2_X1 U862 ( .A(G140), .B(n1188), .ZN(G42) );
NAND4_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1041), .A4(n1200), .ZN(n1188) );
AND2_X1 U864 ( .A1(n1049), .A2(n1037), .ZN(n1200) );
NAND2_X1 U865 ( .A1(n1201), .A2(n1202), .ZN(G39) );
NAND2_X1 U866 ( .A1(n1203), .A2(n1185), .ZN(n1202) );
XNOR2_X1 U867 ( .A(KEYINPUT41), .B(n1204), .ZN(n1203) );
NAND2_X1 U868 ( .A1(n1205), .A2(n1206), .ZN(n1201) );
INV_X1 U869 ( .A(n1185), .ZN(n1206) );
NAND3_X1 U870 ( .A1(n1195), .A2(n1198), .A3(n1021), .ZN(n1185) );
XNOR2_X1 U871 ( .A(G137), .B(n1207), .ZN(n1205) );
XNOR2_X1 U872 ( .A(KEYINPUT6), .B(KEYINPUT56), .ZN(n1207) );
XOR2_X1 U873 ( .A(G134), .B(n1208), .Z(G36) );
AND3_X1 U874 ( .A1(n1192), .A2(n1198), .A3(n1048), .ZN(n1208) );
XOR2_X1 U875 ( .A(G131), .B(n1209), .Z(G33) );
NOR2_X1 U876 ( .A1(n1035), .A2(n1210), .ZN(n1209) );
XOR2_X1 U877 ( .A(KEYINPUT20), .B(n1211), .Z(n1210) );
AND2_X1 U878 ( .A1(n1049), .A2(n1192), .ZN(n1211) );
NOR3_X1 U879 ( .A1(n1212), .A2(n1193), .A3(n1038), .ZN(n1192) );
INV_X1 U880 ( .A(n1198), .ZN(n1035) );
NAND2_X1 U881 ( .A1(n1213), .A2(n1214), .ZN(n1198) );
OR2_X1 U882 ( .A1(n1172), .A2(KEYINPUT36), .ZN(n1214) );
NAND3_X1 U883 ( .A1(n1215), .A2(n1032), .A3(KEYINPUT36), .ZN(n1213) );
XNOR2_X1 U884 ( .A(G128), .B(n1183), .ZN(G30) );
NAND3_X1 U885 ( .A1(n1008), .A2(n1048), .A3(n1195), .ZN(n1183) );
NOR4_X1 U886 ( .A1(n1216), .A2(n1212), .A3(n1072), .A4(n1193), .ZN(n1195) );
XOR2_X1 U887 ( .A(n1217), .B(n1169), .Z(G3) );
AND3_X1 U888 ( .A1(n1021), .A2(n1041), .A3(n1218), .ZN(n1169) );
NAND2_X1 U889 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1217) );
XOR2_X1 U890 ( .A(n1182), .B(n1219), .Z(G27) );
NAND2_X1 U891 ( .A1(n1220), .A2(KEYINPUT32), .ZN(n1219) );
XNOR2_X1 U892 ( .A(G125), .B(KEYINPUT42), .ZN(n1220) );
NAND4_X1 U893 ( .A1(n1221), .A2(n1037), .A3(n1222), .A4(n1049), .ZN(n1182) );
NOR2_X1 U894 ( .A1(n1193), .A2(n1172), .ZN(n1222) );
INV_X1 U895 ( .A(n1199), .ZN(n1193) );
NAND2_X1 U896 ( .A1(n1223), .A2(n1016), .ZN(n1199) );
NAND2_X1 U897 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
INV_X1 U898 ( .A(G900), .ZN(n1225) );
XOR2_X1 U899 ( .A(G122), .B(n1226), .Z(G24) );
NOR2_X1 U900 ( .A1(n1227), .A2(n1172), .ZN(n1226) );
XOR2_X1 U901 ( .A(n1174), .B(KEYINPUT29), .Z(n1227) );
NAND4_X1 U902 ( .A1(n1197), .A2(n1228), .A3(n1196), .A4(n1229), .ZN(n1174) );
NOR2_X1 U903 ( .A1(n1029), .A2(n1025), .ZN(n1229) );
NAND2_X1 U904 ( .A1(n1072), .A2(n1216), .ZN(n1029) );
XNOR2_X1 U905 ( .A(G119), .B(n1230), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1231), .A2(n1008), .A3(KEYINPUT28), .ZN(n1230) );
INV_X1 U907 ( .A(n1175), .ZN(n1231) );
NAND3_X1 U908 ( .A1(n1232), .A2(n1021), .A3(n1233), .ZN(n1175) );
NOR3_X1 U909 ( .A1(n1025), .A2(n1234), .A3(n1072), .ZN(n1233) );
INV_X1 U910 ( .A(n1221), .ZN(n1025) );
XNOR2_X1 U911 ( .A(G116), .B(n1167), .ZN(G18) );
NAND3_X1 U912 ( .A1(n1221), .A2(n1048), .A3(n1218), .ZN(n1167) );
NOR2_X1 U913 ( .A1(n1196), .A2(n1071), .ZN(n1048) );
INV_X1 U914 ( .A(n1197), .ZN(n1071) );
XNOR2_X1 U915 ( .A(G113), .B(n1166), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1221), .A2(n1049), .A3(n1218), .ZN(n1166) );
NOR3_X1 U917 ( .A1(n1172), .A2(n1234), .A3(n1038), .ZN(n1218) );
NAND2_X1 U918 ( .A1(n1232), .A2(n1072), .ZN(n1038) );
NOR2_X1 U919 ( .A1(n1197), .A2(n1235), .ZN(n1049) );
INV_X1 U920 ( .A(n1196), .ZN(n1235) );
NOR2_X1 U921 ( .A1(n1042), .A2(n1057), .ZN(n1221) );
XOR2_X1 U922 ( .A(G110), .B(n1236), .Z(G12) );
NOR2_X1 U923 ( .A1(n1237), .A2(n1172), .ZN(n1236) );
INV_X1 U924 ( .A(n1008), .ZN(n1172) );
NOR2_X1 U925 ( .A1(n1215), .A2(n1056), .ZN(n1008) );
INV_X1 U926 ( .A(n1032), .ZN(n1056) );
NAND2_X1 U927 ( .A1(G214), .A2(n1238), .ZN(n1032) );
INV_X1 U928 ( .A(n1033), .ZN(n1215) );
XNOR2_X1 U929 ( .A(n1239), .B(n1164), .ZN(n1033) );
AND2_X1 U930 ( .A1(G210), .A2(n1238), .ZN(n1164) );
NAND2_X1 U931 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
XNOR2_X1 U932 ( .A(G237), .B(KEYINPUT44), .ZN(n1240) );
NAND2_X1 U933 ( .A1(n1242), .A2(n1241), .ZN(n1239) );
XOR2_X1 U934 ( .A(n1243), .B(n1161), .Z(n1242) );
XNOR2_X1 U935 ( .A(n1244), .B(n1104), .ZN(n1161) );
XNOR2_X1 U936 ( .A(n1245), .B(n1246), .ZN(n1104) );
XOR2_X1 U937 ( .A(G110), .B(n1247), .Z(n1246) );
XNOR2_X1 U938 ( .A(KEYINPUT54), .B(n1248), .ZN(n1247) );
XOR2_X1 U939 ( .A(n1249), .B(n1250), .Z(n1245) );
XOR2_X1 U940 ( .A(n1251), .B(n1252), .Z(n1249) );
NAND2_X1 U941 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
NAND2_X1 U942 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U943 ( .A(KEYINPUT25), .B(n1257), .ZN(n1256) );
XNOR2_X1 U944 ( .A(KEYINPUT11), .B(G116), .ZN(n1255) );
XOR2_X1 U945 ( .A(n1258), .B(KEYINPUT58), .Z(n1253) );
NAND2_X1 U946 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U947 ( .A(KEYINPUT11), .B(G116), .Z(n1260) );
XNOR2_X1 U948 ( .A(KEYINPUT25), .B(G119), .ZN(n1259) );
NAND2_X1 U949 ( .A1(G224), .A2(n1079), .ZN(n1244) );
NOR2_X1 U950 ( .A1(n1261), .A2(n1262), .ZN(n1243) );
NOR3_X1 U951 ( .A1(n1263), .A2(n1264), .A3(n1089), .ZN(n1262) );
INV_X1 U952 ( .A(KEYINPUT50), .ZN(n1263) );
NOR2_X1 U953 ( .A1(KEYINPUT50), .A2(n1160), .ZN(n1261) );
XNOR2_X1 U954 ( .A(n1089), .B(n1264), .ZN(n1160) );
XOR2_X1 U955 ( .A(n1173), .B(KEYINPUT57), .Z(n1237) );
NAND3_X1 U956 ( .A1(n1037), .A2(n1176), .A3(n1021), .ZN(n1173) );
NOR2_X1 U957 ( .A1(n1197), .A2(n1196), .ZN(n1021) );
XNOR2_X1 U958 ( .A(n1265), .B(n1266), .ZN(n1196) );
XOR2_X1 U959 ( .A(KEYINPUT23), .B(n1073), .Z(n1266) );
NOR2_X1 U960 ( .A1(n1123), .A2(G902), .ZN(n1073) );
XNOR2_X1 U961 ( .A(n1267), .B(n1268), .ZN(n1123) );
XOR2_X1 U962 ( .A(G122), .B(n1269), .Z(n1268) );
XOR2_X1 U963 ( .A(G143), .B(G131), .Z(n1269) );
XOR2_X1 U964 ( .A(n1270), .B(G104), .Z(n1267) );
NAND2_X1 U965 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U966 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
INV_X1 U967 ( .A(n1275), .ZN(n1274) );
XOR2_X1 U968 ( .A(KEYINPUT33), .B(n1276), .Z(n1273) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1275), .ZN(n1271) );
XOR2_X1 U970 ( .A(G125), .B(n1278), .Z(n1275) );
XNOR2_X1 U971 ( .A(n1279), .B(G140), .ZN(n1278) );
XOR2_X1 U972 ( .A(KEYINPUT35), .B(n1276), .Z(n1277) );
XNOR2_X1 U973 ( .A(n1280), .B(n1281), .ZN(n1276) );
AND3_X1 U974 ( .A1(G214), .A2(n1079), .A3(n1282), .ZN(n1281) );
NAND2_X1 U975 ( .A1(KEYINPUT34), .A2(n1248), .ZN(n1280) );
INV_X1 U976 ( .A(G113), .ZN(n1248) );
NAND2_X1 U977 ( .A1(KEYINPUT0), .A2(n1074), .ZN(n1265) );
XOR2_X1 U978 ( .A(G475), .B(KEYINPUT63), .Z(n1074) );
XNOR2_X1 U979 ( .A(n1283), .B(G478), .ZN(n1197) );
NAND2_X1 U980 ( .A1(n1116), .A2(n1241), .ZN(n1283) );
XOR2_X1 U981 ( .A(n1284), .B(n1285), .Z(n1116) );
XOR2_X1 U982 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U983 ( .A(G134), .B(n1288), .ZN(n1287) );
XOR2_X1 U984 ( .A(KEYINPUT9), .B(G143), .Z(n1286) );
XOR2_X1 U985 ( .A(n1289), .B(n1250), .Z(n1284) );
XNOR2_X1 U986 ( .A(n1290), .B(G122), .ZN(n1250) );
INV_X1 U987 ( .A(G107), .ZN(n1290) );
XOR2_X1 U988 ( .A(n1291), .B(G116), .Z(n1289) );
NAND2_X1 U989 ( .A1(G217), .A2(n1292), .ZN(n1291) );
NOR2_X1 U990 ( .A1(n1212), .A2(n1234), .ZN(n1176) );
INV_X1 U991 ( .A(n1228), .ZN(n1234) );
NAND2_X1 U992 ( .A1(n1293), .A2(n1016), .ZN(n1228) );
NAND3_X1 U993 ( .A1(n1294), .A2(n1079), .A3(G952), .ZN(n1016) );
NAND2_X1 U994 ( .A1(n1224), .A2(n1295), .ZN(n1293) );
INV_X1 U995 ( .A(G898), .ZN(n1295) );
AND3_X1 U996 ( .A1(G902), .A2(n1294), .A3(G953), .ZN(n1224) );
NAND2_X1 U997 ( .A1(G234), .A2(G237), .ZN(n1294) );
INV_X1 U998 ( .A(n1041), .ZN(n1212) );
NOR2_X1 U999 ( .A1(n1296), .A2(n1057), .ZN(n1041) );
INV_X1 U1000 ( .A(n1043), .ZN(n1057) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1297), .ZN(n1043) );
INV_X1 U1002 ( .A(n1042), .ZN(n1296) );
XOR2_X1 U1003 ( .A(n1064), .B(n1063), .Z(n1042) );
INV_X1 U1004 ( .A(G469), .ZN(n1063) );
NAND2_X1 U1005 ( .A1(n1298), .A2(n1241), .ZN(n1064) );
XOR2_X1 U1006 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1007 ( .A(n1301), .B(n1302), .ZN(n1300) );
NOR2_X1 U1008 ( .A1(KEYINPUT18), .A2(n1139), .ZN(n1302) );
NAND3_X1 U1009 ( .A1(n1303), .A2(n1304), .A3(KEYINPUT26), .ZN(n1301) );
NAND2_X1 U1010 ( .A1(KEYINPUT40), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U1011 ( .A(n1154), .B(n1149), .ZN(n1305) );
OR3_X1 U1012 ( .A1(n1149), .A2(n1152), .A3(KEYINPUT40), .ZN(n1303) );
INV_X1 U1013 ( .A(n1154), .ZN(n1152) );
NAND2_X1 U1014 ( .A1(G227), .A2(n1079), .ZN(n1154) );
XNOR2_X1 U1015 ( .A(G110), .B(G140), .ZN(n1149) );
XNOR2_X1 U1016 ( .A(n1144), .B(n1087), .ZN(n1299) );
XOR2_X1 U1017 ( .A(G128), .B(n1306), .Z(n1087) );
NOR2_X1 U1018 ( .A1(KEYINPUT52), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1019 ( .A(n1308), .B(n1252), .ZN(n1144) );
XNOR2_X1 U1020 ( .A(G104), .B(n1133), .ZN(n1252) );
INV_X1 U1021 ( .A(G101), .ZN(n1133) );
XNOR2_X1 U1022 ( .A(G107), .B(KEYINPUT59), .ZN(n1308) );
NOR2_X1 U1023 ( .A1(n1232), .A2(n1072), .ZN(n1037) );
XOR2_X1 U1024 ( .A(n1309), .B(n1112), .Z(n1072) );
AND2_X1 U1025 ( .A1(G217), .A2(n1297), .ZN(n1112) );
NAND2_X1 U1026 ( .A1(G234), .A2(n1241), .ZN(n1297) );
NAND2_X1 U1027 ( .A1(n1108), .A2(n1241), .ZN(n1309) );
XOR2_X1 U1028 ( .A(n1310), .B(n1311), .Z(n1108) );
XNOR2_X1 U1029 ( .A(KEYINPUT53), .B(n1204), .ZN(n1311) );
INV_X1 U1030 ( .A(G137), .ZN(n1204) );
XOR2_X1 U1031 ( .A(n1312), .B(n1313), .Z(n1310) );
XOR2_X1 U1032 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1033 ( .A(n1089), .B(G119), .ZN(n1315) );
INV_X1 U1034 ( .A(G125), .ZN(n1089) );
XNOR2_X1 U1035 ( .A(KEYINPUT13), .B(n1288), .ZN(n1314) );
XOR2_X1 U1036 ( .A(n1316), .B(n1317), .Z(n1312) );
XNOR2_X1 U1037 ( .A(G110), .B(n1318), .ZN(n1317) );
NAND2_X1 U1038 ( .A1(KEYINPUT38), .A2(n1279), .ZN(n1318) );
XNOR2_X1 U1039 ( .A(n1319), .B(n1320), .ZN(n1316) );
NAND2_X1 U1040 ( .A1(KEYINPUT55), .A2(G140), .ZN(n1320) );
NAND3_X1 U1041 ( .A1(G221), .A2(n1292), .A3(KEYINPUT37), .ZN(n1319) );
AND2_X1 U1042 ( .A1(G234), .A2(n1079), .ZN(n1292) );
INV_X1 U1043 ( .A(n1216), .ZN(n1232) );
NAND2_X1 U1044 ( .A1(n1321), .A2(n1322), .ZN(n1216) );
NAND2_X1 U1045 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
INV_X1 U1046 ( .A(KEYINPUT21), .ZN(n1324) );
NAND2_X1 U1047 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND2_X1 U1048 ( .A1(n1068), .A2(n1327), .ZN(n1326) );
INV_X1 U1049 ( .A(n1065), .ZN(n1325) );
NOR2_X1 U1050 ( .A1(n1068), .A2(n1327), .ZN(n1065) );
INV_X1 U1051 ( .A(G472), .ZN(n1327) );
NAND2_X1 U1052 ( .A1(n1328), .A2(KEYINPUT21), .ZN(n1321) );
XNOR2_X1 U1053 ( .A(G472), .B(n1068), .ZN(n1328) );
NAND2_X1 U1054 ( .A1(n1329), .A2(n1241), .ZN(n1068) );
INV_X1 U1055 ( .A(G902), .ZN(n1241) );
XNOR2_X1 U1056 ( .A(n1330), .B(n1331), .ZN(n1329) );
INV_X1 U1057 ( .A(n1132), .ZN(n1331) );
XNOR2_X1 U1058 ( .A(n1332), .B(n1333), .ZN(n1132) );
XNOR2_X1 U1059 ( .A(n1264), .B(n1139), .ZN(n1333) );
XOR2_X1 U1060 ( .A(n1334), .B(n1335), .Z(n1139) );
NOR2_X1 U1061 ( .A1(KEYINPUT12), .A2(n1094), .ZN(n1335) );
XOR2_X1 U1062 ( .A(G134), .B(KEYINPUT17), .Z(n1094) );
XNOR2_X1 U1063 ( .A(G131), .B(G137), .ZN(n1334) );
XOR2_X1 U1064 ( .A(n1336), .B(n1288), .Z(n1264) );
INV_X1 U1065 ( .A(G128), .ZN(n1288) );
NAND2_X1 U1066 ( .A1(KEYINPUT3), .A2(n1307), .ZN(n1336) );
XNOR2_X1 U1067 ( .A(G143), .B(n1279), .ZN(n1307) );
INV_X1 U1068 ( .A(G146), .ZN(n1279) );
XNOR2_X1 U1069 ( .A(G113), .B(n1337), .ZN(n1332) );
XNOR2_X1 U1070 ( .A(n1257), .B(G116), .ZN(n1337) );
INV_X1 U1071 ( .A(G119), .ZN(n1257) );
XOR2_X1 U1072 ( .A(n1134), .B(n1338), .Z(n1330) );
NOR2_X1 U1073 ( .A1(G101), .A2(KEYINPUT19), .ZN(n1338) );
NAND3_X1 U1074 ( .A1(n1282), .A2(n1079), .A3(G210), .ZN(n1134) );
INV_X1 U1075 ( .A(G953), .ZN(n1079) );
INV_X1 U1076 ( .A(G237), .ZN(n1282) );
endmodule


