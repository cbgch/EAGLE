//Key = 0110000010100110001010001000111010010100100010000110010010111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408;

XOR2_X1 U755 ( .A(n1056), .B(n1057), .Z(G9) );
NOR2_X1 U756 ( .A1(KEYINPUT52), .A2(n1058), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR3_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR3_X1 U759 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NAND3_X1 U761 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1061) );
NAND3_X1 U762 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U765 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
OR2_X1 U766 ( .A1(n1066), .A2(KEYINPUT50), .ZN(n1080) );
NAND3_X1 U767 ( .A1(n1082), .A2(n1083), .A3(KEYINPUT50), .ZN(n1079) );
INV_X1 U768 ( .A(n1064), .ZN(n1077) );
NAND3_X1 U769 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1064) );
NAND3_X1 U770 ( .A1(n1087), .A2(n1088), .A3(n1086), .ZN(n1075) );
INV_X1 U771 ( .A(n1089), .ZN(n1086) );
NAND3_X1 U772 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1093), .ZN(n1092) );
NAND2_X1 U774 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND3_X1 U775 ( .A1(n1084), .A2(n1096), .A3(n1097), .ZN(n1090) );
NOR3_X1 U776 ( .A1(n1098), .A2(G953), .A3(G952), .ZN(n1059) );
INV_X1 U777 ( .A(n1069), .ZN(n1098) );
NAND4_X1 U778 ( .A1(n1074), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1069) );
NOR3_X1 U779 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
XNOR2_X1 U780 ( .A(n1105), .B(KEYINPUT49), .ZN(n1104) );
NOR2_X1 U781 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND3_X1 U782 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1102) );
NAND2_X1 U783 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND4_X1 U784 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1111) );
NAND2_X1 U785 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U786 ( .A1(G469), .A2(n1119), .ZN(n1118) );
NAND2_X1 U787 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U788 ( .A1(n1122), .A2(n1123), .ZN(n1114) );
NAND2_X1 U789 ( .A1(n1124), .A2(n1107), .ZN(n1113) );
NOR4_X1 U790 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1100) );
NOR2_X1 U791 ( .A1(G469), .A2(n1119), .ZN(n1128) );
INV_X1 U792 ( .A(KEYINPUT27), .ZN(n1119) );
NOR3_X1 U793 ( .A1(KEYINPUT27), .A2(n1129), .A3(n1130), .ZN(n1127) );
INV_X1 U794 ( .A(G469), .ZN(n1130) );
AND3_X1 U795 ( .A1(KEYINPUT28), .A2(n1131), .A3(n1132), .ZN(n1126) );
NOR2_X1 U796 ( .A1(KEYINPUT28), .A2(n1132), .ZN(n1125) );
XNOR2_X1 U797 ( .A(KEYINPUT32), .B(n1133), .ZN(n1099) );
XOR2_X1 U798 ( .A(n1134), .B(n1135), .Z(G72) );
NOR2_X1 U799 ( .A1(n1136), .A2(n1070), .ZN(n1135) );
AND2_X1 U800 ( .A1(G227), .A2(G900), .ZN(n1136) );
NAND2_X1 U801 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND3_X1 U802 ( .A1(n1139), .A2(n1070), .A3(n1140), .ZN(n1138) );
INV_X1 U803 ( .A(n1141), .ZN(n1140) );
NAND3_X1 U804 ( .A1(n1142), .A2(n1143), .A3(n1141), .ZN(n1137) );
XNOR2_X1 U805 ( .A(n1144), .B(n1145), .ZN(n1141) );
XNOR2_X1 U806 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U807 ( .A1(KEYINPUT22), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U808 ( .A(KEYINPUT21), .B(n1149), .ZN(n1148) );
INV_X1 U809 ( .A(G125), .ZN(n1146) );
NAND2_X1 U810 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U811 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U812 ( .A(KEYINPUT2), .B(n1154), .Z(n1150) );
NOR2_X1 U813 ( .A1(n1152), .A2(n1153), .ZN(n1154) );
XNOR2_X1 U814 ( .A(n1155), .B(n1156), .ZN(n1153) );
NOR2_X1 U815 ( .A1(KEYINPUT26), .A2(n1157), .ZN(n1156) );
XOR2_X1 U816 ( .A(G137), .B(n1158), .Z(n1157) );
NOR2_X1 U817 ( .A1(KEYINPUT6), .A2(n1159), .ZN(n1158) );
XNOR2_X1 U818 ( .A(KEYINPUT51), .B(n1139), .ZN(n1142) );
XOR2_X1 U819 ( .A(n1160), .B(n1161), .Z(G69) );
NOR2_X1 U820 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U821 ( .A(n1164), .B(KEYINPUT37), .Z(n1163) );
NAND2_X1 U822 ( .A1(G953), .A2(n1165), .ZN(n1164) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1165) );
NOR2_X1 U824 ( .A1(n1166), .A2(G953), .ZN(n1162) );
NOR2_X1 U825 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U826 ( .A(KEYINPUT25), .B(n1169), .Z(n1168) );
NAND2_X1 U827 ( .A1(n1170), .A2(n1171), .ZN(n1160) );
NAND2_X1 U828 ( .A1(n1172), .A2(G953), .ZN(n1171) );
XOR2_X1 U829 ( .A(n1173), .B(n1174), .Z(n1170) );
XOR2_X1 U830 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U831 ( .A(KEYINPUT61), .B(KEYINPUT56), .Z(n1176) );
XOR2_X1 U832 ( .A(n1177), .B(n1178), .Z(n1173) );
NOR2_X1 U833 ( .A1(n1179), .A2(n1180), .ZN(G66) );
XOR2_X1 U834 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U835 ( .A1(n1107), .A2(n1183), .ZN(n1182) );
NAND2_X1 U836 ( .A1(KEYINPUT44), .A2(n1124), .ZN(n1181) );
NOR2_X1 U837 ( .A1(n1179), .A2(n1184), .ZN(G63) );
XOR2_X1 U838 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U839 ( .A1(n1123), .A2(n1183), .ZN(n1186) );
NAND2_X1 U840 ( .A1(KEYINPUT10), .A2(n1122), .ZN(n1185) );
NOR2_X1 U841 ( .A1(n1179), .A2(n1187), .ZN(G60) );
XOR2_X1 U842 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U843 ( .A1(n1190), .A2(G475), .ZN(n1188) );
XOR2_X1 U844 ( .A(G104), .B(n1169), .Z(G6) );
NOR2_X1 U845 ( .A1(n1179), .A2(n1191), .ZN(G57) );
XOR2_X1 U846 ( .A(n1192), .B(n1193), .Z(n1191) );
NAND2_X1 U847 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NAND4_X1 U848 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
NOR2_X1 U849 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XNOR2_X1 U850 ( .A(n1202), .B(n1203), .ZN(n1196) );
NAND2_X1 U851 ( .A1(n1204), .A2(n1205), .ZN(n1194) );
NAND2_X1 U852 ( .A1(n1198), .A2(n1197), .ZN(n1205) );
XNOR2_X1 U853 ( .A(KEYINPUT8), .B(n1206), .ZN(n1198) );
NAND3_X1 U854 ( .A1(n1207), .A2(n1208), .A3(G472), .ZN(n1204) );
NAND2_X1 U855 ( .A1(KEYINPUT58), .A2(n1183), .ZN(n1208) );
INV_X1 U856 ( .A(n1190), .ZN(n1183) );
NAND2_X1 U857 ( .A1(n1209), .A2(n1202), .ZN(n1207) );
INV_X1 U858 ( .A(KEYINPUT58), .ZN(n1202) );
OR2_X1 U859 ( .A1(n1201), .A2(n1063), .ZN(n1209) );
INV_X1 U860 ( .A(n1203), .ZN(n1063) );
NOR2_X1 U861 ( .A1(n1179), .A2(n1210), .ZN(G54) );
XOR2_X1 U862 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U863 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR3_X1 U864 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
NOR3_X1 U865 ( .A1(G140), .A2(G110), .A3(n1218), .ZN(n1217) );
NOR2_X1 U866 ( .A1(n1149), .A2(n1219), .ZN(n1216) );
XNOR2_X1 U867 ( .A(n1218), .B(n1220), .ZN(n1219) );
XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n1221), .ZN(n1220) );
NAND2_X1 U869 ( .A1(n1222), .A2(n1223), .ZN(n1213) );
NAND2_X1 U870 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U871 ( .A(KEYINPUT1), .B(n1226), .Z(n1222) );
NOR2_X1 U872 ( .A1(n1224), .A2(n1225), .ZN(n1226) );
XNOR2_X1 U873 ( .A(n1227), .B(n1228), .ZN(n1224) );
NAND2_X1 U874 ( .A1(n1190), .A2(G469), .ZN(n1211) );
NOR2_X1 U875 ( .A1(n1179), .A2(n1229), .ZN(G51) );
XOR2_X1 U876 ( .A(n1230), .B(n1120), .Z(n1229) );
XOR2_X1 U877 ( .A(n1231), .B(KEYINPUT17), .Z(n1230) );
NAND2_X1 U878 ( .A1(n1190), .A2(n1132), .ZN(n1231) );
INV_X1 U879 ( .A(n1121), .ZN(n1132) );
NOR2_X1 U880 ( .A1(n1201), .A2(n1203), .ZN(n1190) );
NOR3_X1 U881 ( .A1(n1167), .A2(n1169), .A3(n1139), .ZN(n1203) );
NAND4_X1 U882 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1139) );
AND4_X1 U883 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NAND2_X1 U884 ( .A1(n1067), .A2(n1240), .ZN(n1234) );
NAND2_X1 U885 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND3_X1 U886 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1242) );
OR2_X1 U887 ( .A1(n1246), .A2(KEYINPUT41), .ZN(n1244) );
NAND2_X1 U888 ( .A1(KEYINPUT41), .A2(n1247), .ZN(n1243) );
NAND2_X1 U889 ( .A1(n1248), .A2(n1066), .ZN(n1247) );
INV_X1 U890 ( .A(n1087), .ZN(n1066) );
NAND2_X1 U891 ( .A1(n1249), .A2(n1250), .ZN(n1241) );
NAND3_X1 U892 ( .A1(n1084), .A2(n1246), .A3(n1251), .ZN(n1233) );
XNOR2_X1 U893 ( .A(n1252), .B(KEYINPUT13), .ZN(n1251) );
NAND3_X1 U894 ( .A1(n1250), .A2(n1245), .A3(n1252), .ZN(n1232) );
AND3_X1 U895 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1169) );
NAND4_X1 U896 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1167) );
NOR4_X1 U897 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1056), .ZN(n1259) );
AND3_X1 U898 ( .A1(n1253), .A2(n1254), .A3(n1245), .ZN(n1056) );
NAND2_X1 U899 ( .A1(n1263), .A2(n1085), .ZN(n1258) );
NAND3_X1 U900 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1257) );
XNOR2_X1 U901 ( .A(n1267), .B(KEYINPUT53), .ZN(n1266) );
NAND2_X1 U902 ( .A1(n1268), .A2(n1267), .ZN(n1256) );
XOR2_X1 U903 ( .A(n1269), .B(KEYINPUT29), .Z(n1268) );
XOR2_X1 U904 ( .A(G902), .B(KEYINPUT14), .Z(n1201) );
NOR2_X1 U905 ( .A1(n1070), .A2(G952), .ZN(n1179) );
XNOR2_X1 U906 ( .A(G146), .B(n1239), .ZN(G48) );
NAND3_X1 U907 ( .A1(n1250), .A2(n1255), .A3(n1252), .ZN(n1239) );
INV_X1 U908 ( .A(n1270), .ZN(n1250) );
XOR2_X1 U909 ( .A(G143), .B(n1271), .Z(G45) );
NOR4_X1 U910 ( .A1(KEYINPUT4), .A2(n1272), .A3(n1270), .A4(n1273), .ZN(n1271) );
XNOR2_X1 U911 ( .A(G140), .B(n1238), .ZN(G42) );
NAND3_X1 U912 ( .A1(n1068), .A2(n1255), .A3(n1246), .ZN(n1238) );
INV_X1 U913 ( .A(n1274), .ZN(n1246) );
XOR2_X1 U914 ( .A(G137), .B(n1275), .Z(G39) );
NOR2_X1 U915 ( .A1(n1274), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U916 ( .A(G134), .B(n1277), .ZN(G36) );
NAND2_X1 U917 ( .A1(n1278), .A2(n1245), .ZN(n1277) );
XNOR2_X1 U918 ( .A(G131), .B(n1237), .ZN(G33) );
NAND2_X1 U919 ( .A1(n1278), .A2(n1255), .ZN(n1237) );
NOR2_X1 U920 ( .A1(n1274), .A2(n1272), .ZN(n1278) );
NAND2_X1 U921 ( .A1(n1248), .A2(n1087), .ZN(n1274) );
NOR2_X1 U922 ( .A1(n1279), .A2(n1082), .ZN(n1087) );
XNOR2_X1 U923 ( .A(n1280), .B(n1281), .ZN(G30) );
NOR3_X1 U924 ( .A1(n1270), .A2(n1282), .A3(n1094), .ZN(n1281) );
XNOR2_X1 U925 ( .A(n1252), .B(KEYINPUT15), .ZN(n1282) );
NAND2_X1 U926 ( .A1(n1248), .A2(n1267), .ZN(n1270) );
AND2_X1 U927 ( .A1(n1253), .A2(n1283), .ZN(n1248) );
XOR2_X1 U928 ( .A(G101), .B(n1284), .Z(G3) );
NOR2_X1 U929 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
INV_X1 U930 ( .A(n1264), .ZN(n1286) );
NOR2_X1 U931 ( .A1(n1091), .A2(n1272), .ZN(n1264) );
XNOR2_X1 U932 ( .A(G125), .B(n1236), .ZN(G27) );
NAND4_X1 U933 ( .A1(n1085), .A2(n1068), .A3(n1287), .A4(n1255), .ZN(n1236) );
INV_X1 U934 ( .A(n1095), .ZN(n1255) );
AND2_X1 U935 ( .A1(n1283), .A2(n1267), .ZN(n1287) );
NAND2_X1 U936 ( .A1(n1089), .A2(n1288), .ZN(n1283) );
NAND3_X1 U937 ( .A1(G902), .A2(n1289), .A3(n1290), .ZN(n1288) );
INV_X1 U938 ( .A(n1143), .ZN(n1290) );
NAND2_X1 U939 ( .A1(n1291), .A2(G953), .ZN(n1143) );
XNOR2_X1 U940 ( .A(G900), .B(KEYINPUT46), .ZN(n1291) );
INV_X1 U941 ( .A(n1292), .ZN(n1068) );
XOR2_X1 U942 ( .A(G122), .B(n1262), .Z(G24) );
AND3_X1 U943 ( .A1(n1085), .A2(n1254), .A3(n1249), .ZN(n1262) );
INV_X1 U944 ( .A(n1273), .ZN(n1249) );
NAND2_X1 U945 ( .A1(n1105), .A2(n1293), .ZN(n1273) );
NOR3_X1 U946 ( .A1(n1294), .A2(n1295), .A3(n1285), .ZN(n1254) );
XNOR2_X1 U947 ( .A(n1296), .B(n1297), .ZN(G21) );
NOR2_X1 U948 ( .A1(n1081), .A2(n1269), .ZN(n1297) );
NAND3_X1 U949 ( .A1(n1085), .A2(n1265), .A3(n1298), .ZN(n1269) );
INV_X1 U950 ( .A(n1276), .ZN(n1298) );
NAND2_X1 U951 ( .A1(n1084), .A2(n1252), .ZN(n1276) );
NOR2_X1 U952 ( .A1(n1072), .A2(n1074), .ZN(n1252) );
INV_X1 U953 ( .A(n1299), .ZN(n1085) );
INV_X1 U954 ( .A(n1267), .ZN(n1081) );
XNOR2_X1 U955 ( .A(n1261), .B(n1300), .ZN(G18) );
NOR2_X1 U956 ( .A1(G116), .A2(KEYINPUT39), .ZN(n1300) );
NOR4_X1 U957 ( .A1(n1272), .A2(n1299), .A3(n1094), .A4(n1285), .ZN(n1261) );
INV_X1 U958 ( .A(n1245), .ZN(n1094) );
NOR2_X1 U959 ( .A1(n1105), .A2(n1301), .ZN(n1245) );
NAND2_X1 U960 ( .A1(n1302), .A2(n1303), .ZN(G15) );
NAND2_X1 U961 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U962 ( .A(KEYINPUT63), .B(n1306), .Z(n1302) );
NOR2_X1 U963 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
AND2_X1 U964 ( .A1(n1263), .A2(n1307), .ZN(n1304) );
XNOR2_X1 U965 ( .A(KEYINPUT42), .B(n1299), .ZN(n1307) );
NAND2_X1 U966 ( .A1(n1096), .A2(n1109), .ZN(n1299) );
NOR3_X1 U967 ( .A1(n1095), .A2(n1285), .A3(n1272), .ZN(n1263) );
INV_X1 U968 ( .A(n1067), .ZN(n1272) );
NOR2_X1 U969 ( .A1(n1074), .A2(n1295), .ZN(n1067) );
INV_X1 U970 ( .A(n1072), .ZN(n1295) );
NAND2_X1 U971 ( .A1(n1301), .A2(n1105), .ZN(n1095) );
INV_X1 U972 ( .A(n1293), .ZN(n1301) );
XNOR2_X1 U973 ( .A(n1221), .B(n1260), .ZN(G12) );
NOR3_X1 U974 ( .A1(n1292), .A2(n1285), .A3(n1091), .ZN(n1260) );
NAND2_X1 U975 ( .A1(n1084), .A2(n1253), .ZN(n1091) );
NOR2_X1 U976 ( .A1(n1096), .A2(n1097), .ZN(n1253) );
INV_X1 U977 ( .A(n1109), .ZN(n1097) );
NAND2_X1 U978 ( .A1(G221), .A2(n1308), .ZN(n1109) );
XOR2_X1 U979 ( .A(G469), .B(n1309), .Z(n1096) );
NOR2_X1 U980 ( .A1(n1129), .A2(KEYINPUT45), .ZN(n1309) );
AND2_X1 U981 ( .A1(n1117), .A2(n1112), .ZN(n1129) );
XNOR2_X1 U982 ( .A(n1310), .B(n1311), .ZN(n1117) );
XOR2_X1 U983 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR3_X1 U984 ( .A1(n1215), .A2(n1314), .A3(n1315), .ZN(n1313) );
NOR3_X1 U985 ( .A1(n1221), .A2(n1149), .A3(n1218), .ZN(n1315) );
NOR2_X1 U986 ( .A1(G110), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U987 ( .A(n1317), .B(n1318), .ZN(n1316) );
XNOR2_X1 U988 ( .A(KEYINPUT19), .B(n1149), .ZN(n1318) );
NOR3_X1 U989 ( .A1(n1317), .A2(G140), .A3(n1221), .ZN(n1215) );
INV_X1 U990 ( .A(n1218), .ZN(n1317) );
NAND2_X1 U991 ( .A1(G227), .A2(n1070), .ZN(n1218) );
NOR4_X1 U992 ( .A1(n1319), .A2(n1320), .A3(KEYINPUT47), .A4(n1321), .ZN(n1312) );
NOR2_X1 U993 ( .A1(n1322), .A2(n1227), .ZN(n1321) );
NOR2_X1 U994 ( .A1(n1152), .A2(n1323), .ZN(n1322) );
AND2_X1 U995 ( .A1(n1152), .A2(KEYINPUT62), .ZN(n1320) );
NOR4_X1 U996 ( .A1(KEYINPUT62), .A2(n1324), .A3(n1152), .A4(n1323), .ZN(n1319) );
XNOR2_X1 U997 ( .A(KEYINPUT23), .B(KEYINPUT20), .ZN(n1323) );
INV_X1 U998 ( .A(n1227), .ZN(n1324) );
XNOR2_X1 U999 ( .A(n1325), .B(n1326), .ZN(n1227) );
XNOR2_X1 U1000 ( .A(G101), .B(G107), .ZN(n1325) );
INV_X1 U1001 ( .A(n1225), .ZN(n1310) );
NOR2_X1 U1002 ( .A1(n1293), .A2(n1105), .ZN(n1084) );
XNOR2_X1 U1003 ( .A(n1327), .B(G475), .ZN(n1105) );
NAND2_X1 U1004 ( .A1(n1328), .A2(n1112), .ZN(n1327) );
XNOR2_X1 U1005 ( .A(n1189), .B(KEYINPUT40), .ZN(n1328) );
XNOR2_X1 U1006 ( .A(n1329), .B(n1330), .ZN(n1189) );
XNOR2_X1 U1007 ( .A(G122), .B(n1305), .ZN(n1330) );
INV_X1 U1008 ( .A(G113), .ZN(n1305) );
XOR2_X1 U1009 ( .A(n1331), .B(n1326), .Z(n1329) );
NAND2_X1 U1010 ( .A1(KEYINPUT59), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1011 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1012 ( .A(n1335), .B(n1336), .ZN(n1334) );
XOR2_X1 U1013 ( .A(n1337), .B(n1338), .Z(n1333) );
XNOR2_X1 U1014 ( .A(KEYINPUT24), .B(n1155), .ZN(n1338) );
INV_X1 U1015 ( .A(G131), .ZN(n1155) );
NAND2_X1 U1016 ( .A1(G214), .A2(n1339), .ZN(n1337) );
NAND2_X1 U1017 ( .A1(n1133), .A2(n1340), .ZN(n1293) );
NAND3_X1 U1018 ( .A1(n1123), .A2(n1112), .A3(n1122), .ZN(n1340) );
INV_X1 U1019 ( .A(G478), .ZN(n1123) );
NAND2_X1 U1020 ( .A1(G478), .A2(n1341), .ZN(n1133) );
NAND2_X1 U1021 ( .A1(n1122), .A2(n1112), .ZN(n1341) );
XOR2_X1 U1022 ( .A(n1342), .B(n1343), .Z(n1122) );
XOR2_X1 U1023 ( .A(n1344), .B(n1345), .Z(n1343) );
NOR2_X1 U1024 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NOR2_X1 U1025 ( .A1(KEYINPUT33), .A2(n1348), .ZN(n1347) );
AND2_X1 U1026 ( .A1(KEYINPUT7), .A2(n1348), .ZN(n1346) );
AND3_X1 U1027 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1348) );
NAND2_X1 U1028 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1029 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XNOR2_X1 U1030 ( .A(G116), .B(G122), .ZN(n1352) );
NAND4_X1 U1031 ( .A1(n1354), .A2(n1355), .A3(n1356), .A4(n1357), .ZN(n1350) );
XNOR2_X1 U1032 ( .A(G122), .B(n1358), .ZN(n1356) );
INV_X1 U1033 ( .A(G116), .ZN(n1358) );
INV_X1 U1034 ( .A(KEYINPUT38), .ZN(n1355) );
OR2_X1 U1035 ( .A1(n1357), .A2(n1354), .ZN(n1349) );
XOR2_X1 U1036 ( .A(G107), .B(KEYINPUT60), .Z(n1354) );
INV_X1 U1037 ( .A(KEYINPUT12), .ZN(n1357) );
AND2_X1 U1038 ( .A1(n1359), .A2(G217), .ZN(n1344) );
XNOR2_X1 U1039 ( .A(G128), .B(n1360), .ZN(n1342) );
XNOR2_X1 U1040 ( .A(G143), .B(n1159), .ZN(n1360) );
INV_X1 U1041 ( .A(G134), .ZN(n1159) );
NAND2_X1 U1042 ( .A1(n1267), .A2(n1265), .ZN(n1285) );
NAND2_X1 U1043 ( .A1(n1361), .A2(n1089), .ZN(n1265) );
NAND3_X1 U1044 ( .A1(n1289), .A2(n1070), .A3(G952), .ZN(n1089) );
NAND4_X1 U1045 ( .A1(n1172), .A2(n1362), .A3(G902), .A4(G953), .ZN(n1361) );
XOR2_X1 U1046 ( .A(n1289), .B(KEYINPUT57), .Z(n1362) );
NAND2_X1 U1047 ( .A1(G237), .A2(G234), .ZN(n1289) );
XNOR2_X1 U1048 ( .A(G898), .B(KEYINPUT43), .ZN(n1172) );
NOR2_X1 U1049 ( .A1(n1083), .A2(n1082), .ZN(n1267) );
INV_X1 U1050 ( .A(n1108), .ZN(n1082) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1363), .ZN(n1108) );
INV_X1 U1052 ( .A(n1279), .ZN(n1083) );
XOR2_X1 U1053 ( .A(n1131), .B(n1121), .Z(n1279) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1363), .ZN(n1121) );
NAND2_X1 U1055 ( .A1(n1364), .A2(n1112), .ZN(n1363) );
INV_X1 U1056 ( .A(G237), .ZN(n1364) );
NAND2_X1 U1057 ( .A1(n1120), .A2(n1112), .ZN(n1131) );
XNOR2_X1 U1058 ( .A(n1365), .B(n1366), .ZN(n1120) );
XOR2_X1 U1059 ( .A(n1367), .B(n1368), .Z(n1366) );
XNOR2_X1 U1060 ( .A(G125), .B(n1369), .ZN(n1368) );
NOR2_X1 U1061 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XNOR2_X1 U1062 ( .A(KEYINPUT0), .B(n1070), .ZN(n1371) );
INV_X1 U1063 ( .A(G224), .ZN(n1370) );
NAND2_X1 U1064 ( .A1(n1372), .A2(n1373), .ZN(n1367) );
NAND2_X1 U1065 ( .A1(n1177), .A2(n1175), .ZN(n1373) );
XOR2_X1 U1066 ( .A(n1374), .B(KEYINPUT11), .Z(n1372) );
OR2_X1 U1067 ( .A1(n1175), .A2(n1177), .ZN(n1374) );
XOR2_X1 U1068 ( .A(n1375), .B(n1376), .Z(n1177) );
XOR2_X1 U1069 ( .A(KEYINPUT16), .B(G101), .Z(n1376) );
NAND2_X1 U1070 ( .A1(n1377), .A2(KEYINPUT35), .ZN(n1375) );
XNOR2_X1 U1071 ( .A(n1378), .B(n1058), .ZN(n1377) );
INV_X1 U1072 ( .A(G107), .ZN(n1058) );
NAND2_X1 U1073 ( .A1(KEYINPUT30), .A2(n1326), .ZN(n1378) );
XOR2_X1 U1074 ( .A(G104), .B(KEYINPUT18), .Z(n1326) );
XNOR2_X1 U1075 ( .A(n1379), .B(n1380), .ZN(n1175) );
NOR2_X1 U1076 ( .A1(KEYINPUT48), .A2(G116), .ZN(n1380) );
XNOR2_X1 U1077 ( .A(G119), .B(G113), .ZN(n1379) );
XNOR2_X1 U1078 ( .A(n1178), .B(n1228), .ZN(n1365) );
XNOR2_X1 U1079 ( .A(G122), .B(n1221), .ZN(n1178) );
NAND2_X1 U1080 ( .A1(n1381), .A2(n1074), .ZN(n1292) );
INV_X1 U1081 ( .A(n1294), .ZN(n1074) );
XOR2_X1 U1082 ( .A(n1382), .B(n1200), .Z(n1294) );
INV_X1 U1083 ( .A(G472), .ZN(n1200) );
NAND2_X1 U1084 ( .A1(n1383), .A2(n1112), .ZN(n1382) );
XNOR2_X1 U1085 ( .A(n1193), .B(n1384), .ZN(n1383) );
XOR2_X1 U1086 ( .A(n1385), .B(KEYINPUT9), .Z(n1384) );
NAND2_X1 U1087 ( .A1(n1197), .A2(n1206), .ZN(n1385) );
NAND2_X1 U1088 ( .A1(n1386), .A2(n1387), .ZN(n1206) );
XNOR2_X1 U1089 ( .A(n1225), .B(n1228), .ZN(n1386) );
NAND2_X1 U1090 ( .A1(n1388), .A2(n1389), .ZN(n1197) );
XNOR2_X1 U1091 ( .A(n1225), .B(n1152), .ZN(n1389) );
INV_X1 U1092 ( .A(n1228), .ZN(n1152) );
XOR2_X1 U1093 ( .A(G128), .B(n1335), .Z(n1228) );
XOR2_X1 U1094 ( .A(G143), .B(G146), .Z(n1335) );
XNOR2_X1 U1095 ( .A(n1390), .B(n1391), .ZN(n1225) );
XOR2_X1 U1096 ( .A(KEYINPUT55), .B(G137), .Z(n1391) );
XNOR2_X1 U1097 ( .A(G131), .B(G134), .ZN(n1390) );
INV_X1 U1098 ( .A(n1387), .ZN(n1388) );
NAND2_X1 U1099 ( .A1(n1392), .A2(n1393), .ZN(n1387) );
NAND2_X1 U1100 ( .A1(G113), .A2(n1394), .ZN(n1393) );
XOR2_X1 U1101 ( .A(n1395), .B(KEYINPUT3), .Z(n1392) );
OR2_X1 U1102 ( .A1(n1394), .A2(G113), .ZN(n1395) );
XOR2_X1 U1103 ( .A(G116), .B(n1396), .Z(n1394) );
XNOR2_X1 U1104 ( .A(KEYINPUT54), .B(n1296), .ZN(n1396) );
INV_X1 U1105 ( .A(G119), .ZN(n1296) );
XNOR2_X1 U1106 ( .A(n1397), .B(G101), .ZN(n1193) );
NAND2_X1 U1107 ( .A1(G210), .A2(n1339), .ZN(n1397) );
NOR2_X1 U1108 ( .A1(G953), .A2(G237), .ZN(n1339) );
XNOR2_X1 U1109 ( .A(n1072), .B(KEYINPUT31), .ZN(n1381) );
XOR2_X1 U1110 ( .A(n1106), .B(n1398), .Z(n1072) );
NOR2_X1 U1111 ( .A1(n1399), .A2(KEYINPUT36), .ZN(n1398) );
INV_X1 U1112 ( .A(n1107), .ZN(n1399) );
NAND2_X1 U1113 ( .A1(G217), .A2(n1308), .ZN(n1107) );
NAND2_X1 U1114 ( .A1(G234), .A2(n1112), .ZN(n1308) );
AND2_X1 U1115 ( .A1(n1124), .A2(n1112), .ZN(n1106) );
INV_X1 U1116 ( .A(G902), .ZN(n1112) );
XNOR2_X1 U1117 ( .A(n1400), .B(n1401), .ZN(n1124) );
XNOR2_X1 U1118 ( .A(n1402), .B(n1336), .ZN(n1401) );
XNOR2_X1 U1119 ( .A(G125), .B(n1149), .ZN(n1336) );
INV_X1 U1120 ( .A(G140), .ZN(n1149) );
NAND2_X1 U1121 ( .A1(G221), .A2(n1359), .ZN(n1402) );
AND2_X1 U1122 ( .A1(G234), .A2(n1070), .ZN(n1359) );
INV_X1 U1123 ( .A(G953), .ZN(n1070) );
XOR2_X1 U1124 ( .A(n1403), .B(n1404), .Z(n1400) );
XOR2_X1 U1125 ( .A(G146), .B(G137), .Z(n1404) );
NAND2_X1 U1126 ( .A1(n1405), .A2(n1406), .ZN(n1403) );
OR2_X1 U1127 ( .A1(n1407), .A2(G110), .ZN(n1406) );
XOR2_X1 U1128 ( .A(n1408), .B(KEYINPUT5), .Z(n1405) );
NAND2_X1 U1129 ( .A1(G110), .A2(n1407), .ZN(n1408) );
XNOR2_X1 U1130 ( .A(G119), .B(n1280), .ZN(n1407) );
INV_X1 U1131 ( .A(G128), .ZN(n1280) );
INV_X1 U1132 ( .A(G110), .ZN(n1221) );
endmodule


