//Key = 1010111111110111000010000110111000101111001001011111100000110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389;

XOR2_X1 U751 ( .A(G107), .B(n1059), .Z(G9) );
NOR2_X1 U752 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U753 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1064), .A2(n1065), .A3(G953), .A4(n1066), .ZN(n1063) );
NOR4_X1 U755 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1065) );
NAND2_X1 U756 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NAND2_X1 U757 ( .A1(n1061), .A2(n1073), .ZN(n1072) );
NAND3_X1 U758 ( .A1(G214), .A2(n1074), .A3(n1075), .ZN(n1073) );
INV_X1 U759 ( .A(n1076), .ZN(n1067) );
NAND2_X1 U760 ( .A1(n1077), .A2(n1078), .ZN(n1064) );
NAND2_X1 U761 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U762 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U763 ( .A1(KEYINPUT3), .A2(n1083), .ZN(n1082) );
NAND4_X1 U764 ( .A1(n1084), .A2(n1085), .A3(n1071), .A4(n1086), .ZN(n1083) );
NAND2_X1 U765 ( .A1(n1084), .A2(n1087), .ZN(n1081) );
NAND2_X1 U766 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U767 ( .A1(n1071), .A2(n1090), .A3(n1085), .ZN(n1089) );
NAND2_X1 U768 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U769 ( .A1(n1086), .A2(n1093), .ZN(n1092) );
INV_X1 U770 ( .A(KEYINPUT3), .ZN(n1093) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1094), .ZN(n1088) );
NAND2_X1 U772 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1097), .ZN(n1096) );
NAND2_X1 U774 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND3_X1 U775 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
INV_X1 U776 ( .A(KEYINPUT22), .ZN(n1101) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1103), .ZN(n1095) );
NAND3_X1 U778 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NAND2_X1 U779 ( .A1(KEYINPUT22), .A2(n1071), .ZN(n1104) );
INV_X1 U780 ( .A(n1070), .ZN(n1084) );
NOR3_X1 U781 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1062) );
AND4_X1 U782 ( .A1(n1107), .A2(n1079), .A3(n1108), .A4(n1109), .ZN(n1066) );
NOR4_X1 U783 ( .A1(n1102), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1109) );
XOR2_X1 U784 ( .A(n1113), .B(G469), .Z(n1110) );
NAND2_X1 U785 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XNOR2_X1 U786 ( .A(KEYINPUT62), .B(KEYINPUT21), .ZN(n1114) );
XNOR2_X1 U787 ( .A(n1116), .B(G475), .ZN(n1108) );
XOR2_X1 U788 ( .A(n1117), .B(G472), .Z(n1107) );
XOR2_X1 U789 ( .A(n1118), .B(n1119), .Z(G72) );
XOR2_X1 U790 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U791 ( .A1(G953), .A2(n1122), .ZN(n1121) );
NOR2_X1 U792 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U793 ( .A(KEYINPUT17), .B(n1125), .Z(n1124) );
NAND2_X1 U794 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NAND2_X1 U795 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XOR2_X1 U796 ( .A(n1129), .B(n1130), .Z(n1126) );
XOR2_X1 U797 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U798 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U799 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1133) );
XNOR2_X1 U800 ( .A(n1135), .B(n1136), .ZN(n1129) );
XOR2_X1 U801 ( .A(KEYINPUT45), .B(G137), .Z(n1136) );
NAND2_X1 U802 ( .A1(G953), .A2(n1137), .ZN(n1118) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1137) );
XOR2_X1 U804 ( .A(n1138), .B(n1139), .Z(G69) );
NAND2_X1 U805 ( .A1(G953), .A2(n1140), .ZN(n1139) );
NAND2_X1 U806 ( .A1(G898), .A2(G224), .ZN(n1140) );
NAND4_X1 U807 ( .A1(KEYINPUT25), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1138) );
NAND3_X1 U808 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
NAND2_X1 U809 ( .A1(G953), .A2(n1147), .ZN(n1142) );
NAND2_X1 U810 ( .A1(G898), .A2(n1144), .ZN(n1147) );
OR2_X1 U811 ( .A1(n1145), .A2(n1144), .ZN(n1141) );
XOR2_X1 U812 ( .A(n1148), .B(n1149), .Z(n1144) );
NAND2_X1 U813 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NAND2_X1 U814 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U815 ( .A(KEYINPUT15), .B(n1154), .Z(n1150) );
NOR2_X1 U816 ( .A1(n1152), .A2(n1153), .ZN(n1154) );
NOR2_X1 U817 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U818 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U819 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NOR2_X1 U820 ( .A1(n1155), .A2(n1161), .ZN(G63) );
XOR2_X1 U821 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND3_X1 U822 ( .A1(n1159), .A2(G478), .A3(KEYINPUT2), .ZN(n1162) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1164), .ZN(G60) );
NOR3_X1 U824 ( .A1(n1116), .A2(n1165), .A3(n1166), .ZN(n1164) );
AND3_X1 U825 ( .A1(n1167), .A2(G475), .A3(n1159), .ZN(n1166) );
NOR2_X1 U826 ( .A1(n1168), .A2(n1167), .ZN(n1165) );
NOR2_X1 U827 ( .A1(n1077), .A2(n1169), .ZN(n1168) );
XNOR2_X1 U828 ( .A(G104), .B(n1170), .ZN(G6) );
NAND4_X1 U829 ( .A1(n1171), .A2(n1071), .A3(n1172), .A4(n1173), .ZN(n1170) );
XNOR2_X1 U830 ( .A(KEYINPUT56), .B(n1091), .ZN(n1172) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1174), .ZN(G57) );
XOR2_X1 U832 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U833 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U834 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U835 ( .A1(KEYINPUT60), .A2(n1181), .ZN(n1180) );
NAND2_X1 U836 ( .A1(n1159), .A2(G472), .ZN(n1179) );
XOR2_X1 U837 ( .A(n1182), .B(n1183), .Z(n1175) );
XNOR2_X1 U838 ( .A(n1184), .B(G101), .ZN(n1183) );
NAND2_X1 U839 ( .A1(KEYINPUT7), .A2(n1185), .ZN(n1182) );
NOR2_X1 U840 ( .A1(n1155), .A2(n1186), .ZN(G54) );
XOR2_X1 U841 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U842 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U843 ( .A(n1191), .B(n1192), .ZN(n1190) );
NAND2_X1 U844 ( .A1(n1159), .A2(G469), .ZN(n1191) );
XOR2_X1 U845 ( .A(n1193), .B(n1194), .Z(n1187) );
XNOR2_X1 U846 ( .A(n1195), .B(KEYINPUT47), .ZN(n1194) );
NAND2_X1 U847 ( .A1(n1196), .A2(KEYINPUT39), .ZN(n1195) );
XOR2_X1 U848 ( .A(n1197), .B(KEYINPUT23), .Z(n1196) );
NAND2_X1 U849 ( .A1(KEYINPUT34), .A2(n1198), .ZN(n1193) );
NOR2_X1 U850 ( .A1(n1155), .A2(n1199), .ZN(G51) );
XOR2_X1 U851 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U852 ( .A(n1202), .B(n1203), .ZN(n1201) );
NAND2_X1 U853 ( .A1(n1159), .A2(n1204), .ZN(n1202) );
NOR2_X1 U854 ( .A1(n1205), .A2(n1077), .ZN(n1159) );
NOR3_X1 U855 ( .A1(n1123), .A2(n1125), .A3(n1145), .ZN(n1077) );
NAND4_X1 U856 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1145) );
AND3_X1 U857 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NAND2_X1 U858 ( .A1(n1213), .A2(n1214), .ZN(n1208) );
NAND3_X1 U859 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
XOR2_X1 U860 ( .A(n1218), .B(KEYINPUT53), .Z(n1217) );
NAND4_X1 U861 ( .A1(n1219), .A2(n1071), .A3(n1220), .A4(n1173), .ZN(n1216) );
XNOR2_X1 U862 ( .A(KEYINPUT9), .B(n1060), .ZN(n1215) );
NAND4_X1 U863 ( .A1(n1071), .A2(n1220), .A3(n1086), .A4(n1173), .ZN(n1060) );
NAND3_X1 U864 ( .A1(n1076), .A2(n1221), .A3(n1222), .ZN(n1206) );
AND2_X1 U865 ( .A1(n1079), .A2(n1223), .ZN(n1125) );
XOR2_X1 U866 ( .A(KEYINPUT46), .B(n1224), .Z(n1223) );
NAND4_X1 U867 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1123) );
AND3_X1 U868 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
NAND2_X1 U869 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
NAND2_X1 U870 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND3_X1 U871 ( .A1(n1236), .A2(n1213), .A3(n1237), .ZN(n1235) );
NAND2_X1 U872 ( .A1(n1079), .A2(n1238), .ZN(n1234) );
XOR2_X1 U873 ( .A(KEYINPUT24), .B(n1086), .Z(n1238) );
XOR2_X1 U874 ( .A(n1239), .B(n1240), .Z(n1200) );
NOR2_X1 U875 ( .A1(KEYINPUT41), .A2(n1241), .ZN(n1240) );
NOR2_X1 U876 ( .A1(n1146), .A2(G952), .ZN(n1155) );
XOR2_X1 U877 ( .A(n1225), .B(n1242), .Z(G48) );
NAND2_X1 U878 ( .A1(KEYINPUT48), .A2(G146), .ZN(n1242) );
NAND3_X1 U879 ( .A1(n1243), .A2(n1213), .A3(n1221), .ZN(n1225) );
XNOR2_X1 U880 ( .A(G143), .B(n1244), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1236), .A2(n1213), .A3(n1237), .A4(n1245), .ZN(n1244) );
NOR3_X1 U882 ( .A1(n1246), .A2(n1105), .A3(n1098), .ZN(n1245) );
XNOR2_X1 U883 ( .A(KEYINPUT32), .B(n1247), .ZN(n1246) );
XNOR2_X1 U884 ( .A(G140), .B(n1226), .ZN(G42) );
NAND3_X1 U885 ( .A1(n1079), .A2(n1248), .A3(n1243), .ZN(n1226) );
XNOR2_X1 U886 ( .A(G137), .B(n1229), .ZN(G39) );
NAND3_X1 U887 ( .A1(n1076), .A2(n1221), .A3(n1249), .ZN(n1229) );
NOR3_X1 U888 ( .A1(n1098), .A2(n1250), .A3(n1251), .ZN(n1249) );
XOR2_X1 U889 ( .A(n1252), .B(G134), .Z(G36) );
NAND2_X1 U890 ( .A1(KEYINPUT26), .A2(n1253), .ZN(n1252) );
NAND3_X1 U891 ( .A1(n1079), .A2(n1086), .A3(n1232), .ZN(n1253) );
NOR3_X1 U892 ( .A1(n1098), .A2(n1250), .A3(n1105), .ZN(n1232) );
INV_X1 U893 ( .A(n1254), .ZN(n1105) );
NAND2_X1 U894 ( .A1(n1255), .A2(n1256), .ZN(G33) );
OR2_X1 U895 ( .A1(n1257), .A2(KEYINPUT29), .ZN(n1256) );
XOR2_X1 U896 ( .A(n1258), .B(n1259), .Z(n1255) );
NAND2_X1 U897 ( .A1(n1224), .A2(n1079), .ZN(n1259) );
INV_X1 U898 ( .A(n1251), .ZN(n1079) );
NAND2_X1 U899 ( .A1(n1075), .A2(n1260), .ZN(n1251) );
NAND2_X1 U900 ( .A1(G214), .A2(n1074), .ZN(n1260) );
AND2_X1 U901 ( .A1(n1254), .A2(n1243), .ZN(n1224) );
NOR3_X1 U902 ( .A1(n1098), .A2(n1250), .A3(n1091), .ZN(n1243) );
INV_X1 U903 ( .A(n1219), .ZN(n1091) );
XOR2_X1 U904 ( .A(n1220), .B(KEYINPUT30), .Z(n1098) );
NAND2_X1 U905 ( .A1(KEYINPUT29), .A2(n1257), .ZN(n1258) );
XOR2_X1 U906 ( .A(n1231), .B(n1261), .Z(G30) );
XNOR2_X1 U907 ( .A(KEYINPUT4), .B(n1262), .ZN(n1261) );
NAND4_X1 U908 ( .A1(n1171), .A2(n1221), .A3(n1086), .A4(n1247), .ZN(n1231) );
XNOR2_X1 U909 ( .A(n1263), .B(n1264), .ZN(G3) );
NOR2_X1 U910 ( .A1(n1061), .A2(n1218), .ZN(n1264) );
NAND4_X1 U911 ( .A1(n1076), .A2(n1254), .A3(n1220), .A4(n1173), .ZN(n1218) );
XNOR2_X1 U912 ( .A(G125), .B(n1230), .ZN(G27) );
NAND4_X1 U913 ( .A1(n1085), .A2(n1219), .A3(n1265), .A4(n1213), .ZN(n1230) );
NOR2_X1 U914 ( .A1(n1250), .A2(n1106), .ZN(n1265) );
INV_X1 U915 ( .A(n1248), .ZN(n1106) );
INV_X1 U916 ( .A(n1247), .ZN(n1250) );
NAND2_X1 U917 ( .A1(n1070), .A2(n1266), .ZN(n1247) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1267), .A4(n1128), .ZN(n1266) );
INV_X1 U919 ( .A(G900), .ZN(n1128) );
XNOR2_X1 U920 ( .A(G122), .B(n1207), .ZN(G24) );
NAND4_X1 U921 ( .A1(n1222), .A2(n1237), .A3(n1236), .A4(n1071), .ZN(n1207) );
NOR2_X1 U922 ( .A1(n1268), .A2(n1269), .ZN(n1071) );
NAND3_X1 U923 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(G21) );
NAND2_X1 U924 ( .A1(G119), .A2(n1273), .ZN(n1272) );
NAND3_X1 U925 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NAND2_X1 U926 ( .A1(KEYINPUT38), .A2(n1277), .ZN(n1276) );
NAND2_X1 U927 ( .A1(KEYINPUT63), .A2(n1278), .ZN(n1275) );
NAND2_X1 U928 ( .A1(n1279), .A2(n1280), .ZN(n1274) );
INV_X1 U929 ( .A(KEYINPUT63), .ZN(n1280) );
NAND2_X1 U930 ( .A1(n1278), .A2(n1281), .ZN(n1279) );
NAND2_X1 U931 ( .A1(KEYINPUT8), .A2(n1282), .ZN(n1281) );
NAND4_X1 U932 ( .A1(n1278), .A2(n1283), .A3(KEYINPUT38), .A4(KEYINPUT8), .ZN(n1271) );
NAND2_X1 U933 ( .A1(n1284), .A2(n1277), .ZN(n1270) );
INV_X1 U934 ( .A(KEYINPUT8), .ZN(n1277) );
NAND2_X1 U935 ( .A1(n1278), .A2(n1285), .ZN(n1284) );
NAND2_X1 U936 ( .A1(n1283), .A2(n1282), .ZN(n1285) );
INV_X1 U937 ( .A(KEYINPUT38), .ZN(n1282) );
AND4_X1 U938 ( .A1(n1076), .A2(n1221), .A3(n1286), .A4(n1287), .ZN(n1278) );
OR2_X1 U939 ( .A1(n1222), .A2(KEYINPUT16), .ZN(n1287) );
NAND2_X1 U940 ( .A1(KEYINPUT16), .A2(n1288), .ZN(n1286) );
NAND3_X1 U941 ( .A1(n1173), .A2(n1061), .A3(n1085), .ZN(n1288) );
INV_X1 U942 ( .A(n1213), .ZN(n1061) );
XNOR2_X1 U943 ( .A(G116), .B(n1210), .ZN(G18) );
NAND3_X1 U944 ( .A1(n1254), .A2(n1086), .A3(n1222), .ZN(n1210) );
AND2_X1 U945 ( .A1(n1236), .A2(n1289), .ZN(n1086) );
XNOR2_X1 U946 ( .A(n1111), .B(KEYINPUT0), .ZN(n1236) );
XNOR2_X1 U947 ( .A(n1212), .B(n1290), .ZN(G15) );
NOR2_X1 U948 ( .A1(KEYINPUT33), .A2(n1291), .ZN(n1290) );
NAND3_X1 U949 ( .A1(n1254), .A2(n1219), .A3(n1222), .ZN(n1212) );
AND3_X1 U950 ( .A1(n1213), .A2(n1173), .A3(n1085), .ZN(n1222) );
INV_X1 U951 ( .A(n1069), .ZN(n1085) );
NAND2_X1 U952 ( .A1(n1100), .A2(n1292), .ZN(n1069) );
NOR2_X1 U953 ( .A1(n1289), .A2(n1111), .ZN(n1219) );
NOR2_X1 U954 ( .A1(n1269), .A2(n1293), .ZN(n1254) );
XNOR2_X1 U955 ( .A(G110), .B(n1211), .ZN(G12) );
NAND4_X1 U956 ( .A1(n1076), .A2(n1171), .A3(n1248), .A4(n1173), .ZN(n1211) );
NAND2_X1 U957 ( .A1(n1294), .A2(n1070), .ZN(n1173) );
NAND3_X1 U958 ( .A1(n1267), .A2(n1146), .A3(G952), .ZN(n1070) );
NAND4_X1 U959 ( .A1(G953), .A2(G902), .A3(n1267), .A4(n1295), .ZN(n1294) );
INV_X1 U960 ( .A(G898), .ZN(n1295) );
NAND2_X1 U961 ( .A1(G234), .A2(G237), .ZN(n1267) );
NAND2_X1 U962 ( .A1(n1296), .A2(n1297), .ZN(n1248) );
NAND2_X1 U963 ( .A1(n1221), .A2(n1298), .ZN(n1297) );
INV_X1 U964 ( .A(KEYINPUT42), .ZN(n1298) );
AND2_X1 U965 ( .A1(n1269), .A2(n1268), .ZN(n1221) );
NAND3_X1 U966 ( .A1(n1293), .A2(n1269), .A3(KEYINPUT42), .ZN(n1296) );
XNOR2_X1 U967 ( .A(n1112), .B(KEYINPUT5), .ZN(n1269) );
XNOR2_X1 U968 ( .A(n1299), .B(n1160), .ZN(n1112) );
AND2_X1 U969 ( .A1(G217), .A2(n1300), .ZN(n1160) );
NAND2_X1 U970 ( .A1(n1158), .A2(n1205), .ZN(n1299) );
XOR2_X1 U971 ( .A(n1301), .B(n1302), .Z(n1158) );
XOR2_X1 U972 ( .A(G137), .B(n1303), .Z(n1302) );
AND3_X1 U973 ( .A1(G221), .A2(n1146), .A3(G234), .ZN(n1303) );
NAND2_X1 U974 ( .A1(n1304), .A2(n1305), .ZN(n1301) );
NAND2_X1 U975 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U976 ( .A(KEYINPUT14), .B(n1308), .Z(n1304) );
NOR2_X1 U977 ( .A1(n1306), .A2(n1307), .ZN(n1308) );
XNOR2_X1 U978 ( .A(n1309), .B(n1310), .ZN(n1307) );
XNOR2_X1 U979 ( .A(KEYINPUT59), .B(n1262), .ZN(n1310) );
INV_X1 U980 ( .A(G128), .ZN(n1262) );
XNOR2_X1 U981 ( .A(G110), .B(G119), .ZN(n1309) );
XOR2_X1 U982 ( .A(n1311), .B(n1312), .Z(n1306) );
XNOR2_X1 U983 ( .A(n1313), .B(KEYINPUT31), .ZN(n1312) );
NAND2_X1 U984 ( .A1(KEYINPUT28), .A2(n1314), .ZN(n1313) );
INV_X1 U985 ( .A(G140), .ZN(n1314) );
INV_X1 U986 ( .A(n1268), .ZN(n1293) );
NAND2_X1 U987 ( .A1(n1315), .A2(n1316), .ZN(n1268) );
NAND2_X1 U988 ( .A1(G472), .A2(n1117), .ZN(n1316) );
XOR2_X1 U989 ( .A(KEYINPUT61), .B(n1317), .Z(n1315) );
NOR2_X1 U990 ( .A1(G472), .A2(n1117), .ZN(n1317) );
NAND2_X1 U991 ( .A1(n1318), .A2(n1205), .ZN(n1117) );
XOR2_X1 U992 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U993 ( .A(n1321), .B(n1185), .ZN(n1320) );
INV_X1 U994 ( .A(n1322), .ZN(n1185) );
XNOR2_X1 U995 ( .A(n1181), .B(n1177), .ZN(n1321) );
XOR2_X1 U996 ( .A(n1323), .B(n1291), .Z(n1181) );
NAND2_X1 U997 ( .A1(KEYINPUT20), .A2(n1324), .ZN(n1323) );
XOR2_X1 U998 ( .A(n1325), .B(n1326), .Z(n1319) );
XNOR2_X1 U999 ( .A(KEYINPUT6), .B(n1263), .ZN(n1326) );
INV_X1 U1000 ( .A(G101), .ZN(n1263) );
NAND2_X1 U1001 ( .A1(KEYINPUT13), .A2(n1184), .ZN(n1325) );
AND3_X1 U1002 ( .A1(n1327), .A2(n1146), .A3(G210), .ZN(n1184) );
AND2_X1 U1003 ( .A1(n1213), .A2(n1220), .ZN(n1171) );
NOR2_X1 U1004 ( .A1(n1100), .A2(n1102), .ZN(n1220) );
INV_X1 U1005 ( .A(n1292), .ZN(n1102) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1300), .ZN(n1292) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1328), .ZN(n1300) );
XNOR2_X1 U1008 ( .A(n1115), .B(n1329), .ZN(n1100) );
XOR2_X1 U1009 ( .A(KEYINPUT11), .B(G469), .Z(n1329) );
NAND2_X1 U1010 ( .A1(n1330), .A2(n1205), .ZN(n1115) );
XOR2_X1 U1011 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1012 ( .A(n1189), .B(n1197), .ZN(n1332) );
XOR2_X1 U1013 ( .A(n1177), .B(n1131), .Z(n1189) );
XNOR2_X1 U1014 ( .A(n1333), .B(n1334), .ZN(n1131) );
NOR2_X1 U1015 ( .A1(G143), .A2(KEYINPUT40), .ZN(n1334) );
XNOR2_X1 U1016 ( .A(n1335), .B(n1336), .ZN(n1177) );
XOR2_X1 U1017 ( .A(G137), .B(G134), .Z(n1336) );
NAND2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1257), .ZN(n1335) );
XOR2_X1 U1019 ( .A(n1198), .B(n1192), .Z(n1331) );
XOR2_X1 U1020 ( .A(G110), .B(G140), .Z(n1192) );
AND2_X1 U1021 ( .A1(G227), .A2(n1146), .ZN(n1198) );
NOR2_X1 U1022 ( .A1(n1075), .A2(n1337), .ZN(n1213) );
AND2_X1 U1023 ( .A1(G214), .A2(n1074), .ZN(n1337) );
XOR2_X1 U1024 ( .A(n1338), .B(n1204), .Z(n1075) );
AND2_X1 U1025 ( .A1(G210), .A2(n1074), .ZN(n1204) );
NAND2_X1 U1026 ( .A1(n1339), .A2(n1328), .ZN(n1074) );
XNOR2_X1 U1027 ( .A(G902), .B(KEYINPUT19), .ZN(n1328) );
XNOR2_X1 U1028 ( .A(G237), .B(KEYINPUT18), .ZN(n1339) );
NAND3_X1 U1029 ( .A1(n1340), .A2(n1205), .A3(n1341), .ZN(n1338) );
XOR2_X1 U1030 ( .A(n1342), .B(KEYINPUT1), .Z(n1341) );
OR2_X1 U1031 ( .A1(n1203), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1032 ( .A1(n1343), .A2(n1203), .ZN(n1340) );
XNOR2_X1 U1033 ( .A(n1344), .B(n1152), .ZN(n1203) );
XNOR2_X1 U1034 ( .A(n1197), .B(KEYINPUT43), .ZN(n1152) );
XNOR2_X1 U1035 ( .A(G101), .B(n1345), .ZN(n1197) );
XOR2_X1 U1036 ( .A(G107), .B(G104), .Z(n1345) );
XNOR2_X1 U1037 ( .A(n1153), .B(n1149), .ZN(n1344) );
XNOR2_X1 U1038 ( .A(n1346), .B(G122), .ZN(n1149) );
INV_X1 U1039 ( .A(G110), .ZN(n1346) );
XOR2_X1 U1040 ( .A(n1347), .B(n1324), .Z(n1153) );
XOR2_X1 U1041 ( .A(n1283), .B(n1348), .Z(n1324) );
INV_X1 U1042 ( .A(G119), .ZN(n1283) );
NAND2_X1 U1043 ( .A1(KEYINPUT49), .A2(G113), .ZN(n1347) );
XOR2_X1 U1044 ( .A(n1241), .B(n1349), .Z(n1343) );
XNOR2_X1 U1045 ( .A(KEYINPUT50), .B(n1239), .ZN(n1349) );
NAND2_X1 U1046 ( .A1(G224), .A2(n1146), .ZN(n1239) );
XNOR2_X1 U1047 ( .A(n1322), .B(n1135), .ZN(n1241) );
INV_X1 U1048 ( .A(G125), .ZN(n1135) );
XOR2_X1 U1049 ( .A(n1350), .B(n1333), .Z(n1322) );
XNOR2_X1 U1050 ( .A(G146), .B(G128), .ZN(n1333) );
NAND2_X1 U1051 ( .A1(KEYINPUT51), .A2(n1351), .ZN(n1350) );
NOR2_X1 U1052 ( .A1(n1111), .A2(n1237), .ZN(n1076) );
INV_X1 U1053 ( .A(n1289), .ZN(n1237) );
NAND3_X1 U1054 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1289) );
NAND2_X1 U1055 ( .A1(KEYINPUT57), .A2(n1116), .ZN(n1354) );
NAND3_X1 U1056 ( .A1(n1355), .A2(n1356), .A3(n1169), .ZN(n1353) );
INV_X1 U1057 ( .A(KEYINPUT57), .ZN(n1356) );
OR2_X1 U1058 ( .A1(n1169), .A2(n1355), .ZN(n1352) );
NOR2_X1 U1059 ( .A1(n1116), .A2(KEYINPUT54), .ZN(n1355) );
NOR2_X1 U1060 ( .A1(n1167), .A2(G902), .ZN(n1116) );
XOR2_X1 U1061 ( .A(n1357), .B(n1358), .Z(n1167) );
XOR2_X1 U1062 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1063 ( .A(n1291), .B(G104), .ZN(n1360) );
INV_X1 U1064 ( .A(G113), .ZN(n1291) );
XNOR2_X1 U1065 ( .A(n1351), .B(G122), .ZN(n1359) );
XOR2_X1 U1066 ( .A(n1311), .B(n1361), .Z(n1357) );
XOR2_X1 U1067 ( .A(n1362), .B(n1134), .Z(n1361) );
XNOR2_X1 U1068 ( .A(n1257), .B(G140), .ZN(n1134) );
INV_X1 U1069 ( .A(G131), .ZN(n1257) );
AND3_X1 U1070 ( .A1(G214), .A2(n1146), .A3(n1327), .ZN(n1362) );
INV_X1 U1071 ( .A(G237), .ZN(n1327) );
XNOR2_X1 U1072 ( .A(G146), .B(G125), .ZN(n1311) );
INV_X1 U1073 ( .A(G475), .ZN(n1169) );
XNOR2_X1 U1074 ( .A(n1363), .B(G478), .ZN(n1111) );
NAND2_X1 U1075 ( .A1(n1163), .A2(n1205), .ZN(n1363) );
INV_X1 U1076 ( .A(G902), .ZN(n1205) );
XNOR2_X1 U1077 ( .A(n1364), .B(n1365), .ZN(n1163) );
AND3_X1 U1078 ( .A1(G217), .A2(n1146), .A3(G234), .ZN(n1365) );
INV_X1 U1079 ( .A(G953), .ZN(n1146) );
NAND2_X1 U1080 ( .A1(KEYINPUT36), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1081 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND3_X1 U1082 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1368) );
XOR2_X1 U1083 ( .A(n1372), .B(KEYINPUT35), .Z(n1367) );
NAND2_X1 U1084 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1085 ( .A1(n1371), .A2(n1369), .ZN(n1374) );
NAND2_X1 U1086 ( .A1(n1375), .A2(n1376), .ZN(n1369) );
XNOR2_X1 U1087 ( .A(n1377), .B(KEYINPUT55), .ZN(n1376) );
XNOR2_X1 U1088 ( .A(G128), .B(G143), .ZN(n1375) );
XNOR2_X1 U1089 ( .A(n1378), .B(KEYINPUT37), .ZN(n1371) );
NAND2_X1 U1090 ( .A1(n1379), .A2(n1377), .ZN(n1378) );
XOR2_X1 U1091 ( .A(G134), .B(KEYINPUT27), .Z(n1377) );
XNOR2_X1 U1092 ( .A(n1351), .B(G128), .ZN(n1379) );
INV_X1 U1093 ( .A(G143), .ZN(n1351) );
INV_X1 U1094 ( .A(n1370), .ZN(n1373) );
NAND3_X1 U1095 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1370) );
OR2_X1 U1096 ( .A1(n1383), .A2(G107), .ZN(n1382) );
NAND2_X1 U1097 ( .A1(n1384), .A2(n1385), .ZN(n1381) );
INV_X1 U1098 ( .A(KEYINPUT52), .ZN(n1385) );
NAND2_X1 U1099 ( .A1(n1386), .A2(G107), .ZN(n1384) );
XNOR2_X1 U1100 ( .A(n1383), .B(KEYINPUT10), .ZN(n1386) );
NAND2_X1 U1101 ( .A1(KEYINPUT52), .A2(n1387), .ZN(n1380) );
NAND2_X1 U1102 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
OR2_X1 U1103 ( .A1(n1383), .A2(KEYINPUT10), .ZN(n1389) );
NAND3_X1 U1104 ( .A1(G107), .A2(n1383), .A3(KEYINPUT10), .ZN(n1388) );
XOR2_X1 U1105 ( .A(G122), .B(n1348), .Z(n1383) );
XOR2_X1 U1106 ( .A(G116), .B(KEYINPUT12), .Z(n1348) );
endmodule


