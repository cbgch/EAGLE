//Key = 0010000011100101000000111100111110111111011100010001001101001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368;

XOR2_X1 U750 ( .A(G107), .B(n1043), .Z(G9) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U752 ( .A1(KEYINPUT49), .A2(n1046), .ZN(n1045) );
NOR2_X1 U753 ( .A1(KEYINPUT37), .A2(n1047), .ZN(n1044) );
NAND4_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(G75) );
NAND3_X1 U755 ( .A1(KEYINPUT21), .A2(n1052), .A3(n1053), .ZN(n1051) );
INV_X1 U756 ( .A(G952), .ZN(n1053) );
NAND2_X1 U757 ( .A1(G952), .A2(n1054), .ZN(n1050) );
NAND4_X1 U758 ( .A1(n1055), .A2(n1056), .A3(n1052), .A4(n1057), .ZN(n1054) );
NAND2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U761 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
INV_X1 U766 ( .A(n1073), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1065) );
NAND2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U769 ( .A1(n1067), .A2(n1078), .A3(n1074), .ZN(n1060) );
NAND3_X1 U770 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND2_X1 U771 ( .A1(n1062), .A2(n1082), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND3_X1 U774 ( .A1(n1087), .A2(n1064), .A3(n1088), .ZN(n1079) );
INV_X1 U775 ( .A(n1089), .ZN(n1058) );
INV_X1 U776 ( .A(n1090), .ZN(n1049) );
OR2_X1 U777 ( .A1(n1052), .A2(KEYINPUT21), .ZN(n1048) );
NAND4_X1 U778 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1052) );
NOR4_X1 U779 ( .A1(n1088), .A2(n1085), .A3(n1095), .A4(n1096), .ZN(n1094) );
XOR2_X1 U780 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U781 ( .A1(KEYINPUT26), .A2(n1099), .ZN(n1098) );
NOR2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U784 ( .A1(KEYINPUT9), .A2(n1104), .ZN(n1103) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(n1092) );
XOR2_X1 U786 ( .A(n1107), .B(G472), .Z(n1091) );
XOR2_X1 U787 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
XOR2_X1 U790 ( .A(KEYINPUT51), .B(G227), .Z(n1113) );
NOR2_X1 U791 ( .A1(KEYINPUT12), .A2(n1114), .ZN(n1108) );
XOR2_X1 U792 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U793 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U794 ( .A(n1119), .B(n1120), .ZN(n1118) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(n1119) );
NOR2_X1 U796 ( .A1(G900), .A2(n1057), .ZN(n1117) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1057), .ZN(n1115) );
NAND3_X1 U798 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
XNOR2_X1 U799 ( .A(KEYINPUT38), .B(n1127), .ZN(n1125) );
XOR2_X1 U800 ( .A(n1128), .B(n1129), .Z(G69) );
XOR2_X1 U801 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U802 ( .A1(n1132), .A2(n1111), .ZN(n1131) );
XNOR2_X1 U803 ( .A(G953), .B(KEYINPUT50), .ZN(n1111) );
NOR2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U805 ( .A(KEYINPUT60), .B(G224), .Z(n1134) );
NAND2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
XOR2_X1 U807 ( .A(KEYINPUT36), .B(n1137), .Z(n1136) );
NOR2_X1 U808 ( .A1(G898), .A2(n1057), .ZN(n1137) );
XOR2_X1 U809 ( .A(n1138), .B(n1139), .Z(n1135) );
NAND2_X1 U810 ( .A1(n1057), .A2(n1140), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1090), .A2(n1141), .ZN(G66) );
XOR2_X1 U812 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U813 ( .A1(n1144), .A2(n1106), .ZN(n1142) );
NOR2_X1 U814 ( .A1(n1090), .A2(n1145), .ZN(G63) );
XOR2_X1 U815 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1148), .ZN(n1146) );
XOR2_X1 U817 ( .A(KEYINPUT6), .B(G478), .Z(n1148) );
NOR2_X1 U818 ( .A1(n1090), .A2(n1149), .ZN(G60) );
XOR2_X1 U819 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U820 ( .A1(n1152), .A2(n1144), .ZN(n1150) );
XNOR2_X1 U821 ( .A(G475), .B(KEYINPUT22), .ZN(n1152) );
XNOR2_X1 U822 ( .A(G104), .B(n1153), .ZN(G6) );
NAND4_X1 U823 ( .A1(n1154), .A2(n1155), .A3(n1074), .A4(n1156), .ZN(n1153) );
XNOR2_X1 U824 ( .A(n1157), .B(KEYINPUT54), .ZN(n1154) );
NOR2_X1 U825 ( .A1(n1090), .A2(n1158), .ZN(G57) );
XOR2_X1 U826 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U827 ( .A(n1161), .B(n1162), .Z(n1159) );
NOR2_X1 U828 ( .A1(KEYINPUT33), .A2(n1163), .ZN(n1162) );
NAND2_X1 U829 ( .A1(n1144), .A2(G472), .ZN(n1161) );
NOR2_X1 U830 ( .A1(n1090), .A2(n1164), .ZN(G54) );
XOR2_X1 U831 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U832 ( .A1(n1144), .A2(G469), .ZN(n1166) );
NAND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1165) );
NAND2_X1 U834 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U835 ( .A(KEYINPUT35), .B(n1171), .Z(n1167) );
NOR2_X1 U836 ( .A1(n1172), .A2(n1170), .ZN(n1171) );
NAND2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U839 ( .A(KEYINPUT39), .B(n1177), .Z(n1175) );
XOR2_X1 U840 ( .A(KEYINPUT15), .B(n1178), .Z(n1173) );
XNOR2_X1 U841 ( .A(KEYINPUT13), .B(n1169), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1179), .A2(n1180), .ZN(n1169) );
OR2_X1 U843 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U844 ( .A1(n1183), .A2(n1182), .ZN(n1179) );
XOR2_X1 U845 ( .A(KEYINPUT53), .B(n1181), .Z(n1183) );
XNOR2_X1 U846 ( .A(n1120), .B(n1184), .ZN(n1181) );
XNOR2_X1 U847 ( .A(KEYINPUT7), .B(n1185), .ZN(n1184) );
NOR2_X1 U848 ( .A1(n1090), .A2(n1186), .ZN(G51) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U850 ( .A1(KEYINPUT55), .A2(n1189), .ZN(n1188) );
NAND2_X1 U851 ( .A1(n1144), .A2(n1104), .ZN(n1187) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1055), .ZN(n1144) );
AND3_X1 U853 ( .A1(n1191), .A2(n1126), .A3(n1192), .ZN(n1055) );
XOR2_X1 U854 ( .A(n1193), .B(KEYINPUT41), .Z(n1192) );
NAND2_X1 U855 ( .A1(n1124), .A2(n1127), .ZN(n1193) );
AND3_X1 U856 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1124) );
OR2_X1 U857 ( .A1(n1080), .A2(n1197), .ZN(n1196) );
NAND3_X1 U858 ( .A1(n1155), .A2(n1198), .A3(n1199), .ZN(n1194) );
AND3_X1 U859 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1126) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1203), .ZN(n1202) );
NAND2_X1 U861 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
OR2_X1 U862 ( .A1(n1197), .A2(n1206), .ZN(n1205) );
NAND2_X1 U863 ( .A1(n1199), .A2(n1207), .ZN(n1204) );
INV_X1 U864 ( .A(n1140), .ZN(n1191) );
NAND4_X1 U865 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1140) );
NOR3_X1 U866 ( .A1(n1212), .A2(n1213), .A3(n1046), .ZN(n1211) );
INV_X1 U867 ( .A(n1047), .ZN(n1046) );
NAND4_X1 U868 ( .A1(n1074), .A2(n1157), .A3(n1156), .A4(n1207), .ZN(n1047) );
INV_X1 U869 ( .A(n1214), .ZN(n1212) );
NAND2_X1 U870 ( .A1(n1215), .A2(n1198), .ZN(n1210) );
XOR2_X1 U871 ( .A(n1216), .B(KEYINPUT32), .Z(n1215) );
NAND2_X1 U872 ( .A1(n1156), .A2(n1217), .ZN(n1208) );
NAND2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U874 ( .A1(n1157), .A2(n1220), .ZN(n1218) );
NAND2_X1 U875 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U876 ( .A1(n1223), .A2(n1067), .ZN(n1222) );
XNOR2_X1 U877 ( .A(KEYINPUT31), .B(n1073), .ZN(n1223) );
NAND2_X1 U878 ( .A1(n1155), .A2(n1074), .ZN(n1221) );
NOR2_X1 U879 ( .A1(n1057), .A2(G952), .ZN(n1090) );
XNOR2_X1 U880 ( .A(G146), .B(n1224), .ZN(G48) );
NAND2_X1 U881 ( .A1(n1198), .A2(n1225), .ZN(n1224) );
XOR2_X1 U882 ( .A(KEYINPUT46), .B(n1226), .Z(n1225) );
NOR2_X1 U883 ( .A1(n1076), .A2(n1227), .ZN(n1226) );
INV_X1 U884 ( .A(n1155), .ZN(n1076) );
NAND2_X1 U885 ( .A1(n1228), .A2(n1229), .ZN(G45) );
NAND2_X1 U886 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U887 ( .A1(G143), .A2(n1232), .ZN(n1228) );
NAND2_X1 U888 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
OR2_X1 U889 ( .A1(n1127), .A2(KEYINPUT30), .ZN(n1234) );
NAND2_X1 U890 ( .A1(KEYINPUT30), .A2(n1235), .ZN(n1233) );
INV_X1 U891 ( .A(n1230), .ZN(n1235) );
NOR2_X1 U892 ( .A1(KEYINPUT58), .A2(n1127), .ZN(n1230) );
NAND4_X1 U893 ( .A1(n1095), .A2(n1236), .A3(n1198), .A4(n1100), .ZN(n1127) );
XNOR2_X1 U894 ( .A(n1237), .B(n1238), .ZN(G42) );
NOR3_X1 U895 ( .A1(n1080), .A2(KEYINPUT56), .A3(n1197), .ZN(n1238) );
NAND2_X1 U896 ( .A1(n1064), .A2(n1157), .ZN(n1080) );
XNOR2_X1 U897 ( .A(G137), .B(n1195), .ZN(G39) );
NAND3_X1 U898 ( .A1(n1064), .A2(n1067), .A3(n1199), .ZN(n1195) );
INV_X1 U899 ( .A(n1227), .ZN(n1199) );
XNOR2_X1 U900 ( .A(G134), .B(n1200), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1064), .A2(n1207), .A3(n1236), .ZN(n1200) );
XNOR2_X1 U902 ( .A(G131), .B(n1201), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1064), .A2(n1155), .A3(n1236), .ZN(n1201) );
AND4_X1 U904 ( .A1(n1071), .A2(n1157), .A3(n1072), .A4(n1239), .ZN(n1236) );
AND2_X1 U905 ( .A1(n1086), .A2(n1240), .ZN(n1064) );
XOR2_X1 U906 ( .A(G128), .B(n1241), .Z(G30) );
NOR4_X1 U907 ( .A1(KEYINPUT17), .A2(n1083), .A3(n1077), .A4(n1227), .ZN(n1241) );
NAND4_X1 U908 ( .A1(n1242), .A2(n1071), .A3(n1157), .A4(n1239), .ZN(n1227) );
INV_X1 U909 ( .A(n1207), .ZN(n1077) );
XNOR2_X1 U910 ( .A(n1243), .B(n1244), .ZN(G3) );
NOR2_X1 U911 ( .A1(n1083), .A2(n1216), .ZN(n1244) );
NAND4_X1 U912 ( .A1(n1071), .A2(n1157), .A3(n1245), .A4(n1067), .ZN(n1216) );
NOR2_X1 U913 ( .A1(n1246), .A2(n1242), .ZN(n1245) );
XOR2_X1 U914 ( .A(G125), .B(n1247), .Z(G27) );
NOR3_X1 U915 ( .A1(n1248), .A2(n1206), .A3(n1197), .ZN(n1247) );
NAND3_X1 U916 ( .A1(n1073), .A2(n1239), .A3(n1155), .ZN(n1197) );
NAND2_X1 U917 ( .A1(n1089), .A2(n1249), .ZN(n1239) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1112), .ZN(n1249) );
INV_X1 U919 ( .A(G900), .ZN(n1112) );
XNOR2_X1 U920 ( .A(KEYINPUT63), .B(n1083), .ZN(n1248) );
XNOR2_X1 U921 ( .A(n1251), .B(n1252), .ZN(G24) );
NOR3_X1 U922 ( .A1(n1219), .A2(n1253), .A3(n1254), .ZN(n1252) );
NOR2_X1 U923 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U924 ( .A(KEYINPUT48), .ZN(n1256) );
NOR2_X1 U925 ( .A1(n1083), .A2(n1257), .ZN(n1255) );
NOR2_X1 U926 ( .A1(KEYINPUT48), .A2(n1156), .ZN(n1253) );
NAND4_X1 U927 ( .A1(n1095), .A2(n1062), .A3(n1074), .A4(n1100), .ZN(n1219) );
XNOR2_X1 U928 ( .A(G119), .B(n1209), .ZN(G21) );
NAND3_X1 U929 ( .A1(n1258), .A2(n1067), .A3(n1242), .ZN(n1209) );
XOR2_X1 U930 ( .A(n1259), .B(G116), .Z(G18) );
NAND2_X1 U931 ( .A1(KEYINPUT29), .A2(n1214), .ZN(n1259) );
NAND3_X1 U932 ( .A1(n1207), .A2(n1072), .A3(n1258), .ZN(n1214) );
NOR2_X1 U933 ( .A1(n1260), .A2(n1095), .ZN(n1207) );
INV_X1 U934 ( .A(n1100), .ZN(n1260) );
XOR2_X1 U935 ( .A(G113), .B(n1213), .Z(G15) );
AND3_X1 U936 ( .A1(n1258), .A2(n1072), .A3(n1155), .ZN(n1213) );
AND3_X1 U937 ( .A1(n1071), .A2(n1156), .A3(n1062), .ZN(n1258) );
INV_X1 U938 ( .A(n1206), .ZN(n1062) );
NAND2_X1 U939 ( .A1(n1087), .A2(n1261), .ZN(n1206) );
NOR2_X1 U940 ( .A1(n1083), .A2(n1246), .ZN(n1156) );
INV_X1 U941 ( .A(n1257), .ZN(n1246) );
INV_X1 U942 ( .A(n1198), .ZN(n1083) );
XNOR2_X1 U943 ( .A(G110), .B(n1262), .ZN(G12) );
NAND4_X1 U944 ( .A1(n1067), .A2(n1073), .A3(n1263), .A4(n1264), .ZN(n1262) );
AND2_X1 U945 ( .A1(n1198), .A2(n1157), .ZN(n1264) );
NOR2_X1 U946 ( .A1(n1087), .A2(n1088), .ZN(n1157) );
INV_X1 U947 ( .A(n1261), .ZN(n1088) );
NAND2_X1 U948 ( .A1(n1265), .A2(G221), .ZN(n1261) );
XOR2_X1 U949 ( .A(n1266), .B(KEYINPUT4), .Z(n1265) );
XOR2_X1 U950 ( .A(n1097), .B(n1099), .Z(n1087) );
XOR2_X1 U951 ( .A(G469), .B(KEYINPUT11), .Z(n1099) );
NAND2_X1 U952 ( .A1(n1267), .A2(n1268), .ZN(n1097) );
XOR2_X1 U953 ( .A(n1269), .B(n1270), .Z(n1267) );
XNOR2_X1 U954 ( .A(n1182), .B(n1120), .ZN(n1270) );
XNOR2_X1 U955 ( .A(n1271), .B(n1272), .ZN(n1120) );
NOR2_X1 U956 ( .A1(G143), .A2(KEYINPUT45), .ZN(n1272) );
XOR2_X1 U957 ( .A(n1273), .B(n1243), .Z(n1182) );
NAND3_X1 U958 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NAND2_X1 U959 ( .A1(G104), .A2(n1277), .ZN(n1276) );
NAND2_X1 U960 ( .A1(n1278), .A2(n1279), .ZN(n1275) );
INV_X1 U961 ( .A(KEYINPUT42), .ZN(n1279) );
NAND2_X1 U962 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
XNOR2_X1 U963 ( .A(KEYINPUT27), .B(n1277), .ZN(n1280) );
NAND2_X1 U964 ( .A1(KEYINPUT42), .A2(n1282), .ZN(n1274) );
NAND2_X1 U965 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
OR3_X1 U966 ( .A1(n1277), .A2(G104), .A3(KEYINPUT27), .ZN(n1284) );
NAND2_X1 U967 ( .A1(KEYINPUT27), .A2(n1277), .ZN(n1283) );
NOR2_X1 U968 ( .A1(n1285), .A2(n1286), .ZN(n1269) );
NOR2_X1 U969 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U970 ( .A(n1177), .B(n1289), .ZN(n1288) );
NOR2_X1 U971 ( .A1(n1290), .A2(n1185), .ZN(n1285) );
NOR2_X1 U972 ( .A1(n1291), .A2(n1178), .ZN(n1290) );
AND2_X1 U973 ( .A1(n1177), .A2(n1289), .ZN(n1178) );
NOR2_X1 U974 ( .A1(n1177), .A2(n1289), .ZN(n1291) );
INV_X1 U975 ( .A(n1176), .ZN(n1289) );
XOR2_X1 U976 ( .A(G140), .B(G110), .Z(n1176) );
AND2_X1 U977 ( .A1(G227), .A2(n1057), .ZN(n1177) );
NOR2_X1 U978 ( .A1(n1086), .A2(n1085), .ZN(n1198) );
INV_X1 U979 ( .A(n1240), .ZN(n1085) );
NAND2_X1 U980 ( .A1(G214), .A2(n1292), .ZN(n1240) );
XNOR2_X1 U981 ( .A(n1102), .B(n1293), .ZN(n1086) );
XOR2_X1 U982 ( .A(KEYINPUT2), .B(n1104), .Z(n1293) );
AND2_X1 U983 ( .A1(G210), .A2(n1292), .ZN(n1104) );
NAND2_X1 U984 ( .A1(n1294), .A2(n1190), .ZN(n1292) );
INV_X1 U985 ( .A(G237), .ZN(n1294) );
NAND2_X1 U986 ( .A1(n1295), .A2(n1268), .ZN(n1102) );
XOR2_X1 U987 ( .A(KEYINPUT10), .B(n1189), .Z(n1295) );
XNOR2_X1 U988 ( .A(n1296), .B(n1297), .ZN(n1189) );
XOR2_X1 U989 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U990 ( .A(G125), .B(n1300), .Z(n1299) );
NOR2_X1 U991 ( .A1(KEYINPUT0), .A2(n1139), .ZN(n1300) );
XNOR2_X1 U992 ( .A(n1301), .B(n1302), .ZN(n1139) );
AND2_X1 U993 ( .A1(n1057), .A2(G224), .ZN(n1298) );
XOR2_X1 U994 ( .A(n1138), .B(n1303), .Z(n1296) );
XOR2_X1 U995 ( .A(n1304), .B(n1305), .Z(n1138) );
XNOR2_X1 U996 ( .A(n1277), .B(n1306), .ZN(n1305) );
NAND2_X1 U997 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U998 ( .A1(n1309), .A2(n1251), .ZN(n1308) );
XNOR2_X1 U999 ( .A(G110), .B(KEYINPUT40), .ZN(n1309) );
NAND2_X1 U1000 ( .A1(n1310), .A2(G122), .ZN(n1307) );
XOR2_X1 U1001 ( .A(KEYINPUT62), .B(G110), .Z(n1310) );
XNOR2_X1 U1002 ( .A(G101), .B(n1311), .ZN(n1304) );
NOR2_X1 U1003 ( .A1(G104), .A2(KEYINPUT14), .ZN(n1311) );
XNOR2_X1 U1004 ( .A(KEYINPUT47), .B(n1257), .ZN(n1263) );
NAND2_X1 U1005 ( .A1(n1089), .A2(n1312), .ZN(n1257) );
NAND4_X1 U1006 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1133), .ZN(n1312) );
INV_X1 U1007 ( .A(G898), .ZN(n1133) );
NAND3_X1 U1008 ( .A1(n1250), .A2(n1057), .A3(G952), .ZN(n1089) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1250) );
NAND2_X1 U1010 ( .A1(n1313), .A2(n1314), .ZN(n1073) );
OR3_X1 U1011 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT59), .ZN(n1314) );
NAND2_X1 U1012 ( .A1(KEYINPUT59), .A2(n1074), .ZN(n1313) );
NOR2_X1 U1013 ( .A1(n1242), .A2(n1071), .ZN(n1074) );
XOR2_X1 U1014 ( .A(n1315), .B(G472), .Z(n1071) );
NAND2_X1 U1015 ( .A1(KEYINPUT57), .A2(n1107), .ZN(n1315) );
NAND2_X1 U1016 ( .A1(n1268), .A2(n1316), .ZN(n1107) );
XNOR2_X1 U1017 ( .A(n1160), .B(n1163), .ZN(n1316) );
AND2_X1 U1018 ( .A1(n1317), .A2(n1318), .ZN(n1163) );
NAND2_X1 U1019 ( .A1(n1319), .A2(n1243), .ZN(n1318) );
INV_X1 U1020 ( .A(G101), .ZN(n1243) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1320), .ZN(n1319) );
NAND3_X1 U1022 ( .A1(G210), .A2(n1320), .A3(G101), .ZN(n1317) );
XNOR2_X1 U1023 ( .A(n1321), .B(n1322), .ZN(n1160) );
XNOR2_X1 U1024 ( .A(n1303), .B(n1185), .ZN(n1322) );
INV_X1 U1025 ( .A(n1287), .ZN(n1185) );
XOR2_X1 U1026 ( .A(G131), .B(n1323), .Z(n1287) );
NOR2_X1 U1027 ( .A1(KEYINPUT3), .A2(n1122), .ZN(n1323) );
XNOR2_X1 U1028 ( .A(G134), .B(G137), .ZN(n1122) );
XNOR2_X1 U1029 ( .A(n1231), .B(n1271), .ZN(n1303) );
XOR2_X1 U1030 ( .A(G128), .B(G146), .Z(n1271) );
INV_X1 U1031 ( .A(G143), .ZN(n1231) );
XOR2_X1 U1032 ( .A(n1324), .B(n1302), .Z(n1321) );
XOR2_X1 U1033 ( .A(G113), .B(G116), .Z(n1302) );
NAND2_X1 U1034 ( .A1(KEYINPUT8), .A2(n1301), .ZN(n1324) );
INV_X1 U1035 ( .A(G119), .ZN(n1301) );
INV_X1 U1036 ( .A(n1072), .ZN(n1242) );
XNOR2_X1 U1037 ( .A(n1105), .B(n1325), .ZN(n1072) );
NOR2_X1 U1038 ( .A1(n1106), .A2(KEYINPUT20), .ZN(n1325) );
AND2_X1 U1039 ( .A1(G217), .A2(n1266), .ZN(n1106) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1190), .ZN(n1266) );
INV_X1 U1041 ( .A(G902), .ZN(n1190) );
NAND2_X1 U1042 ( .A1(n1268), .A2(n1143), .ZN(n1105) );
XNOR2_X1 U1043 ( .A(n1326), .B(n1327), .ZN(n1143) );
XOR2_X1 U1044 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1045 ( .A(n1330), .B(n1331), .Z(n1329) );
NAND2_X1 U1046 ( .A1(KEYINPUT61), .A2(n1237), .ZN(n1331) );
NAND2_X1 U1047 ( .A1(n1332), .A2(n1333), .ZN(n1330) );
NAND2_X1 U1048 ( .A1(G110), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1049 ( .A(n1335), .B(KEYINPUT1), .Z(n1332) );
OR2_X1 U1050 ( .A1(n1334), .A2(G110), .ZN(n1335) );
XNOR2_X1 U1051 ( .A(n1336), .B(n1337), .ZN(n1334) );
NOR2_X1 U1052 ( .A1(KEYINPUT16), .A2(G128), .ZN(n1337) );
XNOR2_X1 U1053 ( .A(G119), .B(KEYINPUT24), .ZN(n1336) );
NOR2_X1 U1054 ( .A1(n1338), .A2(n1339), .ZN(n1328) );
INV_X1 U1055 ( .A(G221), .ZN(n1339) );
XOR2_X1 U1056 ( .A(n1340), .B(n1341), .Z(n1326) );
NOR2_X1 U1057 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1341) );
XNOR2_X1 U1058 ( .A(G137), .B(G125), .ZN(n1340) );
NAND2_X1 U1059 ( .A1(n1342), .A2(n1343), .ZN(n1067) );
OR3_X1 U1060 ( .A1(n1095), .A2(n1100), .A3(KEYINPUT44), .ZN(n1343) );
INV_X1 U1061 ( .A(n1344), .ZN(n1095) );
NAND2_X1 U1062 ( .A1(KEYINPUT44), .A2(n1155), .ZN(n1342) );
NOR2_X1 U1063 ( .A1(n1344), .A2(n1100), .ZN(n1155) );
XNOR2_X1 U1064 ( .A(n1345), .B(G478), .ZN(n1100) );
NAND2_X1 U1065 ( .A1(n1147), .A2(n1268), .ZN(n1345) );
XOR2_X1 U1066 ( .A(n1346), .B(n1347), .Z(n1147) );
NOR2_X1 U1067 ( .A1(n1338), .A2(n1348), .ZN(n1347) );
INV_X1 U1068 ( .A(G217), .ZN(n1348) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1057), .ZN(n1338) );
INV_X1 U1070 ( .A(G953), .ZN(n1057) );
NAND2_X1 U1071 ( .A1(n1349), .A2(n1350), .ZN(n1346) );
NAND2_X1 U1072 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1073 ( .A(KEYINPUT28), .B(n1353), .Z(n1349) );
NOR2_X1 U1074 ( .A1(n1351), .A2(n1352), .ZN(n1353) );
XOR2_X1 U1075 ( .A(n1354), .B(n1355), .Z(n1352) );
XOR2_X1 U1076 ( .A(G128), .B(n1356), .Z(n1355) );
NOR2_X1 U1077 ( .A1(KEYINPUT52), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1078 ( .A(G134), .B(KEYINPUT43), .ZN(n1357) );
XNOR2_X1 U1079 ( .A(G143), .B(KEYINPUT25), .ZN(n1354) );
XOR2_X1 U1080 ( .A(n1358), .B(n1277), .Z(n1351) );
XOR2_X1 U1081 ( .A(G107), .B(KEYINPUT23), .Z(n1277) );
XNOR2_X1 U1082 ( .A(G116), .B(G122), .ZN(n1358) );
XNOR2_X1 U1083 ( .A(n1359), .B(n1360), .ZN(n1344) );
XOR2_X1 U1084 ( .A(KEYINPUT34), .B(G475), .Z(n1360) );
NAND2_X1 U1085 ( .A1(n1151), .A2(n1268), .ZN(n1359) );
XNOR2_X1 U1086 ( .A(G902), .B(KEYINPUT19), .ZN(n1268) );
XOR2_X1 U1087 ( .A(n1361), .B(n1362), .Z(n1151) );
XOR2_X1 U1088 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1089 ( .A(G113), .B(n1281), .ZN(n1364) );
INV_X1 U1090 ( .A(G104), .ZN(n1281) );
XNOR2_X1 U1091 ( .A(G146), .B(n1251), .ZN(n1363) );
INV_X1 U1092 ( .A(G122), .ZN(n1251) );
XOR2_X1 U1093 ( .A(n1365), .B(n1121), .Z(n1361) );
XOR2_X1 U1094 ( .A(G125), .B(n1366), .Z(n1121) );
XNOR2_X1 U1095 ( .A(n1237), .B(G131), .ZN(n1366) );
INV_X1 U1096 ( .A(G140), .ZN(n1237) );
XOR2_X1 U1097 ( .A(n1367), .B(n1368), .Z(n1365) );
NOR2_X1 U1098 ( .A1(KEYINPUT5), .A2(G143), .ZN(n1368) );
NAND2_X1 U1099 ( .A1(G214), .A2(n1320), .ZN(n1367) );
NOR2_X1 U1100 ( .A1(G953), .A2(G237), .ZN(n1320) );
endmodule


