//Key = 0101011001001101010110100111001111011011100000110010000111011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337;

XNOR2_X1 U741 ( .A(G107), .B(n1015), .ZN(G9) );
NAND4_X1 U742 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1015) );
NOR3_X1 U743 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
XNOR2_X1 U744 ( .A(n1023), .B(KEYINPUT12), .ZN(n1018) );
NOR2_X1 U745 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND3_X1 U747 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1026) );
NAND2_X1 U748 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND3_X1 U752 ( .A1(n1023), .A2(n1040), .A3(n1017), .ZN(n1039) );
NAND4_X1 U753 ( .A1(n1041), .A2(n1040), .A3(n1042), .A4(n1043), .ZN(n1038) );
NAND2_X1 U754 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U755 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1042) );
NAND4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1017), .A4(n1051), .ZN(n1034) );
AND2_X1 U757 ( .A1(n1048), .A2(n1041), .ZN(n1051) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND2_X1 U759 ( .A1(n1040), .A2(n1054), .ZN(n1052) );
NAND2_X1 U760 ( .A1(n1021), .A2(n1055), .ZN(n1054) );
OR3_X1 U761 ( .A1(n1016), .A2(n1056), .A3(n1053), .ZN(n1049) );
INV_X1 U762 ( .A(n1057), .ZN(n1032) );
NOR3_X1 U763 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1024) );
INV_X1 U764 ( .A(n1029), .ZN(n1058) );
NAND4_X1 U765 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1029) );
NOR4_X1 U766 ( .A1(n1021), .A2(n1044), .A3(n1063), .A4(n1064), .ZN(n1062) );
XOR2_X1 U767 ( .A(n1065), .B(KEYINPUT47), .Z(n1063) );
NOR3_X1 U768 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1061) );
NOR2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U770 ( .A(n1071), .B(KEYINPUT44), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1072), .A2(n1073), .ZN(n1067) );
XNOR2_X1 U772 ( .A(n1071), .B(KEYINPUT25), .ZN(n1073) );
XOR2_X1 U773 ( .A(n1074), .B(n1075), .Z(G72) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1030), .ZN(n1077) );
AND2_X1 U776 ( .A1(G227), .A2(G900), .ZN(n1078) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NAND2_X1 U778 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1082), .B(n1083), .Z(n1079) );
XOR2_X1 U780 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U781 ( .A(G125), .B(n1086), .ZN(n1085) );
NOR2_X1 U782 ( .A1(KEYINPUT16), .A2(n1087), .ZN(n1086) );
XNOR2_X1 U783 ( .A(G134), .B(n1088), .ZN(n1087) );
NOR2_X1 U784 ( .A1(KEYINPUT54), .A2(n1089), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1084) );
XNOR2_X1 U786 ( .A(KEYINPUT8), .B(KEYINPUT10), .ZN(n1090) );
XOR2_X1 U787 ( .A(G131), .B(n1092), .Z(n1082) );
XOR2_X1 U788 ( .A(KEYINPUT15), .B(G140), .Z(n1092) );
NAND2_X1 U789 ( .A1(n1030), .A2(n1028), .ZN(n1074) );
NAND2_X1 U790 ( .A1(n1093), .A2(n1094), .ZN(G69) );
NAND2_X1 U791 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U792 ( .A1(G953), .A2(n1097), .ZN(n1095) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1097) );
NAND2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
NAND2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U796 ( .A1(G953), .A2(n1102), .ZN(n1101) );
INV_X1 U797 ( .A(n1103), .ZN(n1100) );
INV_X1 U798 ( .A(n1096), .ZN(n1098) );
NAND2_X1 U799 ( .A1(n1104), .A2(KEYINPUT1), .ZN(n1096) );
XOR2_X1 U800 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR3_X1 U801 ( .A1(n1103), .A2(n1107), .A3(n1108), .ZN(n1106) );
NOR2_X1 U802 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U803 ( .A(KEYINPUT52), .B(n1111), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1112), .A2(n1111), .ZN(n1107) );
NAND2_X1 U805 ( .A1(n1030), .A2(n1027), .ZN(n1105) );
NOR2_X1 U806 ( .A1(n1113), .A2(n1114), .ZN(G66) );
XOR2_X1 U807 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U808 ( .A1(n1117), .A2(G217), .ZN(n1115) );
NOR2_X1 U809 ( .A1(n1113), .A2(n1118), .ZN(G63) );
XOR2_X1 U810 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U811 ( .A1(n1117), .A2(G478), .ZN(n1119) );
NOR2_X1 U812 ( .A1(n1113), .A2(n1121), .ZN(G60) );
XOR2_X1 U813 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U814 ( .A1(n1117), .A2(G475), .ZN(n1122) );
XNOR2_X1 U815 ( .A(n1124), .B(n1125), .ZN(G6) );
NOR2_X1 U816 ( .A1(G104), .A2(KEYINPUT18), .ZN(n1125) );
NOR2_X1 U817 ( .A1(n1113), .A2(n1126), .ZN(G57) );
XOR2_X1 U818 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U819 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U820 ( .A1(n1131), .A2(KEYINPUT60), .ZN(n1129) );
XNOR2_X1 U821 ( .A(n1132), .B(n1133), .ZN(n1131) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(n1127) );
NOR2_X1 U823 ( .A1(KEYINPUT11), .A2(n1136), .ZN(n1135) );
XNOR2_X1 U824 ( .A(G101), .B(n1137), .ZN(n1134) );
NOR3_X1 U825 ( .A1(n1138), .A2(KEYINPUT14), .A3(n1139), .ZN(n1137) );
NOR2_X1 U826 ( .A1(n1113), .A2(n1140), .ZN(G54) );
XOR2_X1 U827 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U829 ( .A1(n1117), .A2(G469), .ZN(n1143) );
XOR2_X1 U830 ( .A(n1145), .B(KEYINPUT32), .Z(n1141) );
NAND2_X1 U831 ( .A1(KEYINPUT3), .A2(n1146), .ZN(n1145) );
XOR2_X1 U832 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U833 ( .A1(KEYINPUT28), .A2(n1133), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1113), .A2(n1149), .ZN(G51) );
NOR2_X1 U835 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U836 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U837 ( .A1(KEYINPUT9), .A2(n1154), .ZN(n1153) );
NAND2_X1 U838 ( .A1(n1117), .A2(n1155), .ZN(n1152) );
INV_X1 U839 ( .A(n1138), .ZN(n1117) );
NAND2_X1 U840 ( .A1(G902), .A2(n1156), .ZN(n1138) );
OR2_X1 U841 ( .A1(n1028), .A2(n1027), .ZN(n1156) );
NAND4_X1 U842 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1027) );
NOR4_X1 U843 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1124), .ZN(n1160) );
AND4_X1 U844 ( .A1(n1164), .A2(n1056), .A3(n1017), .A4(n1165), .ZN(n1124) );
OR2_X1 U845 ( .A1(n1166), .A2(KEYINPUT51), .ZN(n1159) );
NAND4_X1 U846 ( .A1(n1164), .A2(n1016), .A3(n1017), .A4(n1165), .ZN(n1158) );
NAND2_X1 U847 ( .A1(n1023), .A2(n1167), .ZN(n1157) );
NAND3_X1 U848 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
XNOR2_X1 U849 ( .A(KEYINPUT27), .B(n1171), .ZN(n1170) );
NAND3_X1 U850 ( .A1(KEYINPUT51), .A2(n1172), .A3(n1173), .ZN(n1169) );
NOR3_X1 U851 ( .A1(n1174), .A2(n1036), .A3(n1022), .ZN(n1173) );
XNOR2_X1 U852 ( .A(KEYINPUT19), .B(n1175), .ZN(n1168) );
NAND2_X1 U853 ( .A1(n1176), .A2(n1177), .ZN(n1028) );
NOR4_X1 U854 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR4_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1176) );
NOR2_X1 U856 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U857 ( .A(n1023), .B(KEYINPUT41), .ZN(n1186) );
INV_X1 U858 ( .A(n1188), .ZN(n1183) );
NOR2_X1 U859 ( .A1(KEYINPUT9), .A2(n1154), .ZN(n1150) );
XNOR2_X1 U860 ( .A(n1189), .B(n1190), .ZN(n1154) );
XNOR2_X1 U861 ( .A(n1132), .B(n1191), .ZN(n1190) );
XNOR2_X1 U862 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U863 ( .A1(KEYINPUT49), .A2(n1194), .ZN(n1193) );
NAND2_X1 U864 ( .A1(KEYINPUT39), .A2(n1195), .ZN(n1192) );
XNOR2_X1 U865 ( .A(n1196), .B(n1197), .ZN(n1189) );
XOR2_X1 U866 ( .A(KEYINPUT24), .B(KEYINPUT2), .Z(n1197) );
NOR2_X1 U867 ( .A1(n1030), .A2(G952), .ZN(n1113) );
XNOR2_X1 U868 ( .A(n1198), .B(n1184), .ZN(G48) );
AND2_X1 U869 ( .A1(n1199), .A2(n1056), .ZN(n1184) );
XNOR2_X1 U870 ( .A(G143), .B(n1188), .ZN(G45) );
NAND3_X1 U871 ( .A1(n1172), .A2(n1164), .A3(n1200), .ZN(n1188) );
NOR3_X1 U872 ( .A1(n1201), .A2(n1202), .A3(n1059), .ZN(n1200) );
XOR2_X1 U873 ( .A(G140), .B(n1178), .Z(G42) );
AND3_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1056), .ZN(n1178) );
XOR2_X1 U875 ( .A(n1205), .B(n1182), .Z(G39) );
AND2_X1 U876 ( .A1(n1206), .A2(n1204), .ZN(n1182) );
XNOR2_X1 U877 ( .A(G137), .B(KEYINPUT5), .ZN(n1205) );
XNOR2_X1 U878 ( .A(n1207), .B(n1181), .ZN(G36) );
AND3_X1 U879 ( .A1(n1204), .A2(n1016), .A3(n1172), .ZN(n1181) );
XNOR2_X1 U880 ( .A(n1180), .B(n1208), .ZN(G33) );
NAND2_X1 U881 ( .A1(KEYINPUT17), .A2(G131), .ZN(n1208) );
AND3_X1 U882 ( .A1(n1056), .A2(n1204), .A3(n1172), .ZN(n1180) );
AND3_X1 U883 ( .A1(n1041), .A2(n1055), .A3(n1209), .ZN(n1204) );
NOR3_X1 U884 ( .A1(n1202), .A2(n1021), .A3(n1044), .ZN(n1209) );
INV_X1 U885 ( .A(n1210), .ZN(n1202) );
XOR2_X1 U886 ( .A(n1211), .B(KEYINPUT55), .Z(n1041) );
XOR2_X1 U887 ( .A(G128), .B(n1179), .Z(G30) );
AND2_X1 U888 ( .A1(n1199), .A2(n1016), .ZN(n1179) );
AND4_X1 U889 ( .A1(n1164), .A2(n1212), .A3(n1210), .A4(n1213), .ZN(n1199) );
NAND2_X1 U890 ( .A1(n1214), .A2(n1215), .ZN(G3) );
NAND2_X1 U891 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U892 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND2_X1 U893 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
OR2_X1 U894 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
INV_X1 U895 ( .A(KEYINPUT50), .ZN(n1221) );
NAND2_X1 U896 ( .A1(G101), .A2(n1222), .ZN(n1214) );
NOR2_X1 U897 ( .A1(n1163), .A2(KEYINPUT48), .ZN(n1222) );
INV_X1 U898 ( .A(n1220), .ZN(n1163) );
NAND2_X1 U899 ( .A1(n1223), .A2(n1172), .ZN(n1220) );
XNOR2_X1 U900 ( .A(n1224), .B(n1225), .ZN(G27) );
NOR2_X1 U901 ( .A1(n1226), .A2(n1187), .ZN(n1225) );
NAND4_X1 U902 ( .A1(n1036), .A2(n1056), .A3(n1203), .A4(n1210), .ZN(n1187) );
NAND2_X1 U903 ( .A1(n1057), .A2(n1227), .ZN(n1210) );
NAND4_X1 U904 ( .A1(G902), .A2(G953), .A3(n1228), .A4(n1081), .ZN(n1227) );
INV_X1 U905 ( .A(G900), .ZN(n1081) );
XOR2_X1 U906 ( .A(G122), .B(n1229), .Z(G24) );
NOR2_X1 U907 ( .A1(n1226), .A2(n1171), .ZN(n1229) );
NAND4_X1 U908 ( .A1(n1230), .A2(n1017), .A3(n1231), .A4(n1232), .ZN(n1171) );
INV_X1 U909 ( .A(n1045), .ZN(n1017) );
NAND2_X1 U910 ( .A1(n1060), .A2(n1233), .ZN(n1045) );
XOR2_X1 U911 ( .A(G119), .B(n1162), .Z(G21) );
AND3_X1 U912 ( .A1(n1206), .A2(n1023), .A3(n1230), .ZN(n1162) );
AND3_X1 U913 ( .A1(n1212), .A2(n1213), .A3(n1040), .ZN(n1206) );
XNOR2_X1 U914 ( .A(G116), .B(n1166), .ZN(G18) );
NAND4_X1 U915 ( .A1(n1230), .A2(n1172), .A3(n1016), .A4(n1023), .ZN(n1166) );
INV_X1 U916 ( .A(n1174), .ZN(n1016) );
NAND2_X1 U917 ( .A1(n1231), .A2(n1234), .ZN(n1174) );
XNOR2_X1 U918 ( .A(n1235), .B(n1232), .ZN(n1234) );
XOR2_X1 U919 ( .A(G113), .B(n1236), .Z(G15) );
NOR2_X1 U920 ( .A1(n1226), .A2(n1175), .ZN(n1236) );
NAND3_X1 U921 ( .A1(n1172), .A2(n1056), .A3(n1230), .ZN(n1175) );
NOR2_X1 U922 ( .A1(n1053), .A2(n1022), .ZN(n1230) );
INV_X1 U923 ( .A(n1165), .ZN(n1022) );
INV_X1 U924 ( .A(n1036), .ZN(n1053) );
NOR2_X1 U925 ( .A1(n1055), .A2(n1021), .ZN(n1036) );
INV_X1 U926 ( .A(n1046), .ZN(n1172) );
NAND2_X1 U927 ( .A1(n1060), .A2(n1212), .ZN(n1046) );
XNOR2_X1 U928 ( .A(n1237), .B(KEYINPUT57), .ZN(n1212) );
INV_X1 U929 ( .A(n1213), .ZN(n1060) );
XNOR2_X1 U930 ( .A(n1238), .B(n1161), .ZN(G12) );
AND2_X1 U931 ( .A1(n1223), .A2(n1203), .ZN(n1161) );
INV_X1 U932 ( .A(n1047), .ZN(n1203) );
NAND2_X1 U933 ( .A1(n1233), .A2(n1213), .ZN(n1047) );
NAND3_X1 U934 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1213) );
OR2_X1 U935 ( .A1(n1242), .A2(n1116), .ZN(n1241) );
NAND3_X1 U936 ( .A1(n1116), .A2(n1242), .A3(n1243), .ZN(n1240) );
NAND2_X1 U937 ( .A1(G217), .A2(n1244), .ZN(n1242) );
XOR2_X1 U938 ( .A(n1245), .B(n1246), .Z(n1116) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U940 ( .A(n1249), .B(n1250), .Z(n1248) );
NOR2_X1 U941 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U942 ( .A(KEYINPUT59), .B(G221), .Z(n1252) );
INV_X1 U943 ( .A(n1253), .ZN(n1251) );
NOR2_X1 U944 ( .A1(G137), .A2(KEYINPUT23), .ZN(n1249) );
XNOR2_X1 U945 ( .A(KEYINPUT43), .B(n1224), .ZN(n1247) );
XOR2_X1 U946 ( .A(n1254), .B(n1255), .Z(n1245) );
XNOR2_X1 U947 ( .A(n1256), .B(n1257), .ZN(n1254) );
NOR2_X1 U948 ( .A1(G119), .A2(KEYINPUT58), .ZN(n1257) );
NAND2_X1 U949 ( .A1(G902), .A2(G217), .ZN(n1239) );
XNOR2_X1 U950 ( .A(KEYINPUT34), .B(n1237), .ZN(n1233) );
XOR2_X1 U951 ( .A(n1065), .B(KEYINPUT22), .Z(n1237) );
XNOR2_X1 U952 ( .A(n1258), .B(n1139), .ZN(n1065) );
INV_X1 U953 ( .A(G472), .ZN(n1139) );
NAND2_X1 U954 ( .A1(n1259), .A2(n1243), .ZN(n1258) );
XNOR2_X1 U955 ( .A(n1136), .B(n1260), .ZN(n1259) );
XNOR2_X1 U956 ( .A(n1217), .B(n1261), .ZN(n1260) );
NOR2_X1 U957 ( .A1(KEYINPUT53), .A2(n1262), .ZN(n1261) );
XOR2_X1 U958 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U959 ( .A(n1130), .B(n1133), .ZN(n1264) );
XNOR2_X1 U960 ( .A(n1265), .B(KEYINPUT4), .ZN(n1263) );
NAND2_X1 U961 ( .A1(KEYINPUT61), .A2(n1132), .ZN(n1265) );
NAND3_X1 U962 ( .A1(n1266), .A2(n1030), .A3(G210), .ZN(n1136) );
AND3_X1 U963 ( .A1(n1040), .A2(n1165), .A3(n1164), .ZN(n1223) );
NOR3_X1 U964 ( .A1(n1020), .A2(n1021), .A3(n1226), .ZN(n1164) );
INV_X1 U965 ( .A(n1023), .ZN(n1226) );
NOR2_X1 U966 ( .A1(n1267), .A2(n1044), .ZN(n1023) );
INV_X1 U967 ( .A(n1048), .ZN(n1044) );
NAND2_X1 U968 ( .A1(G214), .A2(n1268), .ZN(n1048) );
INV_X1 U969 ( .A(n1211), .ZN(n1267) );
XOR2_X1 U970 ( .A(n1066), .B(KEYINPUT7), .Z(n1211) );
XOR2_X1 U971 ( .A(n1155), .B(n1269), .Z(n1066) );
NOR2_X1 U972 ( .A1(G902), .A2(n1270), .ZN(n1269) );
XOR2_X1 U973 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U974 ( .A(n1195), .B(n1273), .Z(n1272) );
NOR2_X1 U975 ( .A1(n1196), .A2(KEYINPUT42), .ZN(n1273) );
AND2_X1 U976 ( .A1(n1274), .A2(n1275), .ZN(n1196) );
NAND3_X1 U977 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1275) );
XNOR2_X1 U978 ( .A(n1279), .B(KEYINPUT36), .ZN(n1278) );
XNOR2_X1 U979 ( .A(KEYINPUT38), .B(n1280), .ZN(n1276) );
NAND3_X1 U980 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1274) );
XNOR2_X1 U981 ( .A(KEYINPUT36), .B(n1111), .ZN(n1283) );
INV_X1 U982 ( .A(n1279), .ZN(n1111) );
XOR2_X1 U983 ( .A(G110), .B(n1284), .Z(n1279) );
OR2_X1 U984 ( .A1(n1280), .A2(KEYINPUT38), .ZN(n1282) );
NAND2_X1 U985 ( .A1(n1109), .A2(KEYINPUT38), .ZN(n1281) );
INV_X1 U986 ( .A(n1112), .ZN(n1109) );
NAND2_X1 U987 ( .A1(n1277), .A2(n1280), .ZN(n1112) );
OR2_X1 U988 ( .A1(n1130), .A2(n1285), .ZN(n1280) );
NAND2_X1 U989 ( .A1(n1285), .A2(n1130), .ZN(n1277) );
XOR2_X1 U990 ( .A(G113), .B(n1286), .Z(n1130) );
XNOR2_X1 U991 ( .A(G119), .B(n1287), .ZN(n1286) );
INV_X1 U992 ( .A(G116), .ZN(n1287) );
XOR2_X1 U993 ( .A(n1288), .B(n1289), .Z(n1285) );
XNOR2_X1 U994 ( .A(G104), .B(G107), .ZN(n1288) );
NOR2_X1 U995 ( .A1(n1102), .A2(G953), .ZN(n1195) );
INV_X1 U996 ( .A(G224), .ZN(n1102) );
XOR2_X1 U997 ( .A(n1132), .B(n1194), .Z(n1271) );
XNOR2_X1 U998 ( .A(n1224), .B(KEYINPUT29), .ZN(n1194) );
XNOR2_X1 U999 ( .A(n1290), .B(n1291), .ZN(n1132) );
INV_X1 U1000 ( .A(n1256), .ZN(n1291) );
NAND2_X1 U1001 ( .A1(KEYINPUT30), .A2(n1292), .ZN(n1290) );
AND2_X1 U1002 ( .A1(G210), .A2(n1268), .ZN(n1155) );
NAND2_X1 U1003 ( .A1(n1266), .A2(n1243), .ZN(n1268) );
AND2_X1 U1004 ( .A1(G221), .A2(n1293), .ZN(n1021) );
NAND2_X1 U1005 ( .A1(G234), .A2(n1243), .ZN(n1293) );
INV_X1 U1006 ( .A(n1055), .ZN(n1020) );
XOR2_X1 U1007 ( .A(n1294), .B(n1295), .Z(n1055) );
INV_X1 U1008 ( .A(n1071), .ZN(n1295) );
XOR2_X1 U1009 ( .A(G469), .B(KEYINPUT63), .Z(n1071) );
XNOR2_X1 U1010 ( .A(n1072), .B(KEYINPUT13), .ZN(n1294) );
INV_X1 U1011 ( .A(n1069), .ZN(n1072) );
NAND2_X1 U1012 ( .A1(n1296), .A2(n1243), .ZN(n1069) );
XNOR2_X1 U1013 ( .A(n1297), .B(n1133), .ZN(n1296) );
XNOR2_X1 U1014 ( .A(G131), .B(n1298), .ZN(n1133) );
NOR2_X1 U1015 ( .A1(KEYINPUT37), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U1016 ( .A(n1089), .B(n1300), .ZN(n1299) );
NOR2_X1 U1017 ( .A1(G134), .A2(KEYINPUT21), .ZN(n1300) );
INV_X1 U1018 ( .A(G137), .ZN(n1089) );
XNOR2_X1 U1019 ( .A(n1148), .B(n1301), .ZN(n1297) );
NOR2_X1 U1020 ( .A1(KEYINPUT0), .A2(n1144), .ZN(n1301) );
XOR2_X1 U1021 ( .A(n1302), .B(n1255), .Z(n1144) );
XNOR2_X1 U1022 ( .A(n1238), .B(G140), .ZN(n1255) );
NAND2_X1 U1023 ( .A1(G227), .A2(n1030), .ZN(n1302) );
XNOR2_X1 U1024 ( .A(n1091), .B(n1303), .ZN(n1148) );
XOR2_X1 U1025 ( .A(n1304), .B(n1305), .Z(n1303) );
NAND2_X1 U1026 ( .A1(KEYINPUT31), .A2(n1289), .ZN(n1305) );
XNOR2_X1 U1027 ( .A(n1217), .B(KEYINPUT56), .ZN(n1289) );
INV_X1 U1028 ( .A(G101), .ZN(n1217) );
NAND2_X1 U1029 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NAND2_X1 U1030 ( .A1(G107), .A2(n1308), .ZN(n1307) );
XOR2_X1 U1031 ( .A(KEYINPUT40), .B(n1309), .Z(n1306) );
NOR2_X1 U1032 ( .A1(G107), .A2(n1308), .ZN(n1309) );
INV_X1 U1033 ( .A(G104), .ZN(n1308) );
XNOR2_X1 U1034 ( .A(n1256), .B(G143), .ZN(n1091) );
XOR2_X1 U1035 ( .A(G146), .B(n1310), .Z(n1256) );
NAND2_X1 U1036 ( .A1(n1057), .A2(n1311), .ZN(n1165) );
NAND3_X1 U1037 ( .A1(n1103), .A2(n1228), .A3(G902), .ZN(n1311) );
NOR2_X1 U1038 ( .A1(n1030), .A2(G898), .ZN(n1103) );
NAND3_X1 U1039 ( .A1(n1228), .A2(n1030), .A3(G952), .ZN(n1057) );
NAND2_X1 U1040 ( .A1(G237), .A2(G234), .ZN(n1228) );
NAND2_X1 U1041 ( .A1(n1312), .A2(n1313), .ZN(n1040) );
NAND2_X1 U1042 ( .A1(n1056), .A2(n1235), .ZN(n1313) );
INV_X1 U1043 ( .A(KEYINPUT35), .ZN(n1235) );
NOR2_X1 U1044 ( .A1(n1059), .A2(n1231), .ZN(n1056) );
INV_X1 U1045 ( .A(n1201), .ZN(n1231) );
NAND3_X1 U1046 ( .A1(n1201), .A2(n1059), .A3(KEYINPUT35), .ZN(n1312) );
INV_X1 U1047 ( .A(n1232), .ZN(n1059) );
XNOR2_X1 U1048 ( .A(n1314), .B(G475), .ZN(n1232) );
NAND2_X1 U1049 ( .A1(n1123), .A2(n1243), .ZN(n1314) );
XNOR2_X1 U1050 ( .A(n1315), .B(n1316), .ZN(n1123) );
XOR2_X1 U1051 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1052 ( .A(n1224), .B(G113), .ZN(n1318) );
INV_X1 U1053 ( .A(G125), .ZN(n1224) );
XNOR2_X1 U1054 ( .A(n1198), .B(G131), .ZN(n1317) );
INV_X1 U1055 ( .A(G146), .ZN(n1198) );
XOR2_X1 U1056 ( .A(n1319), .B(n1320), .Z(n1315) );
XOR2_X1 U1057 ( .A(n1321), .B(n1284), .Z(n1320) );
NOR2_X1 U1058 ( .A1(G140), .A2(KEYINPUT62), .ZN(n1321) );
XNOR2_X1 U1059 ( .A(G104), .B(n1322), .ZN(n1319) );
NOR2_X1 U1060 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1061 ( .A(n1325), .B(KEYINPUT26), .Z(n1324) );
NAND2_X1 U1062 ( .A1(n1292), .A2(n1326), .ZN(n1325) );
NOR2_X1 U1063 ( .A1(n1292), .A2(n1326), .ZN(n1323) );
NAND3_X1 U1064 ( .A1(n1266), .A2(n1030), .A3(G214), .ZN(n1326) );
INV_X1 U1065 ( .A(G953), .ZN(n1030) );
INV_X1 U1066 ( .A(G237), .ZN(n1266) );
INV_X1 U1067 ( .A(G143), .ZN(n1292) );
XOR2_X1 U1068 ( .A(n1064), .B(KEYINPUT33), .Z(n1201) );
XNOR2_X1 U1069 ( .A(n1327), .B(G478), .ZN(n1064) );
NAND2_X1 U1070 ( .A1(n1120), .A2(n1243), .ZN(n1327) );
INV_X1 U1071 ( .A(G902), .ZN(n1243) );
XOR2_X1 U1072 ( .A(n1328), .B(n1329), .Z(n1120) );
XOR2_X1 U1073 ( .A(n1330), .B(n1331), .Z(n1329) );
NAND2_X1 U1074 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1075 ( .A1(G143), .A2(n1310), .ZN(n1333) );
XOR2_X1 U1076 ( .A(n1334), .B(KEYINPUT45), .Z(n1332) );
OR2_X1 U1077 ( .A1(n1310), .A2(G143), .ZN(n1334) );
XOR2_X1 U1078 ( .A(G128), .B(KEYINPUT20), .Z(n1310) );
NAND2_X1 U1079 ( .A1(n1335), .A2(KEYINPUT46), .ZN(n1330) );
XNOR2_X1 U1080 ( .A(G116), .B(n1284), .ZN(n1335) );
XOR2_X1 U1081 ( .A(G122), .B(KEYINPUT6), .Z(n1284) );
XOR2_X1 U1082 ( .A(n1336), .B(n1337), .Z(n1328) );
XNOR2_X1 U1083 ( .A(n1207), .B(G107), .ZN(n1337) );
INV_X1 U1084 ( .A(G134), .ZN(n1207) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1253), .ZN(n1336) );
NOR2_X1 U1086 ( .A1(n1244), .A2(G953), .ZN(n1253) );
INV_X1 U1087 ( .A(G234), .ZN(n1244) );
INV_X1 U1088 ( .A(G110), .ZN(n1238) );
endmodule


