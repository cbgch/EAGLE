//Key = 0110010110100110101111001100001100011011101000101001101000000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;

XOR2_X1 U745 ( .A(n1035), .B(n1036), .Z(G9) );
XNOR2_X1 U746 ( .A(G107), .B(KEYINPUT9), .ZN(n1036) );
NAND3_X1 U747 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1035) );
NOR3_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
XOR2_X1 U749 ( .A(n1043), .B(KEYINPUT25), .Z(n1041) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U751 ( .A1(G953), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
NOR2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR3_X1 U754 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NOR3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1054) );
NOR2_X1 U756 ( .A1(n1040), .A2(n1059), .ZN(n1058) );
NOR3_X1 U757 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1057) );
XOR2_X1 U758 ( .A(n1059), .B(KEYINPUT34), .Z(n1061) );
NAND3_X1 U759 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1056) );
NAND3_X1 U760 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND3_X1 U761 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT56), .ZN(n1064) );
NAND2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1063) );
INV_X1 U763 ( .A(KEYINPUT56), .ZN(n1072) );
NOR3_X1 U764 ( .A1(n1070), .A2(n1073), .A3(n1059), .ZN(n1051) );
NOR2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1053), .ZN(n1075) );
NOR2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U768 ( .A1(n1079), .A2(n1055), .ZN(n1074) );
NOR2_X1 U769 ( .A1(n1037), .A2(n1080), .ZN(n1079) );
NOR3_X1 U770 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1044) );
AND4_X1 U771 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1046) );
NOR4_X1 U772 ( .A1(n1085), .A2(n1068), .A3(n1086), .A4(n1087), .ZN(n1084) );
XOR2_X1 U773 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U774 ( .A(KEYINPUT18), .B(n1090), .Z(n1089) );
XNOR2_X1 U775 ( .A(n1091), .B(n1092), .ZN(n1086) );
NAND2_X1 U776 ( .A1(KEYINPUT31), .A2(n1093), .ZN(n1091) );
INV_X1 U777 ( .A(n1094), .ZN(n1068) );
XNOR2_X1 U778 ( .A(G472), .B(n1095), .ZN(n1083) );
NAND2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(G72) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U781 ( .A(n1100), .B(n1101), .ZN(n1099) );
XOR2_X1 U782 ( .A(KEYINPUT52), .B(n1102), .Z(n1098) );
XOR2_X1 U783 ( .A(n1103), .B(KEYINPUT55), .Z(n1096) );
NAND2_X1 U784 ( .A1(n1104), .A2(n1102), .ZN(n1103) );
AND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND2_X1 U786 ( .A1(G900), .A2(G227), .ZN(n1106) );
XOR2_X1 U787 ( .A(KEYINPUT57), .B(G953), .Z(n1105) );
XOR2_X1 U788 ( .A(n1101), .B(n1100), .Z(n1104) );
AND2_X1 U789 ( .A1(n1107), .A2(n1108), .ZN(n1100) );
NAND2_X1 U790 ( .A1(G953), .A2(n1109), .ZN(n1108) );
XOR2_X1 U791 ( .A(KEYINPUT36), .B(G900), .Z(n1109) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(n1107) );
XOR2_X1 U793 ( .A(KEYINPUT1), .B(G140), .Z(n1111) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1110) );
NAND3_X1 U795 ( .A1(KEYINPUT2), .A2(n1114), .A3(n1115), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1116), .B(KEYINPUT60), .Z(n1115) );
OR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
XNOR2_X1 U799 ( .A(n1119), .B(n1120), .ZN(n1117) );
NOR2_X1 U800 ( .A1(G134), .A2(KEYINPUT26), .ZN(n1120) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1101) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(G69) );
XOR2_X1 U803 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U804 ( .A1(n1127), .A2(n1121), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U807 ( .A1(KEYINPUT37), .A2(n1132), .ZN(n1131) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1133), .ZN(n1128) );
XOR2_X1 U809 ( .A(KEYINPUT47), .B(G898), .Z(n1133) );
NOR2_X1 U810 ( .A1(n1134), .A2(n1121), .ZN(n1123) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(G66) );
NOR3_X1 U813 ( .A1(n1090), .A2(n1139), .A3(n1140), .ZN(n1138) );
NOR3_X1 U814 ( .A1(n1141), .A2(n1088), .A3(n1142), .ZN(n1140) );
NOR2_X1 U815 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NOR2_X1 U816 ( .A1(n1145), .A2(n1088), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1137), .A2(n1146), .ZN(G63) );
NOR2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U819 ( .A(n1149), .B(KEYINPUT13), .Z(n1148) );
NAND2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
AND2_X1 U822 ( .A1(n1152), .A2(G478), .ZN(n1150) );
NOR3_X1 U823 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(G60) );
AND2_X1 U824 ( .A1(KEYINPUT62), .A2(n1137), .ZN(n1155) );
NOR3_X1 U825 ( .A1(KEYINPUT62), .A2(G953), .A3(G952), .ZN(n1154) );
XNOR2_X1 U826 ( .A(n1156), .B(n1157), .ZN(n1153) );
AND2_X1 U827 ( .A1(G475), .A2(n1152), .ZN(n1157) );
XNOR2_X1 U828 ( .A(G104), .B(n1158), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1137), .A2(n1159), .ZN(G57) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U831 ( .A(n1162), .B(n1163), .ZN(n1161) );
NAND2_X1 U832 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U833 ( .A1(KEYINPUT14), .A2(n1166), .ZN(n1165) );
OR2_X1 U834 ( .A1(KEYINPUT46), .A2(n1166), .ZN(n1164) );
AND2_X1 U835 ( .A1(n1152), .A2(G472), .ZN(n1166) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1160) );
INV_X1 U837 ( .A(n1169), .ZN(n1168) );
NOR2_X1 U838 ( .A1(n1137), .A2(n1170), .ZN(G54) );
XOR2_X1 U839 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U840 ( .A(n1173), .B(n1169), .Z(n1172) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1169) );
NAND2_X1 U842 ( .A1(n1176), .A2(KEYINPUT51), .ZN(n1173) );
XOR2_X1 U843 ( .A(n1177), .B(G101), .Z(n1176) );
XOR2_X1 U844 ( .A(n1178), .B(n1179), .Z(n1171) );
NOR3_X1 U845 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NOR2_X1 U846 ( .A1(KEYINPUT54), .A2(n1183), .ZN(n1182) );
NOR3_X1 U847 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1181) );
INV_X1 U848 ( .A(KEYINPUT54), .ZN(n1184) );
AND2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1180) );
NAND2_X1 U850 ( .A1(KEYINPUT35), .A2(n1183), .ZN(n1186) );
XOR2_X1 U851 ( .A(G140), .B(G110), .Z(n1183) );
NAND3_X1 U852 ( .A1(n1187), .A2(n1188), .A3(G469), .ZN(n1178) );
OR2_X1 U853 ( .A1(n1152), .A2(KEYINPUT50), .ZN(n1188) );
INV_X1 U854 ( .A(n1142), .ZN(n1152) );
NAND2_X1 U855 ( .A1(KEYINPUT50), .A2(n1189), .ZN(n1187) );
NAND2_X1 U856 ( .A1(n1145), .A2(G902), .ZN(n1189) );
NOR2_X1 U857 ( .A1(n1137), .A2(n1190), .ZN(G51) );
XOR2_X1 U858 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U859 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND2_X1 U860 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U861 ( .A1(n1113), .A2(n1197), .ZN(n1196) );
INV_X1 U862 ( .A(KEYINPUT28), .ZN(n1197) );
NAND3_X1 U863 ( .A1(G125), .A2(n1175), .A3(KEYINPUT28), .ZN(n1195) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1191) );
NOR2_X1 U865 ( .A1(n1092), .A2(n1142), .ZN(n1199) );
NAND2_X1 U866 ( .A1(G902), .A2(n1048), .ZN(n1142) );
INV_X1 U867 ( .A(n1145), .ZN(n1048) );
NOR2_X1 U868 ( .A1(n1122), .A2(n1127), .ZN(n1145) );
NAND4_X1 U869 ( .A1(n1200), .A2(n1158), .A3(n1201), .A4(n1202), .ZN(n1127) );
AND4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR3_X1 U871 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1201) );
NOR2_X1 U872 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
INV_X1 U873 ( .A(KEYINPUT42), .ZN(n1210) );
NOR3_X1 U874 ( .A1(KEYINPUT42), .A2(n1212), .A3(n1213), .ZN(n1208) );
NOR2_X1 U875 ( .A1(n1070), .A2(n1214), .ZN(n1207) );
NAND3_X1 U876 ( .A1(n1080), .A2(n1038), .A3(n1215), .ZN(n1158) );
NAND3_X1 U877 ( .A1(n1037), .A2(n1038), .A3(n1215), .ZN(n1200) );
NAND4_X1 U878 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1122) );
NOR4_X1 U879 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
NOR2_X1 U880 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
INV_X1 U881 ( .A(n1226), .ZN(n1225) );
NOR3_X1 U882 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1224) );
NOR2_X1 U883 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1232), .B(KEYINPUT29), .Z(n1230) );
NOR2_X1 U885 ( .A1(n1053), .A2(n1233), .ZN(n1227) );
AND2_X1 U886 ( .A1(KEYINPUT39), .A2(n1234), .ZN(n1221) );
NOR3_X1 U887 ( .A1(KEYINPUT39), .A2(n1080), .A3(n1235), .ZN(n1220) );
NOR2_X1 U888 ( .A1(n1121), .A2(G952), .ZN(n1137) );
XOR2_X1 U889 ( .A(G146), .B(n1222), .Z(G48) );
AND3_X1 U890 ( .A1(n1236), .A2(n1237), .A3(n1080), .ZN(n1222) );
XNOR2_X1 U891 ( .A(G143), .B(n1218), .ZN(G45) );
NAND4_X1 U892 ( .A1(n1077), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1218) );
INV_X1 U893 ( .A(n1240), .ZN(n1238) );
XOR2_X1 U894 ( .A(n1241), .B(n1242), .Z(G42) );
NAND3_X1 U895 ( .A1(n1080), .A2(n1226), .A3(n1078), .ZN(n1242) );
XOR2_X1 U896 ( .A(n1119), .B(n1243), .Z(G39) );
NAND3_X1 U897 ( .A1(n1226), .A2(n1082), .A3(n1244), .ZN(n1243) );
XOR2_X1 U898 ( .A(n1233), .B(KEYINPUT8), .Z(n1244) );
XNOR2_X1 U899 ( .A(G134), .B(n1216), .ZN(G36) );
NAND3_X1 U900 ( .A1(n1226), .A2(n1037), .A3(n1077), .ZN(n1216) );
XOR2_X1 U901 ( .A(n1118), .B(n1245), .Z(G33) );
NAND3_X1 U902 ( .A1(n1246), .A2(n1247), .A3(n1228), .ZN(n1245) );
OR2_X1 U903 ( .A1(n1226), .A2(KEYINPUT49), .ZN(n1247) );
NOR3_X1 U904 ( .A1(n1040), .A2(n1248), .A3(n1059), .ZN(n1226) );
NAND2_X1 U905 ( .A1(KEYINPUT49), .A2(n1249), .ZN(n1246) );
NAND3_X1 U906 ( .A1(n1059), .A2(n1250), .A3(n1251), .ZN(n1249) );
INV_X1 U907 ( .A(n1040), .ZN(n1251) );
NAND2_X1 U908 ( .A1(n1252), .A2(n1094), .ZN(n1059) );
XOR2_X1 U909 ( .A(n1066), .B(KEYINPUT12), .Z(n1252) );
XOR2_X1 U910 ( .A(n1253), .B(n1217), .Z(G30) );
NAND3_X1 U911 ( .A1(n1237), .A2(n1037), .A3(n1236), .ZN(n1217) );
NOR3_X1 U912 ( .A1(n1213), .A2(n1248), .A3(n1040), .ZN(n1237) );
INV_X1 U913 ( .A(n1250), .ZN(n1248) );
XOR2_X1 U914 ( .A(n1254), .B(n1206), .Z(G3) );
NAND3_X1 U915 ( .A1(n1077), .A2(n1082), .A3(n1215), .ZN(n1206) );
XOR2_X1 U916 ( .A(G125), .B(n1234), .Z(G27) );
NOR2_X1 U917 ( .A1(n1235), .A2(n1232), .ZN(n1234) );
NAND3_X1 U918 ( .A1(n1078), .A2(n1250), .A3(n1071), .ZN(n1235) );
NAND2_X1 U919 ( .A1(n1050), .A2(n1255), .ZN(n1250) );
NAND4_X1 U920 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1257), .ZN(n1255) );
INV_X1 U921 ( .A(G900), .ZN(n1257) );
NAND2_X1 U922 ( .A1(n1258), .A2(n1259), .ZN(G24) );
NAND2_X1 U923 ( .A1(G122), .A2(n1211), .ZN(n1259) );
NAND2_X1 U924 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
XNOR2_X1 U925 ( .A(KEYINPUT32), .B(n1211), .ZN(n1261) );
NAND2_X1 U926 ( .A1(n1212), .A2(n1069), .ZN(n1211) );
INV_X1 U927 ( .A(n1213), .ZN(n1069) );
AND3_X1 U928 ( .A1(n1067), .A2(n1038), .A3(n1262), .ZN(n1212) );
NOR3_X1 U929 ( .A1(n1240), .A2(n1263), .A3(n1264), .ZN(n1262) );
INV_X1 U930 ( .A(n1055), .ZN(n1038) );
NAND2_X1 U931 ( .A1(n1265), .A2(n1266), .ZN(n1055) );
INV_X1 U932 ( .A(n1267), .ZN(n1266) );
INV_X1 U933 ( .A(n1070), .ZN(n1067) );
XOR2_X1 U934 ( .A(KEYINPUT40), .B(G122), .Z(n1260) );
XNOR2_X1 U935 ( .A(G119), .B(n1205), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1071), .A2(n1236), .A3(n1082), .A4(n1043), .ZN(n1205) );
INV_X1 U937 ( .A(n1233), .ZN(n1236) );
NAND2_X1 U938 ( .A1(n1267), .A2(n1268), .ZN(n1233) );
XNOR2_X1 U939 ( .A(G116), .B(n1204), .ZN(G18) );
NAND4_X1 U940 ( .A1(n1071), .A2(n1077), .A3(n1037), .A4(n1043), .ZN(n1204) );
NOR2_X1 U941 ( .A1(n1239), .A2(n1240), .ZN(n1037) );
NOR2_X1 U942 ( .A1(n1070), .A2(n1213), .ZN(n1071) );
XOR2_X1 U943 ( .A(n1042), .B(KEYINPUT11), .Z(n1213) );
XOR2_X1 U944 ( .A(G113), .B(n1269), .Z(G15) );
NOR2_X1 U945 ( .A1(n1270), .A2(n1214), .ZN(n1269) );
NAND3_X1 U946 ( .A1(n1271), .A2(n1043), .A3(n1228), .ZN(n1214) );
AND2_X1 U947 ( .A1(n1080), .A2(n1077), .ZN(n1228) );
NOR2_X1 U948 ( .A1(n1265), .A2(n1267), .ZN(n1077) );
INV_X1 U949 ( .A(n1232), .ZN(n1080) );
NAND2_X1 U950 ( .A1(n1240), .A2(n1239), .ZN(n1232) );
INV_X1 U951 ( .A(n1264), .ZN(n1239) );
INV_X1 U952 ( .A(n1042), .ZN(n1271) );
XOR2_X1 U953 ( .A(n1070), .B(KEYINPUT22), .Z(n1270) );
NAND2_X1 U954 ( .A1(n1081), .A2(n1272), .ZN(n1070) );
XOR2_X1 U955 ( .A(n1273), .B(n1203), .Z(G12) );
NAND3_X1 U956 ( .A1(n1078), .A2(n1082), .A3(n1215), .ZN(n1203) );
NOR3_X1 U957 ( .A1(n1042), .A2(n1263), .A3(n1040), .ZN(n1215) );
NAND2_X1 U958 ( .A1(n1060), .A2(n1272), .ZN(n1040) );
XOR2_X1 U959 ( .A(n1085), .B(KEYINPUT16), .Z(n1272) );
INV_X1 U960 ( .A(n1062), .ZN(n1085) );
NAND2_X1 U961 ( .A1(G221), .A2(n1274), .ZN(n1062) );
INV_X1 U962 ( .A(n1081), .ZN(n1060) );
XOR2_X1 U963 ( .A(n1275), .B(G469), .Z(n1081) );
NAND2_X1 U964 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U965 ( .A(n1278), .B(n1279), .Z(n1276) );
XOR2_X1 U966 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U967 ( .A(n1185), .B(n1282), .ZN(n1281) );
NOR2_X1 U968 ( .A1(KEYINPUT15), .A2(n1283), .ZN(n1282) );
NAND2_X1 U969 ( .A1(G227), .A2(n1121), .ZN(n1185) );
XOR2_X1 U970 ( .A(KEYINPUT10), .B(G140), .Z(n1280) );
XOR2_X1 U971 ( .A(n1284), .B(n1285), .Z(n1278) );
INV_X1 U972 ( .A(n1177), .ZN(n1285) );
XNOR2_X1 U973 ( .A(KEYINPUT0), .B(n1286), .ZN(n1177) );
NOR2_X1 U974 ( .A1(KEYINPUT45), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U975 ( .A(n1288), .B(n1175), .ZN(n1284) );
INV_X1 U976 ( .A(n1043), .ZN(n1263) );
NAND2_X1 U977 ( .A1(n1050), .A2(n1289), .ZN(n1043) );
NAND4_X1 U978 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1136), .ZN(n1289) );
INV_X1 U979 ( .A(G898), .ZN(n1136) );
NAND3_X1 U980 ( .A1(n1256), .A2(n1121), .A3(G952), .ZN(n1050) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n1256) );
NAND2_X1 U982 ( .A1(n1290), .A2(n1094), .ZN(n1042) );
NAND2_X1 U983 ( .A1(G214), .A2(n1291), .ZN(n1094) );
INV_X1 U984 ( .A(n1066), .ZN(n1290) );
XNOR2_X1 U985 ( .A(n1093), .B(n1092), .ZN(n1066) );
NAND2_X1 U986 ( .A1(G210), .A2(n1291), .ZN(n1092) );
NAND2_X1 U987 ( .A1(n1292), .A2(n1277), .ZN(n1291) );
INV_X1 U988 ( .A(G237), .ZN(n1292) );
NAND4_X1 U989 ( .A1(n1293), .A2(n1277), .A3(n1294), .A4(n1295), .ZN(n1093) );
NAND2_X1 U990 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
INV_X1 U991 ( .A(KEYINPUT38), .ZN(n1297) );
NAND2_X1 U992 ( .A1(n1193), .A2(n1298), .ZN(n1296) );
XNOR2_X1 U993 ( .A(KEYINPUT61), .B(n1299), .ZN(n1298) );
NAND2_X1 U994 ( .A1(KEYINPUT38), .A2(n1300), .ZN(n1294) );
NAND2_X1 U995 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND3_X1 U996 ( .A1(KEYINPUT61), .A2(n1193), .A3(n1299), .ZN(n1302) );
OR2_X1 U997 ( .A1(n1299), .A2(KEYINPUT61), .ZN(n1301) );
OR2_X1 U998 ( .A1(n1299), .A2(n1193), .ZN(n1293) );
XNOR2_X1 U999 ( .A(n1130), .B(n1132), .ZN(n1193) );
XNOR2_X1 U1000 ( .A(n1303), .B(n1304), .ZN(n1132) );
NOR2_X1 U1001 ( .A1(KEYINPUT53), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1002 ( .A(n1306), .B(n1288), .Z(n1130) );
XOR2_X1 U1003 ( .A(n1254), .B(n1273), .Z(n1288) );
XOR2_X1 U1004 ( .A(G122), .B(n1287), .Z(n1306) );
XNOR2_X1 U1005 ( .A(G104), .B(G107), .ZN(n1287) );
XNOR2_X1 U1006 ( .A(n1198), .B(n1113), .ZN(n1299) );
XOR2_X1 U1007 ( .A(G125), .B(n1175), .Z(n1113) );
NOR2_X1 U1008 ( .A1(n1135), .A2(G953), .ZN(n1198) );
INV_X1 U1009 ( .A(G224), .ZN(n1135) );
INV_X1 U1010 ( .A(n1053), .ZN(n1082) );
NAND2_X1 U1011 ( .A1(n1240), .A2(n1264), .ZN(n1053) );
XOR2_X1 U1012 ( .A(n1307), .B(G475), .Z(n1264) );
NAND2_X1 U1013 ( .A1(n1156), .A2(n1277), .ZN(n1307) );
XNOR2_X1 U1014 ( .A(n1308), .B(n1309), .ZN(n1156) );
XOR2_X1 U1015 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1016 ( .A(n1312), .B(n1313), .Z(n1311) );
AND2_X1 U1017 ( .A1(n1314), .A2(G214), .ZN(n1313) );
NOR2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1315), .ZN(n1312) );
XOR2_X1 U1019 ( .A(G104), .B(n1316), .Z(n1315) );
NOR2_X1 U1020 ( .A1(KEYINPUT17), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1021 ( .A(G113), .B(G122), .ZN(n1317) );
NOR2_X1 U1022 ( .A1(G143), .A2(KEYINPUT23), .ZN(n1310) );
XOR2_X1 U1023 ( .A(n1318), .B(n1319), .Z(n1308) );
XOR2_X1 U1024 ( .A(G146), .B(G140), .Z(n1319) );
XOR2_X1 U1025 ( .A(n1118), .B(G125), .Z(n1318) );
XOR2_X1 U1026 ( .A(n1320), .B(n1321), .Z(n1240) );
XOR2_X1 U1027 ( .A(KEYINPUT6), .B(G478), .Z(n1321) );
OR2_X1 U1028 ( .A1(n1151), .A2(G902), .ZN(n1320) );
XNOR2_X1 U1029 ( .A(n1322), .B(n1323), .ZN(n1151) );
XOR2_X1 U1030 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1031 ( .A(G122), .B(G116), .Z(n1325) );
XOR2_X1 U1032 ( .A(KEYINPUT24), .B(G143), .Z(n1324) );
XOR2_X1 U1033 ( .A(n1326), .B(n1327), .Z(n1322) );
XOR2_X1 U1034 ( .A(G107), .B(n1328), .Z(n1327) );
NOR2_X1 U1035 ( .A1(KEYINPUT44), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1036 ( .A(KEYINPUT59), .B(G134), .Z(n1329) );
XOR2_X1 U1037 ( .A(n1330), .B(n1331), .Z(n1326) );
NOR2_X1 U1038 ( .A1(G128), .A2(KEYINPUT3), .ZN(n1331) );
NAND3_X1 U1039 ( .A1(G217), .A2(n1121), .A3(G234), .ZN(n1330) );
INV_X1 U1040 ( .A(n1231), .ZN(n1078) );
NAND2_X1 U1041 ( .A1(n1267), .A2(n1265), .ZN(n1231) );
INV_X1 U1042 ( .A(n1268), .ZN(n1265) );
XNOR2_X1 U1043 ( .A(G472), .B(n1332), .ZN(n1268) );
NOR2_X1 U1044 ( .A1(n1095), .A2(KEYINPUT43), .ZN(n1332) );
AND2_X1 U1045 ( .A1(n1333), .A2(n1277), .ZN(n1095) );
XOR2_X1 U1046 ( .A(n1334), .B(n1335), .Z(n1333) );
NAND2_X1 U1047 ( .A1(KEYINPUT48), .A2(n1162), .ZN(n1335) );
AND2_X1 U1048 ( .A1(n1336), .A2(n1337), .ZN(n1162) );
NAND2_X1 U1049 ( .A1(n1338), .A2(n1254), .ZN(n1337) );
INV_X1 U1050 ( .A(G101), .ZN(n1254) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1314), .ZN(n1338) );
NAND3_X1 U1052 ( .A1(G210), .A2(n1314), .A3(G101), .ZN(n1336) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1314) );
NAND2_X1 U1054 ( .A1(n1339), .A2(n1340), .ZN(n1334) );
NAND2_X1 U1055 ( .A1(n1341), .A2(n1167), .ZN(n1340) );
XOR2_X1 U1056 ( .A(KEYINPUT19), .B(n1342), .Z(n1339) );
NOR2_X1 U1057 ( .A1(n1167), .A2(n1341), .ZN(n1342) );
XNOR2_X1 U1058 ( .A(n1175), .B(n1343), .ZN(n1341) );
NOR2_X1 U1059 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NOR2_X1 U1060 ( .A1(KEYINPUT5), .A2(n1283), .ZN(n1345) );
INV_X1 U1061 ( .A(n1174), .ZN(n1283) );
NOR2_X1 U1062 ( .A1(KEYINPUT4), .A2(n1174), .ZN(n1344) );
XOR2_X1 U1063 ( .A(n1118), .B(n1346), .Z(n1174) );
XOR2_X1 U1064 ( .A(G137), .B(G134), .Z(n1346) );
INV_X1 U1065 ( .A(G131), .ZN(n1118) );
XNOR2_X1 U1066 ( .A(n1347), .B(n1348), .ZN(n1175) );
XOR2_X1 U1067 ( .A(KEYINPUT21), .B(G146), .Z(n1348) );
XOR2_X1 U1068 ( .A(n1253), .B(G143), .Z(n1347) );
XOR2_X1 U1069 ( .A(n1305), .B(n1349), .Z(n1167) );
XOR2_X1 U1070 ( .A(KEYINPUT20), .B(n1303), .Z(n1349) );
XOR2_X1 U1071 ( .A(G113), .B(G119), .Z(n1303) );
XOR2_X1 U1072 ( .A(G116), .B(KEYINPUT41), .Z(n1305) );
XOR2_X1 U1073 ( .A(n1088), .B(n1350), .Z(n1267) );
NOR2_X1 U1074 ( .A1(n1090), .A2(KEYINPUT33), .ZN(n1350) );
NOR2_X1 U1075 ( .A1(n1143), .A2(G902), .ZN(n1090) );
INV_X1 U1076 ( .A(n1141), .ZN(n1143) );
NAND2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1141) );
NAND2_X1 U1078 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1079 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
INV_X1 U1080 ( .A(n1357), .ZN(n1353) );
XOR2_X1 U1081 ( .A(KEYINPUT7), .B(n1358), .Z(n1351) );
AND3_X1 U1082 ( .A1(n1357), .A2(n1356), .A3(n1355), .ZN(n1358) );
NAND2_X1 U1083 ( .A1(n1359), .A2(n1360), .ZN(n1355) );
NAND2_X1 U1084 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XNOR2_X1 U1085 ( .A(G146), .B(n1363), .ZN(n1359) );
NAND3_X1 U1086 ( .A1(n1364), .A2(n1362), .A3(n1361), .ZN(n1356) );
XOR2_X1 U1087 ( .A(n1365), .B(KEYINPUT63), .Z(n1361) );
NAND2_X1 U1088 ( .A1(n1366), .A2(n1273), .ZN(n1365) );
XOR2_X1 U1089 ( .A(G119), .B(n1253), .Z(n1366) );
INV_X1 U1090 ( .A(G128), .ZN(n1253) );
NAND2_X1 U1091 ( .A1(G110), .A2(n1367), .ZN(n1362) );
XOR2_X1 U1092 ( .A(G128), .B(G119), .Z(n1367) );
XOR2_X1 U1093 ( .A(n1363), .B(G146), .Z(n1364) );
NAND2_X1 U1094 ( .A1(n1368), .A2(n1369), .ZN(n1363) );
NAND2_X1 U1095 ( .A1(G140), .A2(G125), .ZN(n1369) );
NAND2_X1 U1096 ( .A1(n1370), .A2(n1241), .ZN(n1368) );
INV_X1 U1097 ( .A(G140), .ZN(n1241) );
XNOR2_X1 U1098 ( .A(G125), .B(KEYINPUT27), .ZN(n1370) );
NAND2_X1 U1099 ( .A1(n1371), .A2(n1372), .ZN(n1357) );
NAND2_X1 U1100 ( .A1(n1373), .A2(n1119), .ZN(n1372) );
INV_X1 U1101 ( .A(G137), .ZN(n1119) );
NAND2_X1 U1102 ( .A1(n1374), .A2(G137), .ZN(n1371) );
XOR2_X1 U1103 ( .A(KEYINPUT30), .B(n1373), .Z(n1374) );
AND3_X1 U1104 ( .A1(G234), .A2(n1121), .A3(G221), .ZN(n1373) );
INV_X1 U1105 ( .A(G953), .ZN(n1121) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1274), .ZN(n1088) );
NAND2_X1 U1107 ( .A1(G234), .A2(n1277), .ZN(n1274) );
INV_X1 U1108 ( .A(G902), .ZN(n1277) );
INV_X1 U1109 ( .A(G110), .ZN(n1273) );
endmodule


