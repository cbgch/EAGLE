//Key = 0010001010110100100010000110101100001011001111001100110011111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320;

XNOR2_X1 U719 ( .A(n994), .B(n995), .ZN(G9) );
XOR2_X1 U720 ( .A(KEYINPUT31), .B(G107), .Z(n995) );
NOR2_X1 U721 ( .A1(n996), .A2(n997), .ZN(G75) );
NOR4_X1 U722 ( .A1(G953), .A2(n998), .A3(n999), .A4(n1000), .ZN(n997) );
NOR2_X1 U723 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U725 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U727 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR2_X1 U728 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U730 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U731 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1011) );
NOR2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR3_X1 U734 ( .A1(n1020), .A2(n1023), .A3(n1014), .ZN(n1007) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR4_X1 U737 ( .A1(n1028), .A2(n1014), .A3(n1020), .A4(n1010), .ZN(n1003) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR3_X1 U739 ( .A1(n998), .A2(G953), .A3(G952), .ZN(n996) );
AND4_X1 U740 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n998) );
NOR4_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
NAND3_X1 U742 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1035) );
NOR3_X1 U743 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1033) );
XNOR2_X1 U744 ( .A(n1045), .B(KEYINPUT36), .ZN(n1044) );
XOR2_X1 U745 ( .A(n1046), .B(KEYINPUT39), .Z(n1042) );
XOR2_X1 U746 ( .A(n1047), .B(n1048), .Z(G72) );
XOR2_X1 U747 ( .A(n1049), .B(n1050), .Z(n1048) );
NOR2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U749 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U750 ( .A(n1055), .B(n1056), .Z(n1054) );
XNOR2_X1 U751 ( .A(n1057), .B(n1058), .ZN(n1053) );
NAND2_X1 U752 ( .A1(n1059), .A2(KEYINPUT42), .ZN(n1057) );
XNOR2_X1 U753 ( .A(G131), .B(n1060), .ZN(n1059) );
NOR2_X1 U754 ( .A1(KEYINPUT5), .A2(n1061), .ZN(n1060) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1049) );
NAND2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U757 ( .A1(G953), .A2(n1066), .ZN(n1047) );
NAND2_X1 U758 ( .A1(G900), .A2(G227), .ZN(n1066) );
XOR2_X1 U759 ( .A(n1067), .B(n1068), .Z(G69) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1063), .ZN(n1069) );
AND2_X1 U762 ( .A1(G224), .A2(G898), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1067) );
NAND2_X1 U764 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U765 ( .A(n1075), .B(n1076), .ZN(n1072) );
NOR2_X1 U766 ( .A1(KEYINPUT24), .A2(n1077), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XNOR2_X1 U768 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1084), .ZN(G63) );
XOR2_X1 U771 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U772 ( .A1(KEYINPUT27), .A2(n1087), .ZN(n1086) );
NAND2_X1 U773 ( .A1(n1088), .A2(G478), .ZN(n1085) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1089), .ZN(G60) );
XOR2_X1 U775 ( .A(n1090), .B(n1091), .Z(n1089) );
AND2_X1 U776 ( .A1(G475), .A2(n1088), .ZN(n1090) );
XNOR2_X1 U777 ( .A(G104), .B(n1092), .ZN(G6) );
NOR3_X1 U778 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(G57) );
AND2_X1 U779 ( .A1(KEYINPUT58), .A2(n1078), .ZN(n1095) );
NOR3_X1 U780 ( .A1(KEYINPUT58), .A2(n1096), .A3(n1063), .ZN(n1094) );
XOR2_X1 U781 ( .A(n1097), .B(n1098), .Z(n1093) );
XOR2_X1 U782 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U783 ( .A(KEYINPUT20), .B(n1101), .Z(n1100) );
NOR3_X1 U784 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1000), .B(KEYINPUT43), .Z(n1103) );
XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n1105), .ZN(n1102) );
XOR2_X1 U787 ( .A(n1106), .B(n1107), .Z(n1097) );
NOR2_X1 U788 ( .A1(KEYINPUT47), .A2(n1108), .ZN(n1107) );
NAND2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
XOR2_X1 U790 ( .A(KEYINPUT57), .B(n1111), .Z(n1109) );
NOR2_X1 U791 ( .A1(n1078), .A2(n1112), .ZN(G54) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U793 ( .A(n1115), .B(n1116), .Z(n1114) );
AND2_X1 U794 ( .A1(G469), .A2(n1088), .ZN(n1115) );
INV_X1 U795 ( .A(n1083), .ZN(n1088) );
XNOR2_X1 U796 ( .A(G110), .B(n1117), .ZN(n1113) );
XNOR2_X1 U797 ( .A(KEYINPUT11), .B(n1118), .ZN(n1117) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1063), .ZN(n1078) );
NOR2_X1 U799 ( .A1(n1120), .A2(n1121), .ZN(G51) );
XOR2_X1 U800 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1122) );
NOR2_X1 U802 ( .A1(n1126), .A2(n1083), .ZN(n1125) );
NAND2_X1 U803 ( .A1(n1127), .A2(n1000), .ZN(n1083) );
NAND3_X1 U804 ( .A1(n1128), .A2(n1129), .A3(n1064), .ZN(n1000) );
AND4_X1 U805 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1064) );
NOR4_X1 U806 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
NOR2_X1 U807 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR3_X1 U809 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
NOR2_X1 U810 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
AND3_X1 U811 ( .A1(KEYINPUT23), .A2(n1020), .A3(n1021), .ZN(n1145) );
NOR2_X1 U812 ( .A1(n1025), .A2(n1147), .ZN(n1143) );
NOR3_X1 U813 ( .A1(n1148), .A2(KEYINPUT30), .A3(n1149), .ZN(n1147) );
INV_X1 U814 ( .A(n1146), .ZN(n1025) );
NOR4_X1 U815 ( .A1(n1150), .A2(n1149), .A3(n1010), .A4(n1151), .ZN(n1140) );
INV_X1 U816 ( .A(n1152), .ZN(n1010) );
XNOR2_X1 U817 ( .A(n1030), .B(KEYINPUT46), .ZN(n1150) );
NAND2_X1 U818 ( .A1(KEYINPUT30), .A2(n1153), .ZN(n1132) );
INV_X1 U819 ( .A(n1154), .ZN(n1153) );
NAND2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1131) );
OR2_X1 U821 ( .A1(n1157), .A2(KEYINPUT23), .ZN(n1130) );
XNOR2_X1 U822 ( .A(KEYINPUT26), .B(n1065), .ZN(n1129) );
INV_X1 U823 ( .A(n1070), .ZN(n1128) );
NAND4_X1 U824 ( .A1(n1158), .A2(n1092), .A3(n1159), .A4(n1160), .ZN(n1070) );
NOR4_X1 U825 ( .A1(n994), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1160) );
AND2_X1 U826 ( .A1(n1029), .A2(n1164), .ZN(n994) );
NAND4_X1 U827 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1159) );
NAND2_X1 U828 ( .A1(n1169), .A2(n1006), .ZN(n1168) );
NAND2_X1 U829 ( .A1(KEYINPUT19), .A2(n1021), .ZN(n1169) );
NAND3_X1 U830 ( .A1(n1170), .A2(n1151), .A3(n1171), .ZN(n1167) );
OR2_X1 U831 ( .A1(n1172), .A2(KEYINPUT19), .ZN(n1170) );
NAND2_X1 U832 ( .A1(n1030), .A2(n1164), .ZN(n1092) );
NOR3_X1 U833 ( .A1(n1014), .A2(n1173), .A3(n1174), .ZN(n1164) );
INV_X1 U834 ( .A(n1175), .ZN(n1014) );
NAND4_X1 U835 ( .A1(n1176), .A2(n1177), .A3(n1175), .A4(n1178), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1046), .A2(n1031), .ZN(n1178) );
OR2_X1 U837 ( .A1(n1179), .A2(KEYINPUT29), .ZN(n1177) );
NAND2_X1 U838 ( .A1(KEYINPUT29), .A2(n1180), .ZN(n1176) );
NAND3_X1 U839 ( .A1(n1166), .A2(n1149), .A3(n1152), .ZN(n1180) );
XNOR2_X1 U840 ( .A(KEYINPUT61), .B(G902), .ZN(n1127) );
NAND3_X1 U841 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1124) );
NAND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
OR3_X1 U843 ( .A1(n1185), .A2(n1184), .A3(KEYINPUT14), .ZN(n1182) );
AND2_X1 U844 ( .A1(KEYINPUT63), .A2(n1186), .ZN(n1184) );
NAND2_X1 U845 ( .A1(KEYINPUT14), .A2(n1187), .ZN(n1181) );
OR2_X1 U846 ( .A1(n1185), .A2(n1186), .ZN(n1187) );
NOR2_X1 U847 ( .A1(n1119), .A2(n1188), .ZN(n1120) );
XNOR2_X1 U848 ( .A(KEYINPUT16), .B(n1063), .ZN(n1188) );
INV_X1 U849 ( .A(n1096), .ZN(n1119) );
XNOR2_X1 U850 ( .A(G952), .B(KEYINPUT33), .ZN(n1096) );
XOR2_X1 U851 ( .A(G146), .B(n1136), .Z(G48) );
AND2_X1 U852 ( .A1(n1189), .A2(n1030), .ZN(n1136) );
XNOR2_X1 U853 ( .A(n1190), .B(n1135), .ZN(G45) );
NOR4_X1 U854 ( .A1(n1046), .A2(n1138), .A3(n1031), .A4(n1191), .ZN(n1135) );
NAND2_X1 U855 ( .A1(n1165), .A2(n1021), .ZN(n1191) );
XNOR2_X1 U856 ( .A(G140), .B(n1065), .ZN(G42) );
NAND3_X1 U857 ( .A1(n1030), .A2(n1192), .A3(n1022), .ZN(n1065) );
XOR2_X1 U858 ( .A(n1193), .B(n1194), .Z(G39) );
XNOR2_X1 U859 ( .A(G137), .B(KEYINPUT1), .ZN(n1194) );
NAND2_X1 U860 ( .A1(n1195), .A2(n1156), .ZN(n1193) );
XNOR2_X1 U861 ( .A(n1155), .B(KEYINPUT13), .ZN(n1195) );
NOR4_X1 U862 ( .A1(n1006), .A2(n1148), .A3(n1146), .A4(n1138), .ZN(n1155) );
XNOR2_X1 U863 ( .A(G134), .B(n1157), .ZN(G36) );
NAND3_X1 U864 ( .A1(n1192), .A2(n1029), .A3(n1021), .ZN(n1157) );
XOR2_X1 U865 ( .A(G131), .B(n1134), .Z(G33) );
AND3_X1 U866 ( .A1(n1030), .A2(n1192), .A3(n1021), .ZN(n1134) );
NOR3_X1 U867 ( .A1(n1146), .A2(n1138), .A3(n1020), .ZN(n1192) );
INV_X1 U868 ( .A(n1156), .ZN(n1020) );
NOR2_X1 U869 ( .A1(n1017), .A2(n1036), .ZN(n1156) );
INV_X1 U870 ( .A(n1018), .ZN(n1036) );
XNOR2_X1 U871 ( .A(G128), .B(n1154), .ZN(G30) );
NAND2_X1 U872 ( .A1(n1189), .A2(n1029), .ZN(n1154) );
INV_X1 U873 ( .A(n1142), .ZN(n1029) );
NOR3_X1 U874 ( .A1(n1174), .A2(n1138), .A3(n1148), .ZN(n1189) );
XNOR2_X1 U875 ( .A(G101), .B(n1196), .ZN(G3) );
NAND4_X1 U876 ( .A1(KEYINPUT49), .A2(n1171), .A3(n1197), .A4(n1021), .ZN(n1196) );
NOR2_X1 U877 ( .A1(n1173), .A2(n1174), .ZN(n1197) );
INV_X1 U878 ( .A(n1165), .ZN(n1174) );
INV_X1 U879 ( .A(n1166), .ZN(n1173) );
XNOR2_X1 U880 ( .A(G125), .B(n1198), .ZN(G27) );
NAND4_X1 U881 ( .A1(n1152), .A2(n1030), .A3(n1022), .A4(n1199), .ZN(n1198) );
NOR3_X1 U882 ( .A1(n1149), .A2(KEYINPUT22), .A3(n1138), .ZN(n1199) );
AND2_X1 U883 ( .A1(n1002), .A2(n1200), .ZN(n1138) );
NAND3_X1 U884 ( .A1(G902), .A2(n1201), .A3(n1051), .ZN(n1200) );
NOR2_X1 U885 ( .A1(n1063), .A2(G900), .ZN(n1051) );
XNOR2_X1 U886 ( .A(G122), .B(n1202), .ZN(G24) );
NAND3_X1 U887 ( .A1(n1179), .A2(n1175), .A3(n1203), .ZN(n1202) );
NOR3_X1 U888 ( .A1(n1031), .A2(KEYINPUT41), .A3(n1046), .ZN(n1203) );
NOR2_X1 U889 ( .A1(n1204), .A2(n1205), .ZN(n1175) );
XOR2_X1 U890 ( .A(G119), .B(n1163), .Z(G21) );
NOR3_X1 U891 ( .A1(n1006), .A2(n1148), .A3(n1206), .ZN(n1163) );
NAND2_X1 U892 ( .A1(n1205), .A2(n1204), .ZN(n1148) );
XNOR2_X1 U893 ( .A(n1162), .B(n1207), .ZN(G18) );
NOR2_X1 U894 ( .A1(G116), .A2(KEYINPUT40), .ZN(n1207) );
NOR3_X1 U895 ( .A1(n1172), .A2(n1142), .A3(n1206), .ZN(n1162) );
NAND2_X1 U896 ( .A1(n1046), .A2(n1208), .ZN(n1142) );
INV_X1 U897 ( .A(n1021), .ZN(n1172) );
XNOR2_X1 U898 ( .A(n1209), .B(n1161), .ZN(G15) );
AND3_X1 U899 ( .A1(n1021), .A2(n1030), .A3(n1179), .ZN(n1161) );
INV_X1 U900 ( .A(n1206), .ZN(n1179) );
NAND3_X1 U901 ( .A1(n1016), .A2(n1166), .A3(n1152), .ZN(n1206) );
NOR2_X1 U902 ( .A1(n1026), .A2(n1037), .ZN(n1152) );
INV_X1 U903 ( .A(n1027), .ZN(n1037) );
INV_X1 U904 ( .A(n1149), .ZN(n1016) );
NOR2_X1 U905 ( .A1(n1208), .A2(n1046), .ZN(n1030) );
NOR2_X1 U906 ( .A1(n1204), .A2(n1032), .ZN(n1021) );
XNOR2_X1 U907 ( .A(G110), .B(n1210), .ZN(G12) );
NAND4_X1 U908 ( .A1(n1171), .A2(n1022), .A3(n1165), .A4(n1211), .ZN(n1210) );
XNOR2_X1 U909 ( .A(KEYINPUT45), .B(n1166), .ZN(n1211) );
NAND2_X1 U910 ( .A1(n1002), .A2(n1212), .ZN(n1166) );
NAND4_X1 U911 ( .A1(n1213), .A2(G953), .A3(G902), .A4(n1074), .ZN(n1212) );
INV_X1 U912 ( .A(G898), .ZN(n1074) );
XOR2_X1 U913 ( .A(n1201), .B(KEYINPUT4), .Z(n1213) );
NAND3_X1 U914 ( .A1(n1201), .A2(n1063), .A3(G952), .ZN(n1002) );
NAND2_X1 U915 ( .A1(G237), .A2(G234), .ZN(n1201) );
NOR2_X1 U916 ( .A1(n1149), .A2(n1146), .ZN(n1165) );
NAND2_X1 U917 ( .A1(n1027), .A2(n1026), .ZN(n1146) );
NAND3_X1 U918 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1026) );
INV_X1 U919 ( .A(n1038), .ZN(n1216) );
NOR2_X1 U920 ( .A1(n1217), .A2(G469), .ZN(n1038) );
OR2_X1 U921 ( .A1(G469), .A2(KEYINPUT53), .ZN(n1215) );
NAND2_X1 U922 ( .A1(n1045), .A2(KEYINPUT53), .ZN(n1214) );
AND2_X1 U923 ( .A1(G469), .A2(n1217), .ZN(n1045) );
NAND2_X1 U924 ( .A1(n1218), .A2(n1105), .ZN(n1217) );
XNOR2_X1 U925 ( .A(n1219), .B(n1116), .ZN(n1218) );
XNOR2_X1 U926 ( .A(n1220), .B(n1221), .ZN(n1116) );
XOR2_X1 U927 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U928 ( .A(n1224), .B(n1225), .Z(n1223) );
NOR2_X1 U929 ( .A1(KEYINPUT15), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U930 ( .A(KEYINPUT7), .B(n1227), .ZN(n1226) );
INV_X1 U931 ( .A(G104), .ZN(n1227) );
NAND2_X1 U932 ( .A1(G227), .A2(n1063), .ZN(n1224) );
XNOR2_X1 U933 ( .A(G101), .B(G107), .ZN(n1222) );
XOR2_X1 U934 ( .A(n1228), .B(n1056), .Z(n1220) );
XNOR2_X1 U935 ( .A(n1229), .B(KEYINPUT44), .ZN(n1056) );
XOR2_X1 U936 ( .A(n1230), .B(n1061), .Z(n1228) );
NAND3_X1 U937 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1219) );
NAND2_X1 U938 ( .A1(n1234), .A2(n1118), .ZN(n1233) );
NAND2_X1 U939 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U940 ( .A(KEYINPUT59), .B(n1237), .ZN(n1235) );
NAND3_X1 U941 ( .A1(G140), .A2(n1237), .A3(n1236), .ZN(n1232) );
INV_X1 U942 ( .A(KEYINPUT55), .ZN(n1236) );
INV_X1 U943 ( .A(G110), .ZN(n1237) );
NAND2_X1 U944 ( .A1(KEYINPUT55), .A2(G110), .ZN(n1231) );
NAND2_X1 U945 ( .A1(G221), .A2(n1238), .ZN(n1027) );
NAND2_X1 U946 ( .A1(n1018), .A2(n1017), .ZN(n1149) );
NAND2_X1 U947 ( .A1(n1239), .A2(n1040), .ZN(n1017) );
NAND2_X1 U948 ( .A1(n1240), .A2(n1126), .ZN(n1040) );
XOR2_X1 U949 ( .A(KEYINPUT2), .B(n1043), .Z(n1239) );
NOR2_X1 U950 ( .A1(n1126), .A2(n1240), .ZN(n1043) );
AND2_X1 U951 ( .A1(n1241), .A2(n1105), .ZN(n1240) );
XOR2_X1 U952 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U953 ( .A(n1185), .B(n1123), .ZN(n1243) );
XOR2_X1 U954 ( .A(n1077), .B(n1075), .Z(n1123) );
XNOR2_X1 U955 ( .A(n1244), .B(KEYINPUT54), .ZN(n1075) );
NAND2_X1 U956 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U957 ( .A1(G110), .A2(n1247), .ZN(n1246) );
XOR2_X1 U958 ( .A(KEYINPUT25), .B(n1248), .Z(n1245) );
NOR2_X1 U959 ( .A1(G110), .A2(n1247), .ZN(n1248) );
XNOR2_X1 U960 ( .A(n1249), .B(n1250), .ZN(n1077) );
XOR2_X1 U961 ( .A(G101), .B(n1251), .Z(n1250) );
NOR2_X1 U962 ( .A1(KEYINPUT34), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U963 ( .A(G104), .B(n1253), .ZN(n1252) );
NOR2_X1 U964 ( .A1(KEYINPUT37), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U965 ( .A(G107), .B(KEYINPUT48), .ZN(n1254) );
XOR2_X1 U966 ( .A(n1255), .B(n1256), .Z(n1249) );
NAND2_X1 U967 ( .A1(KEYINPUT8), .A2(n1209), .ZN(n1255) );
INV_X1 U968 ( .A(G113), .ZN(n1209) );
XNOR2_X1 U969 ( .A(G125), .B(n1257), .ZN(n1185) );
NAND2_X1 U970 ( .A1(n1258), .A2(n1259), .ZN(n1242) );
NAND2_X1 U971 ( .A1(KEYINPUT38), .A2(n1260), .ZN(n1259) );
NAND2_X1 U972 ( .A1(KEYINPUT21), .A2(n1186), .ZN(n1258) );
INV_X1 U973 ( .A(n1260), .ZN(n1186) );
NAND2_X1 U974 ( .A1(G224), .A2(n1063), .ZN(n1260) );
NAND2_X1 U975 ( .A1(G210), .A2(n1261), .ZN(n1126) );
NAND2_X1 U976 ( .A1(G214), .A2(n1261), .ZN(n1018) );
NAND2_X1 U977 ( .A1(n1262), .A2(n1105), .ZN(n1261) );
INV_X1 U978 ( .A(G237), .ZN(n1262) );
INV_X1 U979 ( .A(n1151), .ZN(n1022) );
NAND2_X1 U980 ( .A1(n1032), .A2(n1204), .ZN(n1151) );
NAND3_X1 U981 ( .A1(n1263), .A2(n1264), .A3(n1041), .ZN(n1204) );
NAND3_X1 U982 ( .A1(n1082), .A2(n1105), .A3(n1080), .ZN(n1041) );
OR2_X1 U983 ( .A1(n1039), .A2(KEYINPUT32), .ZN(n1264) );
OR2_X1 U984 ( .A1(n1082), .A2(n1265), .ZN(n1039) );
AND2_X1 U985 ( .A1(n1105), .A2(n1080), .ZN(n1265) );
NAND3_X1 U986 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1080) );
OR2_X1 U987 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U988 ( .A1(KEYINPUT0), .A2(n1271), .ZN(n1267) );
NAND2_X1 U989 ( .A1(n1270), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U990 ( .A(KEYINPUT6), .B(n1269), .ZN(n1272) );
NAND2_X1 U991 ( .A1(n1273), .A2(n1274), .ZN(n1266) );
INV_X1 U992 ( .A(KEYINPUT0), .ZN(n1274) );
NAND2_X1 U993 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND3_X1 U994 ( .A1(KEYINPUT6), .A2(n1270), .A3(n1269), .ZN(n1276) );
XOR2_X1 U995 ( .A(n1277), .B(n1278), .Z(n1270) );
XOR2_X1 U996 ( .A(n1279), .B(n1055), .Z(n1278) );
NOR2_X1 U997 ( .A1(G146), .A2(KEYINPUT62), .ZN(n1279) );
XOR2_X1 U998 ( .A(n1280), .B(n1281), .Z(n1277) );
NOR2_X1 U999 ( .A1(KEYINPUT18), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U1000 ( .A(G119), .B(G128), .ZN(n1282) );
XNOR2_X1 U1001 ( .A(G110), .B(KEYINPUT12), .ZN(n1280) );
OR2_X1 U1002 ( .A1(n1269), .A2(KEYINPUT6), .ZN(n1275) );
XOR2_X1 U1003 ( .A(n1283), .B(G137), .Z(n1269) );
NAND2_X1 U1004 ( .A1(G221), .A2(n1284), .ZN(n1283) );
NAND2_X1 U1005 ( .A1(KEYINPUT32), .A2(n1082), .ZN(n1263) );
NAND2_X1 U1006 ( .A1(G217), .A2(n1238), .ZN(n1082) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1105), .ZN(n1238) );
INV_X1 U1008 ( .A(n1205), .ZN(n1032) );
XOR2_X1 U1009 ( .A(n1285), .B(n1104), .Z(n1205) );
INV_X1 U1010 ( .A(G472), .ZN(n1104) );
NAND2_X1 U1011 ( .A1(n1286), .A2(n1105), .ZN(n1285) );
INV_X1 U1012 ( .A(G902), .ZN(n1105) );
XOR2_X1 U1013 ( .A(n1287), .B(n1101), .Z(n1286) );
AND2_X1 U1014 ( .A1(n1288), .A2(n1289), .ZN(n1101) );
NAND2_X1 U1015 ( .A1(G113), .A2(n1256), .ZN(n1289) );
XOR2_X1 U1016 ( .A(n1290), .B(KEYINPUT35), .Z(n1288) );
OR2_X1 U1017 ( .A1(n1256), .A2(G113), .ZN(n1290) );
XOR2_X1 U1018 ( .A(G116), .B(G119), .Z(n1256) );
XOR2_X1 U1019 ( .A(n1291), .B(n1292), .Z(n1287) );
NOR2_X1 U1020 ( .A1(KEYINPUT3), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1021 ( .A(n1108), .B(KEYINPUT10), .ZN(n1293) );
XNOR2_X1 U1022 ( .A(n1294), .B(G101), .ZN(n1108) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1024 ( .A1(n1296), .A2(n1110), .ZN(n1291) );
NAND2_X1 U1025 ( .A1(n1297), .A2(n1257), .ZN(n1110) );
XOR2_X1 U1026 ( .A(KEYINPUT28), .B(n1111), .Z(n1296) );
NOR2_X1 U1027 ( .A1(n1297), .A2(n1257), .ZN(n1111) );
XOR2_X1 U1028 ( .A(n1229), .B(n1298), .Z(n1257) );
NOR3_X1 U1029 ( .A1(KEYINPUT9), .A2(n1299), .A3(n1300), .ZN(n1298) );
AND2_X1 U1030 ( .A1(n1301), .A2(n1058), .ZN(n1300) );
NOR2_X1 U1031 ( .A1(n1302), .A2(n1301), .ZN(n1299) );
INV_X1 U1032 ( .A(KEYINPUT50), .ZN(n1301) );
NOR2_X1 U1033 ( .A1(G146), .A2(n1190), .ZN(n1302) );
INV_X1 U1034 ( .A(G128), .ZN(n1229) );
XNOR2_X1 U1035 ( .A(n1061), .B(G131), .ZN(n1297) );
XOR2_X1 U1036 ( .A(G137), .B(n1303), .Z(n1061) );
INV_X1 U1037 ( .A(n1006), .ZN(n1171) );
NAND2_X1 U1038 ( .A1(n1031), .A2(n1046), .ZN(n1006) );
XOR2_X1 U1039 ( .A(n1304), .B(n1305), .Z(n1046) );
XOR2_X1 U1040 ( .A(KEYINPUT17), .B(G475), .Z(n1305) );
OR2_X1 U1041 ( .A1(n1091), .A2(G902), .ZN(n1304) );
XNOR2_X1 U1042 ( .A(n1306), .B(n1307), .ZN(n1091) );
XOR2_X1 U1043 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1295), .ZN(n1309) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1295) );
NAND2_X1 U1046 ( .A1(n1310), .A2(KEYINPUT56), .ZN(n1308) );
XNOR2_X1 U1047 ( .A(G104), .B(n1311), .ZN(n1310) );
XNOR2_X1 U1048 ( .A(n1247), .B(G113), .ZN(n1311) );
XOR2_X1 U1049 ( .A(n1230), .B(n1055), .Z(n1306) );
XNOR2_X1 U1050 ( .A(G125), .B(n1118), .ZN(n1055) );
INV_X1 U1051 ( .A(G140), .ZN(n1118) );
XNOR2_X1 U1052 ( .A(G131), .B(n1058), .ZN(n1230) );
XOR2_X1 U1053 ( .A(G143), .B(G146), .Z(n1058) );
INV_X1 U1054 ( .A(n1208), .ZN(n1031) );
XNOR2_X1 U1055 ( .A(n1312), .B(G478), .ZN(n1208) );
OR2_X1 U1056 ( .A1(n1087), .A2(G902), .ZN(n1312) );
XNOR2_X1 U1057 ( .A(n1313), .B(n1314), .ZN(n1087) );
XOR2_X1 U1058 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1059 ( .A(G116), .B(G107), .Z(n1316) );
XNOR2_X1 U1060 ( .A(KEYINPUT51), .B(n1247), .ZN(n1315) );
INV_X1 U1061 ( .A(G122), .ZN(n1247) );
XNOR2_X1 U1062 ( .A(n1303), .B(n1317), .ZN(n1313) );
XOR2_X1 U1063 ( .A(n1318), .B(n1319), .Z(n1317) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1284), .ZN(n1319) );
AND2_X1 U1065 ( .A1(G234), .A2(n1063), .ZN(n1284) );
INV_X1 U1066 ( .A(G953), .ZN(n1063) );
NAND2_X1 U1067 ( .A1(KEYINPUT60), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1068 ( .A(n1190), .B(G128), .ZN(n1320) );
INV_X1 U1069 ( .A(G143), .ZN(n1190) );
XOR2_X1 U1070 ( .A(G134), .B(KEYINPUT52), .Z(n1303) );
endmodule


