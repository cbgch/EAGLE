//Key = 1101101110011111000111111110111000101001011101111011111101011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351;

XOR2_X1 U738 ( .A(n1028), .B(n1029), .Z(G9) );
NAND2_X1 U739 ( .A1(KEYINPUT14), .A2(n1030), .ZN(n1028) );
INV_X1 U740 ( .A(G107), .ZN(n1030) );
NOR2_X1 U741 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR4_X1 U742 ( .A1(G953), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR3_X1 U745 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
AND2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR3_X1 U752 ( .A1(n1046), .A2(n1055), .A3(n1050), .ZN(n1038) );
NOR3_X1 U753 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NOR3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
XOR2_X1 U755 ( .A(KEYINPUT47), .B(n1062), .Z(n1059) );
NOR2_X1 U756 ( .A1(n1063), .A2(n1042), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U758 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U759 ( .A1(n1033), .A2(G953), .A3(G952), .ZN(n1031) );
AND4_X1 U760 ( .A1(n1060), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1033) );
NOR4_X1 U761 ( .A1(n1071), .A2(n1054), .A3(n1072), .A4(n1073), .ZN(n1070) );
AND2_X1 U762 ( .A1(n1074), .A2(G472), .ZN(n1073) );
NOR2_X1 U763 ( .A1(n1050), .A2(n1075), .ZN(n1069) );
XOR2_X1 U764 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U765 ( .A(n1078), .B(KEYINPUT62), .Z(n1077) );
XOR2_X1 U766 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1079) );
NAND3_X1 U770 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND2_X1 U771 ( .A1(G953), .A2(n1084), .ZN(n1088) );
XOR2_X1 U772 ( .A(n1090), .B(KEYINPUT12), .Z(n1087) );
NAND3_X1 U773 ( .A1(n1090), .A2(n1082), .A3(n1091), .ZN(n1085) );
INV_X1 U774 ( .A(n1089), .ZN(n1091) );
XOR2_X1 U775 ( .A(n1092), .B(n1093), .Z(n1089) );
XOR2_X1 U776 ( .A(KEYINPUT13), .B(n1094), .Z(n1093) );
NOR2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U778 ( .A(n1097), .B(KEYINPUT15), .Z(n1096) );
NAND2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U780 ( .A(G131), .B(KEYINPUT7), .ZN(n1098) );
NOR2_X1 U781 ( .A1(G131), .A2(n1099), .ZN(n1095) );
XOR2_X1 U782 ( .A(KEYINPUT56), .B(n1100), .Z(n1099) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1092) );
NAND2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1090) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(G69) );
NOR2_X1 U786 ( .A1(n1107), .A2(n1082), .ZN(n1106) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1107) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U790 ( .A(KEYINPUT58), .B(n1112), .Z(n1110) );
NOR2_X1 U791 ( .A1(G953), .A2(n1113), .ZN(n1112) );
NAND3_X1 U792 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1108) );
INV_X1 U793 ( .A(n1116), .ZN(n1114) );
XNOR2_X1 U794 ( .A(n1117), .B(n1118), .ZN(n1113) );
XNOR2_X1 U795 ( .A(n1119), .B(KEYINPUT9), .ZN(n1117) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XNOR2_X1 U797 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U799 ( .A1(n1120), .A2(n1126), .ZN(G63) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U801 ( .A1(n1129), .A2(n1125), .ZN(n1127) );
INV_X1 U802 ( .A(G478), .ZN(n1129) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1130), .ZN(G60) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1125), .ZN(n1131) );
INV_X1 U806 ( .A(G475), .ZN(n1133) );
XNOR2_X1 U807 ( .A(G104), .B(n1134), .ZN(G6) );
NAND2_X1 U808 ( .A1(n1135), .A2(n1065), .ZN(n1134) );
XOR2_X1 U809 ( .A(n1136), .B(KEYINPUT20), .Z(n1135) );
NOR2_X1 U810 ( .A1(n1120), .A2(n1137), .ZN(G57) );
XOR2_X1 U811 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U812 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U813 ( .A(n1142), .B(n1143), .ZN(n1141) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(n1138) );
XOR2_X1 U815 ( .A(KEYINPUT34), .B(KEYINPUT32), .Z(n1145) );
XOR2_X1 U816 ( .A(n1146), .B(n1147), .Z(n1144) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1125), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1120), .A2(n1149), .ZN(G54) );
XOR2_X1 U819 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U820 ( .A1(n1078), .A2(n1125), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1152), .A2(KEYINPUT22), .ZN(n1150) );
XOR2_X1 U822 ( .A(n1153), .B(KEYINPUT17), .Z(n1152) );
NOR2_X1 U823 ( .A1(n1120), .A2(n1154), .ZN(G51) );
XOR2_X1 U824 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U826 ( .A(n1159), .B(n1143), .ZN(n1158) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1125), .ZN(n1159) );
NAND2_X1 U828 ( .A1(G902), .A2(n1035), .ZN(n1125) );
NAND3_X1 U829 ( .A1(n1115), .A2(n1103), .A3(n1161), .ZN(n1035) );
XOR2_X1 U830 ( .A(n1104), .B(KEYINPUT44), .Z(n1161) );
AND4_X1 U831 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1103) );
NOR3_X1 U832 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
AND3_X1 U833 ( .A1(n1057), .A2(n1048), .A3(n1169), .ZN(n1168) );
NOR2_X1 U834 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1047), .A2(n1172), .ZN(n1170) );
XOR2_X1 U836 ( .A(KEYINPUT33), .B(n1048), .Z(n1172) );
INV_X1 U837 ( .A(n1111), .ZN(n1115) );
NAND4_X1 U838 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1111) );
NOR4_X1 U839 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR2_X1 U840 ( .A1(n1181), .A2(n1136), .ZN(n1180) );
NAND4_X1 U841 ( .A1(n1048), .A2(n1052), .A3(n1182), .A4(n1183), .ZN(n1136) );
NOR4_X1 U842 ( .A1(n1184), .A2(n1042), .A3(n1185), .A4(n1186), .ZN(n1179) );
NAND3_X1 U843 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1184) );
NAND2_X1 U844 ( .A1(KEYINPUT48), .A2(n1190), .ZN(n1188) );
NAND2_X1 U845 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
INV_X1 U846 ( .A(KEYINPUT48), .ZN(n1192) );
NAND2_X1 U847 ( .A1(n1183), .A2(n1181), .ZN(n1191) );
INV_X1 U848 ( .A(n1193), .ZN(n1178) );
NOR2_X1 U849 ( .A1(n1194), .A2(n1029), .ZN(n1175) );
AND4_X1 U850 ( .A1(n1052), .A2(n1182), .A3(n1195), .A4(n1047), .ZN(n1029) );
XOR2_X1 U851 ( .A(n1196), .B(n1197), .Z(n1155) );
XOR2_X1 U852 ( .A(KEYINPUT59), .B(G125), .Z(n1197) );
NOR2_X1 U853 ( .A1(n1082), .A2(G952), .ZN(n1120) );
XOR2_X1 U854 ( .A(n1198), .B(n1199), .Z(G48) );
NOR2_X1 U855 ( .A1(KEYINPUT35), .A2(n1200), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1201), .A2(n1171), .ZN(n1198) );
INV_X1 U857 ( .A(n1202), .ZN(n1171) );
XOR2_X1 U858 ( .A(G143), .B(n1167), .Z(G45) );
NOR4_X1 U859 ( .A1(n1203), .A2(n1204), .A3(n1186), .A4(n1185), .ZN(n1167) );
XNOR2_X1 U860 ( .A(G140), .B(n1104), .ZN(G42) );
NAND3_X1 U861 ( .A1(n1169), .A2(n1062), .A3(n1205), .ZN(n1104) );
XOR2_X1 U862 ( .A(n1162), .B(n1206), .Z(G39) );
XOR2_X1 U863 ( .A(KEYINPUT57), .B(G137), .Z(n1206) );
NAND4_X1 U864 ( .A1(n1169), .A2(n1062), .A3(n1207), .A4(n1061), .ZN(n1162) );
INV_X1 U865 ( .A(n1040), .ZN(n1062) );
NAND2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(G36) );
OR2_X1 U867 ( .A1(n1210), .A2(G134), .ZN(n1209) );
NAND2_X1 U868 ( .A1(G134), .A2(n1211), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
OR2_X1 U870 ( .A1(n1163), .A2(KEYINPUT46), .ZN(n1213) );
NAND2_X1 U871 ( .A1(KEYINPUT46), .A2(n1210), .ZN(n1212) );
NAND2_X1 U872 ( .A1(n1214), .A2(n1215), .ZN(n1210) );
INV_X1 U873 ( .A(n1163), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1169), .A2(n1047), .A3(n1057), .ZN(n1163) );
XNOR2_X1 U875 ( .A(KEYINPUT26), .B(KEYINPUT11), .ZN(n1214) );
XNOR2_X1 U876 ( .A(G131), .B(n1216), .ZN(G33) );
NAND4_X1 U877 ( .A1(n1057), .A2(n1048), .A3(n1052), .A4(n1217), .ZN(n1216) );
XNOR2_X1 U878 ( .A(KEYINPUT4), .B(n1218), .ZN(n1217) );
NOR3_X1 U879 ( .A1(n1203), .A2(n1219), .A3(n1040), .ZN(n1057) );
NAND2_X1 U880 ( .A1(n1068), .A2(n1220), .ZN(n1040) );
XNOR2_X1 U881 ( .A(G128), .B(n1221), .ZN(G30) );
NAND2_X1 U882 ( .A1(n1202), .A2(n1047), .ZN(n1221) );
NOR2_X1 U883 ( .A1(n1204), .A2(n1060), .ZN(n1202) );
NAND3_X1 U884 ( .A1(n1065), .A2(n1061), .A3(n1169), .ZN(n1204) );
AND2_X1 U885 ( .A1(n1052), .A2(n1218), .ZN(n1169) );
XNOR2_X1 U886 ( .A(n1194), .B(n1222), .ZN(G3) );
NAND2_X1 U887 ( .A1(KEYINPUT60), .A2(G101), .ZN(n1222) );
AND4_X1 U888 ( .A1(n1223), .A2(n1052), .A3(n1224), .A4(n1195), .ZN(n1194) );
NOR2_X1 U889 ( .A1(n1219), .A2(n1203), .ZN(n1224) );
INV_X1 U890 ( .A(n1060), .ZN(n1203) );
INV_X1 U891 ( .A(n1050), .ZN(n1223) );
NAND2_X1 U892 ( .A1(n1225), .A2(n1226), .ZN(G27) );
NAND2_X1 U893 ( .A1(G125), .A2(n1227), .ZN(n1226) );
NAND2_X1 U894 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U895 ( .A1(KEYINPUT45), .A2(n1230), .ZN(n1229) );
INV_X1 U896 ( .A(KEYINPUT55), .ZN(n1230) );
NAND3_X1 U897 ( .A1(n1231), .A2(n1232), .A3(KEYINPUT55), .ZN(n1225) );
OR2_X1 U898 ( .A1(n1164), .A2(KEYINPUT45), .ZN(n1232) );
NAND2_X1 U899 ( .A1(KEYINPUT45), .A2(n1233), .ZN(n1231) );
NAND2_X1 U900 ( .A1(n1228), .A2(n1234), .ZN(n1233) );
INV_X1 U901 ( .A(n1164), .ZN(n1228) );
NAND4_X1 U902 ( .A1(n1205), .A2(n1189), .A3(n1065), .A4(n1218), .ZN(n1164) );
NAND2_X1 U903 ( .A1(n1037), .A2(n1235), .ZN(n1218) );
NAND4_X1 U904 ( .A1(G902), .A2(G953), .A3(n1236), .A4(n1084), .ZN(n1235) );
INV_X1 U905 ( .A(G900), .ZN(n1084) );
INV_X1 U906 ( .A(n1046), .ZN(n1189) );
NOR3_X1 U907 ( .A1(n1061), .A2(n1060), .A3(n1201), .ZN(n1205) );
INV_X1 U908 ( .A(n1219), .ZN(n1061) );
XOR2_X1 U909 ( .A(n1237), .B(n1238), .Z(G24) );
NAND3_X1 U910 ( .A1(n1239), .A2(n1182), .A3(n1240), .ZN(n1238) );
NOR3_X1 U911 ( .A1(n1190), .A2(n1185), .A3(n1186), .ZN(n1240) );
INV_X1 U912 ( .A(n1042), .ZN(n1182) );
NAND2_X1 U913 ( .A1(n1219), .A2(n1060), .ZN(n1042) );
XOR2_X1 U914 ( .A(n1046), .B(KEYINPUT25), .Z(n1239) );
XOR2_X1 U915 ( .A(n1241), .B(G119), .Z(G21) );
NAND2_X1 U916 ( .A1(KEYINPUT30), .A2(n1193), .ZN(n1241) );
NAND2_X1 U917 ( .A1(n1242), .A2(n1207), .ZN(n1193) );
XOR2_X1 U918 ( .A(G116), .B(n1177), .Z(G18) );
AND3_X1 U919 ( .A1(n1060), .A2(n1047), .A3(n1242), .ZN(n1177) );
NOR2_X1 U920 ( .A1(n1243), .A2(n1186), .ZN(n1047) );
XOR2_X1 U921 ( .A(n1244), .B(n1173), .Z(G15) );
NAND3_X1 U922 ( .A1(n1060), .A2(n1242), .A3(n1048), .ZN(n1173) );
INV_X1 U923 ( .A(n1201), .ZN(n1048) );
NAND2_X1 U924 ( .A1(n1186), .A2(n1243), .ZN(n1201) );
INV_X1 U925 ( .A(n1185), .ZN(n1243) );
NOR3_X1 U926 ( .A1(n1190), .A2(n1219), .A3(n1046), .ZN(n1242) );
NAND2_X1 U927 ( .A1(n1245), .A2(n1246), .ZN(n1046) );
XOR2_X1 U928 ( .A(n1053), .B(KEYINPUT38), .Z(n1245) );
XOR2_X1 U929 ( .A(n1247), .B(n1174), .Z(G12) );
NAND4_X1 U930 ( .A1(n1207), .A2(n1052), .A3(n1195), .A4(n1219), .ZN(n1174) );
NOR2_X1 U931 ( .A1(n1248), .A2(n1071), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1074), .A2(G472), .ZN(n1071) );
AND2_X1 U933 ( .A1(n1249), .A2(n1074), .ZN(n1248) );
NAND2_X1 U934 ( .A1(n1250), .A2(n1251), .ZN(n1074) );
XOR2_X1 U935 ( .A(n1252), .B(n1253), .Z(n1250) );
XOR2_X1 U936 ( .A(n1142), .B(n1254), .Z(n1253) );
XOR2_X1 U937 ( .A(n1255), .B(n1244), .Z(n1142) );
XOR2_X1 U938 ( .A(n1256), .B(n1257), .Z(n1252) );
NOR2_X1 U939 ( .A1(KEYINPUT18), .A2(n1143), .ZN(n1257) );
NAND2_X1 U940 ( .A1(n1258), .A2(KEYINPUT41), .ZN(n1256) );
XOR2_X1 U941 ( .A(n1146), .B(G101), .Z(n1258) );
NAND2_X1 U942 ( .A1(G210), .A2(n1259), .ZN(n1146) );
XOR2_X1 U943 ( .A(n1148), .B(KEYINPUT1), .Z(n1249) );
INV_X1 U944 ( .A(G472), .ZN(n1148) );
INV_X1 U945 ( .A(n1190), .ZN(n1195) );
NAND2_X1 U946 ( .A1(n1065), .A2(n1183), .ZN(n1190) );
NAND2_X1 U947 ( .A1(n1037), .A2(n1260), .ZN(n1183) );
NAND3_X1 U948 ( .A1(n1116), .A2(n1236), .A3(G902), .ZN(n1260) );
NOR2_X1 U949 ( .A1(n1082), .A2(G898), .ZN(n1116) );
NAND3_X1 U950 ( .A1(n1236), .A2(n1082), .A3(G952), .ZN(n1037) );
NAND2_X1 U951 ( .A1(G237), .A2(G234), .ZN(n1236) );
INV_X1 U952 ( .A(n1181), .ZN(n1065) );
NAND2_X1 U953 ( .A1(n1220), .A2(n1067), .ZN(n1181) );
INV_X1 U954 ( .A(n1068), .ZN(n1067) );
XNOR2_X1 U955 ( .A(n1261), .B(n1160), .ZN(n1068) );
NAND2_X1 U956 ( .A1(G210), .A2(n1262), .ZN(n1160) );
NAND2_X1 U957 ( .A1(n1263), .A2(n1251), .ZN(n1261) );
XOR2_X1 U958 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U959 ( .A(n1266), .B(n1143), .Z(n1265) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1143) );
INV_X1 U961 ( .A(n1269), .ZN(n1268) );
XOR2_X1 U962 ( .A(G143), .B(n1200), .Z(n1267) );
NAND2_X1 U963 ( .A1(KEYINPUT29), .A2(n1157), .ZN(n1266) );
XNOR2_X1 U964 ( .A(n1270), .B(n1119), .ZN(n1157) );
XNOR2_X1 U965 ( .A(n1271), .B(n1272), .ZN(n1119) );
XOR2_X1 U966 ( .A(KEYINPUT61), .B(G113), .Z(n1272) );
XOR2_X1 U967 ( .A(n1273), .B(n1274), .Z(n1271) );
NAND2_X1 U968 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U970 ( .A(KEYINPUT6), .ZN(n1278) );
XOR2_X1 U971 ( .A(n1279), .B(G101), .Z(n1277) );
NAND2_X1 U972 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U973 ( .A1(n1282), .A2(KEYINPUT6), .ZN(n1275) );
XOR2_X1 U974 ( .A(G101), .B(n1255), .Z(n1282) );
XNOR2_X1 U975 ( .A(n1281), .B(n1280), .ZN(n1255) );
XOR2_X1 U976 ( .A(G116), .B(KEYINPUT27), .Z(n1280) );
NAND2_X1 U977 ( .A1(KEYINPUT21), .A2(n1118), .ZN(n1270) );
XOR2_X1 U978 ( .A(G110), .B(G122), .Z(n1118) );
XOR2_X1 U979 ( .A(n1196), .B(n1283), .Z(n1264) );
NOR2_X1 U980 ( .A1(KEYINPUT37), .A2(n1234), .ZN(n1283) );
INV_X1 U981 ( .A(G125), .ZN(n1234) );
AND2_X1 U982 ( .A1(G224), .A2(n1082), .ZN(n1196) );
XOR2_X1 U983 ( .A(n1072), .B(KEYINPUT23), .Z(n1220) );
INV_X1 U984 ( .A(n1066), .ZN(n1072) );
NAND2_X1 U985 ( .A1(G214), .A2(n1262), .ZN(n1066) );
NAND2_X1 U986 ( .A1(n1284), .A2(n1251), .ZN(n1262) );
INV_X1 U987 ( .A(G237), .ZN(n1284) );
NOR2_X1 U988 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U989 ( .A(n1246), .ZN(n1054) );
NAND2_X1 U990 ( .A1(G221), .A2(n1285), .ZN(n1246) );
XOR2_X1 U991 ( .A(n1286), .B(n1287), .Z(n1053) );
XNOR2_X1 U992 ( .A(KEYINPUT42), .B(n1076), .ZN(n1287) );
NAND2_X1 U993 ( .A1(n1288), .A2(n1251), .ZN(n1076) );
XOR2_X1 U994 ( .A(n1153), .B(n1289), .Z(n1288) );
XOR2_X1 U995 ( .A(KEYINPUT54), .B(KEYINPUT3), .Z(n1289) );
XOR2_X1 U996 ( .A(n1290), .B(n1291), .Z(n1153) );
XOR2_X1 U997 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U998 ( .A(G110), .B(n1294), .Z(n1293) );
NOR2_X1 U999 ( .A1(G953), .A2(n1083), .ZN(n1294) );
INV_X1 U1000 ( .A(G227), .ZN(n1083) );
XOR2_X1 U1001 ( .A(KEYINPUT24), .B(G140), .Z(n1292) );
XOR2_X1 U1002 ( .A(n1101), .B(n1295), .Z(n1290) );
XNOR2_X1 U1003 ( .A(n1274), .B(n1140), .ZN(n1295) );
XNOR2_X1 U1004 ( .A(n1254), .B(G101), .ZN(n1140) );
XOR2_X1 U1005 ( .A(G131), .B(n1100), .Z(n1254) );
XOR2_X1 U1006 ( .A(G137), .B(G134), .Z(n1100) );
XOR2_X1 U1007 ( .A(G104), .B(n1296), .Z(n1274) );
XOR2_X1 U1008 ( .A(n1269), .B(n1297), .Z(n1101) );
XNOR2_X1 U1009 ( .A(n1298), .B(KEYINPUT39), .ZN(n1297) );
NAND2_X1 U1010 ( .A1(n1299), .A2(KEYINPUT51), .ZN(n1298) );
XOR2_X1 U1011 ( .A(n1200), .B(n1300), .Z(n1299) );
NOR2_X1 U1012 ( .A1(KEYINPUT40), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U1013 ( .A(G143), .B(KEYINPUT5), .ZN(n1301) );
INV_X1 U1014 ( .A(G146), .ZN(n1200) );
NAND2_X1 U1015 ( .A1(KEYINPUT52), .A2(n1078), .ZN(n1286) );
INV_X1 U1016 ( .A(G469), .ZN(n1078) );
NOR2_X1 U1017 ( .A1(n1050), .A2(n1060), .ZN(n1207) );
XNOR2_X1 U1018 ( .A(n1302), .B(n1124), .ZN(n1060) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1285), .ZN(n1124) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1251), .ZN(n1285) );
NAND2_X1 U1021 ( .A1(n1122), .A2(n1251), .ZN(n1302) );
INV_X1 U1022 ( .A(G902), .ZN(n1251) );
XNOR2_X1 U1023 ( .A(n1303), .B(n1304), .ZN(n1122) );
XNOR2_X1 U1024 ( .A(n1305), .B(n1102), .ZN(n1304) );
XOR2_X1 U1025 ( .A(G140), .B(G125), .Z(n1102) );
NAND2_X1 U1026 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
OR2_X1 U1027 ( .A1(n1308), .A2(n1247), .ZN(n1307) );
XOR2_X1 U1028 ( .A(n1309), .B(KEYINPUT2), .Z(n1306) );
NAND2_X1 U1029 ( .A1(n1308), .A2(n1247), .ZN(n1309) );
XOR2_X1 U1030 ( .A(n1281), .B(n1269), .Z(n1308) );
INV_X1 U1031 ( .A(G119), .ZN(n1281) );
XOR2_X1 U1032 ( .A(n1310), .B(n1311), .Z(n1303) );
XOR2_X1 U1033 ( .A(G146), .B(G137), .Z(n1311) );
NAND2_X1 U1034 ( .A1(n1312), .A2(G221), .ZN(n1310) );
NAND2_X1 U1035 ( .A1(n1186), .A2(n1185), .ZN(n1050) );
XOR2_X1 U1036 ( .A(n1313), .B(G475), .Z(n1185) );
OR2_X1 U1037 ( .A1(n1132), .A2(G902), .ZN(n1313) );
XNOR2_X1 U1038 ( .A(n1314), .B(n1315), .ZN(n1132) );
XOR2_X1 U1039 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND3_X1 U1040 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1317) );
NAND2_X1 U1041 ( .A1(G140), .A2(n1321), .ZN(n1320) );
OR3_X1 U1042 ( .A1(n1321), .A2(G140), .A3(KEYINPUT10), .ZN(n1319) );
OR2_X1 U1043 ( .A1(G125), .A2(KEYINPUT49), .ZN(n1321) );
NAND2_X1 U1044 ( .A1(KEYINPUT10), .A2(G125), .ZN(n1318) );
NAND2_X1 U1045 ( .A1(KEYINPUT43), .A2(n1322), .ZN(n1316) );
XNOR2_X1 U1046 ( .A(G104), .B(n1323), .ZN(n1322) );
NAND3_X1 U1047 ( .A1(n1324), .A2(n1325), .A3(n1326), .ZN(n1323) );
NAND2_X1 U1048 ( .A1(G113), .A2(n1237), .ZN(n1326) );
NAND2_X1 U1049 ( .A1(KEYINPUT63), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1050 ( .A1(n1328), .A2(n1244), .ZN(n1327) );
XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n1237), .Z(n1328) );
NAND2_X1 U1052 ( .A1(n1329), .A2(n1330), .ZN(n1324) );
INV_X1 U1053 ( .A(KEYINPUT63), .ZN(n1330) );
NAND2_X1 U1054 ( .A1(n1331), .A2(n1332), .ZN(n1329) );
OR2_X1 U1055 ( .A1(G122), .A2(KEYINPUT53), .ZN(n1332) );
NAND3_X1 U1056 ( .A1(G122), .A2(n1244), .A3(KEYINPUT53), .ZN(n1331) );
INV_X1 U1057 ( .A(G113), .ZN(n1244) );
XOR2_X1 U1058 ( .A(n1333), .B(G146), .Z(n1314) );
NAND2_X1 U1059 ( .A1(KEYINPUT36), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1060 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1061 ( .A(G131), .B(G143), .ZN(n1336) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1259), .ZN(n1335) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1259) );
XOR2_X1 U1064 ( .A(n1337), .B(G478), .Z(n1186) );
OR2_X1 U1065 ( .A1(n1128), .A2(G902), .ZN(n1337) );
XNOR2_X1 U1066 ( .A(n1338), .B(n1339), .ZN(n1128) );
XOR2_X1 U1067 ( .A(n1340), .B(n1341), .Z(n1339) );
NAND2_X1 U1068 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1069 ( .A1(G122), .A2(n1344), .ZN(n1343) );
INV_X1 U1070 ( .A(G116), .ZN(n1344) );
XOR2_X1 U1071 ( .A(n1345), .B(KEYINPUT31), .Z(n1342) );
NAND2_X1 U1072 ( .A1(G116), .A2(n1237), .ZN(n1345) );
INV_X1 U1073 ( .A(G122), .ZN(n1237) );
NAND2_X1 U1074 ( .A1(n1346), .A2(n1312), .ZN(n1340) );
AND2_X1 U1075 ( .A1(G234), .A2(n1082), .ZN(n1312) );
INV_X1 U1076 ( .A(G953), .ZN(n1082) );
XNOR2_X1 U1077 ( .A(G217), .B(KEYINPUT28), .ZN(n1346) );
XNOR2_X1 U1078 ( .A(n1347), .B(n1348), .ZN(n1338) );
NAND2_X1 U1079 ( .A1(KEYINPUT50), .A2(n1296), .ZN(n1348) );
XOR2_X1 U1080 ( .A(G107), .B(KEYINPUT8), .Z(n1296) );
NAND2_X1 U1081 ( .A1(n1349), .A2(KEYINPUT19), .ZN(n1347) );
XOR2_X1 U1082 ( .A(n1269), .B(n1350), .Z(n1349) );
XOR2_X1 U1083 ( .A(G134), .B(n1351), .Z(n1350) );
NOR2_X1 U1084 ( .A1(G143), .A2(KEYINPUT16), .ZN(n1351) );
XNOR2_X1 U1085 ( .A(G128), .B(KEYINPUT0), .ZN(n1269) );
INV_X1 U1086 ( .A(G110), .ZN(n1247) );
endmodule


