//Key = 1110010010000111110100110111111010110010000110010010111011011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430, n1431;

XNOR2_X1 U783 ( .A(G107), .B(n1085), .ZN(G9) );
NOR2_X1 U784 ( .A1(n1086), .A2(n1087), .ZN(G75) );
AND3_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NOR3_X1 U786 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1086) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR3_X1 U788 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1094) );
NOR3_X1 U789 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1097) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U796 ( .A1(KEYINPUT31), .A2(n1115), .ZN(n1113) );
NOR2_X1 U797 ( .A1(n1116), .A2(n1101), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1096) );
INV_X1 U800 ( .A(KEYINPUT31), .ZN(n1120) );
NOR3_X1 U801 ( .A1(n1115), .A2(n1099), .A3(n1106), .ZN(n1119) );
INV_X1 U802 ( .A(n1121), .ZN(n1106) );
INV_X1 U803 ( .A(n1122), .ZN(n1099) );
INV_X1 U804 ( .A(n1123), .ZN(n1115) );
NAND3_X1 U805 ( .A1(n1124), .A2(n1089), .A3(n1088), .ZN(n1091) );
NAND4_X1 U806 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1088) );
NOR3_X1 U807 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
XNOR2_X1 U808 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U809 ( .A1(KEYINPUT30), .A2(n1134), .ZN(n1132) );
NOR2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NAND3_X1 U811 ( .A1(n1105), .A2(n1137), .A3(n1138), .ZN(n1129) );
NOR3_X1 U812 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U814 ( .A(KEYINPUT36), .B(n1144), .Z(n1143) );
NOR2_X1 U815 ( .A1(G478), .A2(n1145), .ZN(n1140) );
XNOR2_X1 U816 ( .A(n1144), .B(KEYINPUT55), .ZN(n1145) );
XNOR2_X1 U817 ( .A(KEYINPUT58), .B(n1146), .ZN(n1139) );
XOR2_X1 U818 ( .A(KEYINPUT17), .B(n1147), .Z(n1126) );
NAND4_X1 U819 ( .A1(n1121), .A2(n1122), .A3(n1148), .A4(n1149), .ZN(n1124) );
NAND2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
OR2_X1 U821 ( .A1(n1137), .A2(n1152), .ZN(n1151) );
NOR2_X1 U822 ( .A1(n1108), .A2(n1112), .ZN(n1122) );
XOR2_X1 U823 ( .A(n1153), .B(n1154), .Z(G72) );
XOR2_X1 U824 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND3_X1 U825 ( .A1(n1157), .A2(n1089), .A3(KEYINPUT56), .ZN(n1156) );
NAND2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1155) );
NAND2_X1 U827 ( .A1(G953), .A2(n1160), .ZN(n1159) );
XOR2_X1 U828 ( .A(n1161), .B(n1162), .Z(n1158) );
XOR2_X1 U829 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U830 ( .A(n1165), .B(n1166), .ZN(n1161) );
XNOR2_X1 U831 ( .A(KEYINPUT0), .B(n1167), .ZN(n1166) );
NOR2_X1 U832 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1167) );
XNOR2_X1 U833 ( .A(G146), .B(n1169), .ZN(n1168) );
NOR3_X1 U834 ( .A1(n1089), .A2(KEYINPUT39), .A3(n1170), .ZN(n1153) );
AND2_X1 U835 ( .A1(G227), .A2(G900), .ZN(n1170) );
NAND2_X1 U836 ( .A1(n1171), .A2(n1172), .ZN(G69) );
NAND2_X1 U837 ( .A1(G953), .A2(n1173), .ZN(n1172) );
NAND2_X1 U838 ( .A1(n1174), .A2(G898), .ZN(n1173) );
XNOR2_X1 U839 ( .A(n1175), .B(G224), .ZN(n1174) );
NAND2_X1 U840 ( .A1(n1176), .A2(n1089), .ZN(n1171) );
XNOR2_X1 U841 ( .A(n1177), .B(n1178), .ZN(n1176) );
INV_X1 U842 ( .A(n1175), .ZN(n1178) );
XOR2_X1 U843 ( .A(n1179), .B(n1180), .Z(n1175) );
NOR2_X1 U844 ( .A1(KEYINPUT42), .A2(n1181), .ZN(n1180) );
XNOR2_X1 U845 ( .A(G122), .B(n1182), .ZN(n1181) );
NAND2_X1 U846 ( .A1(KEYINPUT44), .A2(n1183), .ZN(n1177) );
NAND2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U848 ( .A(n1186), .B(KEYINPUT24), .Z(n1184) );
NOR3_X1 U849 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(G66) );
AND2_X1 U850 ( .A1(KEYINPUT14), .A2(n1190), .ZN(n1189) );
NOR3_X1 U851 ( .A1(KEYINPUT14), .A2(n1089), .A3(n1090), .ZN(n1188) );
INV_X1 U852 ( .A(G952), .ZN(n1090) );
XOR2_X1 U853 ( .A(n1191), .B(n1192), .Z(n1187) );
NOR2_X1 U854 ( .A1(n1136), .A2(n1193), .ZN(n1192) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1194), .ZN(G63) );
NOR3_X1 U856 ( .A1(n1144), .A2(n1195), .A3(n1196), .ZN(n1194) );
NOR3_X1 U857 ( .A1(n1197), .A2(n1142), .A3(n1193), .ZN(n1196) );
INV_X1 U858 ( .A(G478), .ZN(n1142) );
NOR2_X1 U859 ( .A1(n1198), .A2(n1199), .ZN(n1195) );
AND2_X1 U860 ( .A1(n1093), .A2(G478), .ZN(n1198) );
NOR2_X1 U861 ( .A1(n1190), .A2(n1200), .ZN(G60) );
XOR2_X1 U862 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND3_X1 U863 ( .A1(n1203), .A2(n1093), .A3(G475), .ZN(n1202) );
XNOR2_X1 U864 ( .A(KEYINPUT18), .B(n1204), .ZN(n1203) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(G6) );
XOR2_X1 U866 ( .A(KEYINPUT9), .B(G104), .Z(n1206) );
NOR3_X1 U867 ( .A1(n1150), .A2(KEYINPUT45), .A3(n1207), .ZN(n1205) );
XNOR2_X1 U868 ( .A(n1208), .B(KEYINPUT4), .ZN(n1207) );
NOR2_X1 U869 ( .A1(n1190), .A2(n1209), .ZN(G57) );
NOR2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U871 ( .A(KEYINPUT7), .B(n1212), .Z(n1211) );
NOR2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
AND2_X1 U873 ( .A1(n1214), .A2(n1213), .ZN(n1210) );
XOR2_X1 U874 ( .A(n1215), .B(G101), .Z(n1213) );
NAND2_X1 U875 ( .A1(KEYINPUT28), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U876 ( .A(n1217), .B(n1218), .ZN(n1214) );
NOR2_X1 U877 ( .A1(n1219), .A2(n1193), .ZN(n1218) );
NOR2_X1 U878 ( .A1(n1190), .A2(n1220), .ZN(G54) );
XOR2_X1 U879 ( .A(n1221), .B(n1222), .Z(n1220) );
NOR2_X1 U880 ( .A1(n1223), .A2(n1193), .ZN(n1222) );
NOR2_X1 U881 ( .A1(n1224), .A2(n1225), .ZN(n1221) );
XOR2_X1 U882 ( .A(KEYINPUT48), .B(n1226), .Z(n1225) );
NOR2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
AND2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1224) );
XOR2_X1 U885 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U886 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
INV_X1 U887 ( .A(n1233), .ZN(n1232) );
XOR2_X1 U888 ( .A(KEYINPUT23), .B(n1234), .Z(n1231) );
NOR3_X1 U889 ( .A1(n1190), .A2(n1235), .A3(n1236), .ZN(G51) );
NOR2_X1 U890 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
INV_X1 U891 ( .A(KEYINPUT51), .ZN(n1238) );
XOR2_X1 U892 ( .A(n1239), .B(n1240), .Z(n1237) );
NAND2_X1 U893 ( .A1(KEYINPUT54), .A2(n1241), .ZN(n1239) );
NOR2_X1 U894 ( .A1(KEYINPUT51), .A2(n1242), .ZN(n1235) );
XOR2_X1 U895 ( .A(n1243), .B(n1240), .Z(n1242) );
XNOR2_X1 U896 ( .A(n1244), .B(n1245), .ZN(n1240) );
NOR2_X1 U897 ( .A1(n1134), .A2(n1193), .ZN(n1245) );
NAND2_X1 U898 ( .A1(G902), .A2(n1093), .ZN(n1193) );
NAND3_X1 U899 ( .A1(n1185), .A2(n1186), .A3(n1246), .ZN(n1093) );
INV_X1 U900 ( .A(n1157), .ZN(n1246) );
NAND4_X1 U901 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1157) );
AND4_X1 U902 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
NAND3_X1 U903 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1249) );
NAND2_X1 U904 ( .A1(n1258), .A2(n1150), .ZN(n1256) );
NAND2_X1 U905 ( .A1(n1117), .A2(n1259), .ZN(n1258) );
INV_X1 U906 ( .A(KEYINPUT1), .ZN(n1259) );
NAND3_X1 U907 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1255) );
NAND2_X1 U908 ( .A1(KEYINPUT1), .A2(n1117), .ZN(n1260) );
NAND3_X1 U909 ( .A1(n1263), .A2(n1103), .A3(n1264), .ZN(n1247) );
NAND2_X1 U910 ( .A1(n1265), .A2(n1262), .ZN(n1186) );
XOR2_X1 U911 ( .A(n1266), .B(KEYINPUT8), .Z(n1265) );
AND4_X1 U912 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1185) );
AND3_X1 U913 ( .A1(n1271), .A2(n1085), .A3(n1272), .ZN(n1270) );
NAND4_X1 U914 ( .A1(n1273), .A2(n1148), .A3(n1103), .A4(n1117), .ZN(n1085) );
NAND2_X1 U915 ( .A1(n1208), .A2(n1262), .ZN(n1269) );
NOR4_X1 U916 ( .A1(n1261), .A2(n1101), .A3(n1274), .A4(n1275), .ZN(n1208) );
NAND4_X1 U917 ( .A1(n1276), .A2(n1277), .A3(n1121), .A4(n1278), .ZN(n1268) );
NOR2_X1 U918 ( .A1(n1279), .A2(n1101), .ZN(n1278) );
OR2_X1 U919 ( .A1(n1280), .A2(n1273), .ZN(n1277) );
NAND2_X1 U920 ( .A1(n1281), .A2(n1280), .ZN(n1276) );
INV_X1 U921 ( .A(KEYINPUT22), .ZN(n1280) );
NAND2_X1 U922 ( .A1(n1282), .A2(n1150), .ZN(n1281) );
NAND3_X1 U923 ( .A1(n1273), .A2(n1283), .A3(n1284), .ZN(n1267) );
NAND3_X1 U924 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1283) );
NAND2_X1 U925 ( .A1(KEYINPUT53), .A2(n1288), .ZN(n1287) );
NAND3_X1 U926 ( .A1(n1114), .A2(n1289), .A3(n1274), .ZN(n1286) );
INV_X1 U927 ( .A(KEYINPUT53), .ZN(n1289) );
NAND2_X1 U928 ( .A1(n1123), .A2(n1103), .ZN(n1285) );
NAND2_X1 U929 ( .A1(n1290), .A2(n1291), .ZN(n1244) );
NAND2_X1 U930 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U931 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U932 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
XNOR2_X1 U933 ( .A(G125), .B(n1298), .ZN(n1296) );
XNOR2_X1 U934 ( .A(KEYINPUT50), .B(KEYINPUT25), .ZN(n1298) );
NAND2_X1 U935 ( .A1(n1299), .A2(n1300), .ZN(n1290) );
NAND2_X1 U936 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
OR2_X1 U937 ( .A1(n1303), .A2(n1295), .ZN(n1302) );
NAND2_X1 U938 ( .A1(n1304), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U939 ( .A(n1297), .B(n1295), .ZN(n1304) );
XNOR2_X1 U940 ( .A(n1305), .B(KEYINPUT61), .ZN(n1295) );
INV_X1 U941 ( .A(KEYINPUT41), .ZN(n1297) );
NAND2_X1 U942 ( .A1(KEYINPUT54), .A2(n1306), .ZN(n1243) );
NOR2_X1 U943 ( .A1(n1089), .A2(G952), .ZN(n1190) );
NAND2_X1 U944 ( .A1(n1307), .A2(n1308), .ZN(G48) );
NAND2_X1 U945 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U946 ( .A(KEYINPUT62), .B(n1311), .Z(n1307) );
NOR2_X1 U947 ( .A1(n1309), .A2(n1310), .ZN(n1311) );
AND4_X1 U948 ( .A1(n1118), .A2(n1262), .A3(n1312), .A4(n1313), .ZN(n1309) );
OR2_X1 U949 ( .A1(n1257), .A2(KEYINPUT21), .ZN(n1313) );
NAND2_X1 U950 ( .A1(KEYINPUT21), .A2(n1314), .ZN(n1312) );
NAND2_X1 U951 ( .A1(n1315), .A2(n1274), .ZN(n1314) );
XNOR2_X1 U952 ( .A(G143), .B(n1248), .ZN(G45) );
NAND3_X1 U953 ( .A1(n1262), .A2(n1316), .A3(n1317), .ZN(n1248) );
XNOR2_X1 U954 ( .A(G140), .B(n1318), .ZN(G42) );
NAND3_X1 U955 ( .A1(n1264), .A2(n1263), .A3(n1319), .ZN(n1318) );
XNOR2_X1 U956 ( .A(n1103), .B(KEYINPUT13), .ZN(n1319) );
XNOR2_X1 U957 ( .A(n1254), .B(n1320), .ZN(G39) );
NOR2_X1 U958 ( .A1(KEYINPUT49), .A2(n1321), .ZN(n1320) );
NAND3_X1 U959 ( .A1(n1264), .A2(n1284), .A3(n1257), .ZN(n1254) );
XNOR2_X1 U960 ( .A(G134), .B(n1253), .ZN(G36) );
NAND3_X1 U961 ( .A1(n1317), .A2(n1117), .A3(n1264), .ZN(n1253) );
XNOR2_X1 U962 ( .A(G131), .B(n1252), .ZN(G33) );
NAND3_X1 U963 ( .A1(n1317), .A2(n1118), .A3(n1264), .ZN(n1252) );
INV_X1 U964 ( .A(n1095), .ZN(n1264) );
NAND2_X1 U965 ( .A1(n1322), .A2(n1137), .ZN(n1095) );
INV_X1 U966 ( .A(n1152), .ZN(n1322) );
AND2_X1 U967 ( .A1(n1288), .A2(n1323), .ZN(n1317) );
XNOR2_X1 U968 ( .A(G128), .B(n1324), .ZN(G30) );
NAND3_X1 U969 ( .A1(n1117), .A2(n1262), .A3(n1257), .ZN(n1324) );
AND2_X1 U970 ( .A1(n1315), .A2(n1103), .ZN(n1257) );
AND3_X1 U971 ( .A1(n1323), .A2(n1325), .A3(n1326), .ZN(n1315) );
XNOR2_X1 U972 ( .A(G101), .B(n1327), .ZN(G3) );
NAND3_X1 U973 ( .A1(n1284), .A2(n1273), .A3(n1288), .ZN(n1327) );
AND2_X1 U974 ( .A1(n1103), .A2(n1114), .ZN(n1288) );
XNOR2_X1 U975 ( .A(G125), .B(n1251), .ZN(G27) );
NAND3_X1 U976 ( .A1(n1121), .A2(n1262), .A3(n1263), .ZN(n1251) );
AND3_X1 U977 ( .A1(n1118), .A2(n1323), .A3(n1123), .ZN(n1263) );
NAND2_X1 U978 ( .A1(n1108), .A2(n1328), .ZN(n1323) );
NAND4_X1 U979 ( .A1(G953), .A2(G902), .A3(n1329), .A4(n1160), .ZN(n1328) );
INV_X1 U980 ( .A(G900), .ZN(n1160) );
INV_X1 U981 ( .A(n1150), .ZN(n1262) );
XOR2_X1 U982 ( .A(G122), .B(n1330), .Z(G24) );
NOR3_X1 U983 ( .A1(n1331), .A2(n1279), .A3(n1101), .ZN(n1330) );
INV_X1 U984 ( .A(n1316), .ZN(n1279) );
NAND2_X1 U985 ( .A1(n1332), .A2(n1333), .ZN(n1316) );
OR2_X1 U986 ( .A1(n1261), .A2(KEYINPUT19), .ZN(n1333) );
NAND2_X1 U987 ( .A1(KEYINPUT19), .A2(n1334), .ZN(n1332) );
NAND2_X1 U988 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
OR3_X1 U989 ( .A1(n1337), .A2(n1146), .A3(KEYINPUT20), .ZN(n1336) );
NAND2_X1 U990 ( .A1(KEYINPUT20), .A2(n1117), .ZN(n1335) );
XOR2_X1 U991 ( .A(G119), .B(n1338), .Z(G21) );
NOR2_X1 U992 ( .A1(n1150), .A2(n1266), .ZN(n1338) );
NAND3_X1 U993 ( .A1(n1121), .A2(n1284), .A3(n1339), .ZN(n1266) );
NOR3_X1 U994 ( .A1(n1125), .A2(n1275), .A3(n1340), .ZN(n1339) );
INV_X1 U995 ( .A(n1326), .ZN(n1125) );
XNOR2_X1 U996 ( .A(G116), .B(n1271), .ZN(G18) );
NAND3_X1 U997 ( .A1(n1117), .A2(n1114), .A3(n1341), .ZN(n1271) );
NOR2_X1 U998 ( .A1(n1342), .A2(n1337), .ZN(n1117) );
XNOR2_X1 U999 ( .A(G113), .B(n1272), .ZN(G15) );
NAND3_X1 U1000 ( .A1(n1118), .A2(n1114), .A3(n1341), .ZN(n1272) );
INV_X1 U1001 ( .A(n1331), .ZN(n1341) );
NAND2_X1 U1002 ( .A1(n1121), .A2(n1273), .ZN(n1331) );
NOR2_X1 U1003 ( .A1(n1104), .A2(n1343), .ZN(n1121) );
INV_X1 U1004 ( .A(n1105), .ZN(n1343) );
NAND2_X1 U1005 ( .A1(n1344), .A2(n1345), .ZN(n1114) );
OR2_X1 U1006 ( .A1(n1101), .A2(KEYINPUT60), .ZN(n1345) );
INV_X1 U1007 ( .A(n1148), .ZN(n1101) );
NOR2_X1 U1008 ( .A1(n1325), .A2(n1326), .ZN(n1148) );
NAND3_X1 U1009 ( .A1(n1340), .A2(n1326), .A3(KEYINPUT60), .ZN(n1344) );
INV_X1 U1010 ( .A(n1261), .ZN(n1118) );
NAND2_X1 U1011 ( .A1(n1337), .A2(n1346), .ZN(n1261) );
XNOR2_X1 U1012 ( .A(KEYINPUT20), .B(n1146), .ZN(n1346) );
XNOR2_X1 U1013 ( .A(G110), .B(n1347), .ZN(G12) );
NAND4_X1 U1014 ( .A1(n1348), .A2(n1284), .A3(n1273), .A4(n1103), .ZN(n1347) );
INV_X1 U1015 ( .A(n1274), .ZN(n1103) );
NAND2_X1 U1016 ( .A1(n1104), .A2(n1105), .ZN(n1274) );
NAND2_X1 U1017 ( .A1(G221), .A2(n1349), .ZN(n1105) );
XNOR2_X1 U1018 ( .A(n1147), .B(KEYINPUT38), .ZN(n1104) );
XOR2_X1 U1019 ( .A(n1350), .B(n1223), .Z(n1147) );
INV_X1 U1020 ( .A(G469), .ZN(n1223) );
NAND2_X1 U1021 ( .A1(n1351), .A2(n1204), .ZN(n1350) );
XNOR2_X1 U1022 ( .A(n1227), .B(n1352), .ZN(n1351) );
XOR2_X1 U1023 ( .A(n1353), .B(KEYINPUT16), .Z(n1352) );
NAND2_X1 U1024 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1025 ( .A1(n1356), .A2(n1230), .ZN(n1355) );
OR2_X1 U1026 ( .A1(n1234), .A2(n1233), .ZN(n1356) );
XOR2_X1 U1027 ( .A(KEYINPUT35), .B(n1357), .Z(n1354) );
NOR3_X1 U1028 ( .A1(n1230), .A2(n1234), .A3(n1233), .ZN(n1357) );
NOR2_X1 U1029 ( .A1(n1182), .A2(G140), .ZN(n1233) );
AND2_X1 U1030 ( .A1(G140), .A2(n1182), .ZN(n1234) );
INV_X1 U1031 ( .A(G110), .ZN(n1182) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1089), .ZN(n1230) );
XNOR2_X1 U1033 ( .A(n1358), .B(n1359), .ZN(n1227) );
XOR2_X1 U1034 ( .A(G143), .B(n1163), .Z(n1359) );
XOR2_X1 U1035 ( .A(n1360), .B(n1361), .Z(n1358) );
NOR2_X1 U1036 ( .A1(n1150), .A2(n1275), .ZN(n1273) );
INV_X1 U1037 ( .A(n1282), .ZN(n1275) );
NAND2_X1 U1038 ( .A1(n1108), .A2(n1362), .ZN(n1282) );
NAND4_X1 U1039 ( .A1(G953), .A2(G902), .A3(n1329), .A4(n1363), .ZN(n1362) );
INV_X1 U1040 ( .A(G898), .ZN(n1363) );
NAND3_X1 U1041 ( .A1(n1329), .A2(n1089), .A3(G952), .ZN(n1108) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1329) );
NAND2_X1 U1043 ( .A1(n1152), .A2(n1137), .ZN(n1150) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1364), .ZN(n1137) );
XOR2_X1 U1045 ( .A(n1133), .B(n1134), .Z(n1152) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1364), .ZN(n1134) );
NAND2_X1 U1047 ( .A1(n1365), .A2(n1204), .ZN(n1364) );
NAND2_X1 U1048 ( .A1(n1366), .A2(n1204), .ZN(n1133) );
XNOR2_X1 U1049 ( .A(n1367), .B(n1241), .ZN(n1366) );
INV_X1 U1050 ( .A(n1306), .ZN(n1241) );
XOR2_X1 U1051 ( .A(n1368), .B(n1369), .Z(n1306) );
INV_X1 U1052 ( .A(n1179), .ZN(n1369) );
XNOR2_X1 U1053 ( .A(n1370), .B(n1371), .ZN(n1179) );
XNOR2_X1 U1054 ( .A(n1361), .B(KEYINPUT3), .ZN(n1370) );
XOR2_X1 U1055 ( .A(G101), .B(n1372), .Z(n1361) );
XOR2_X1 U1056 ( .A(G107), .B(G104), .Z(n1372) );
NAND2_X1 U1057 ( .A1(n1373), .A2(KEYINPUT2), .ZN(n1368) );
XNOR2_X1 U1058 ( .A(G110), .B(G122), .ZN(n1373) );
XOR2_X1 U1059 ( .A(n1374), .B(KEYINPUT26), .Z(n1367) );
NAND2_X1 U1060 ( .A1(n1375), .A2(KEYINPUT57), .ZN(n1374) );
XNOR2_X1 U1061 ( .A(n1292), .B(n1376), .ZN(n1375) );
XNOR2_X1 U1062 ( .A(G125), .B(n1305), .ZN(n1376) );
NAND2_X1 U1063 ( .A1(G224), .A2(n1089), .ZN(n1305) );
INV_X1 U1064 ( .A(n1300), .ZN(n1292) );
XOR2_X1 U1065 ( .A(n1377), .B(n1378), .Z(n1300) );
INV_X1 U1066 ( .A(n1112), .ZN(n1284) );
NAND2_X1 U1067 ( .A1(n1337), .A2(n1146), .ZN(n1112) );
INV_X1 U1068 ( .A(n1342), .ZN(n1146) );
XNOR2_X1 U1069 ( .A(n1379), .B(G475), .ZN(n1342) );
NAND2_X1 U1070 ( .A1(n1204), .A2(n1201), .ZN(n1379) );
NAND2_X1 U1071 ( .A1(n1380), .A2(n1381), .ZN(n1201) );
NAND2_X1 U1072 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
XOR2_X1 U1073 ( .A(n1384), .B(n1385), .Z(n1383) );
XOR2_X1 U1074 ( .A(n1386), .B(G104), .Z(n1382) );
XOR2_X1 U1075 ( .A(n1387), .B(KEYINPUT10), .Z(n1380) );
NAND2_X1 U1076 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
XNOR2_X1 U1077 ( .A(G104), .B(n1386), .ZN(n1389) );
NAND2_X1 U1078 ( .A1(n1390), .A2(n1391), .ZN(n1386) );
NAND2_X1 U1079 ( .A1(G122), .A2(n1392), .ZN(n1391) );
XOR2_X1 U1080 ( .A(KEYINPUT27), .B(n1393), .Z(n1390) );
NOR2_X1 U1081 ( .A1(G122), .A2(n1392), .ZN(n1393) );
INV_X1 U1082 ( .A(G113), .ZN(n1392) );
XNOR2_X1 U1083 ( .A(n1384), .B(n1385), .ZN(n1388) );
XNOR2_X1 U1084 ( .A(n1394), .B(n1395), .ZN(n1385) );
NOR2_X1 U1085 ( .A1(G131), .A2(KEYINPUT46), .ZN(n1395) );
XNOR2_X1 U1086 ( .A(G143), .B(n1396), .ZN(n1394) );
NOR2_X1 U1087 ( .A1(KEYINPUT12), .A2(n1397), .ZN(n1396) );
XNOR2_X1 U1088 ( .A(KEYINPUT29), .B(n1310), .ZN(n1397) );
XNOR2_X1 U1089 ( .A(n1398), .B(n1165), .ZN(n1384) );
XNOR2_X1 U1090 ( .A(G140), .B(n1303), .ZN(n1165) );
INV_X1 U1091 ( .A(G125), .ZN(n1303) );
NAND3_X1 U1092 ( .A1(n1365), .A2(n1089), .A3(G214), .ZN(n1398) );
XNOR2_X1 U1093 ( .A(n1144), .B(G478), .ZN(n1337) );
NOR2_X1 U1094 ( .A1(n1199), .A2(G902), .ZN(n1144) );
INV_X1 U1095 ( .A(n1197), .ZN(n1199) );
XNOR2_X1 U1096 ( .A(n1399), .B(n1400), .ZN(n1197) );
XOR2_X1 U1097 ( .A(G107), .B(n1401), .Z(n1400) );
XNOR2_X1 U1098 ( .A(G122), .B(n1402), .ZN(n1401) );
INV_X1 U1099 ( .A(G116), .ZN(n1402) );
XOR2_X1 U1100 ( .A(n1403), .B(n1404), .Z(n1399) );
NOR4_X1 U1101 ( .A1(KEYINPUT33), .A2(G953), .A3(n1405), .A4(n1406), .ZN(n1404) );
XOR2_X1 U1102 ( .A(KEYINPUT43), .B(G234), .Z(n1406) );
INV_X1 U1103 ( .A(G217), .ZN(n1405) );
NAND2_X1 U1104 ( .A1(n1407), .A2(n1408), .ZN(n1403) );
NAND2_X1 U1105 ( .A1(G134), .A2(n1169), .ZN(n1408) );
XOR2_X1 U1106 ( .A(KEYINPUT5), .B(n1409), .Z(n1407) );
NOR2_X1 U1107 ( .A1(G134), .A2(n1169), .ZN(n1409) );
XNOR2_X1 U1108 ( .A(n1378), .B(G143), .ZN(n1169) );
INV_X1 U1109 ( .A(G128), .ZN(n1378) );
XNOR2_X1 U1110 ( .A(n1123), .B(KEYINPUT52), .ZN(n1348) );
NOR2_X1 U1111 ( .A1(n1326), .A2(n1340), .ZN(n1123) );
INV_X1 U1112 ( .A(n1325), .ZN(n1340) );
NAND2_X1 U1113 ( .A1(n1410), .A2(n1411), .ZN(n1325) );
OR2_X1 U1114 ( .A1(n1136), .A2(n1135), .ZN(n1411) );
XOR2_X1 U1115 ( .A(n1138), .B(KEYINPUT6), .Z(n1410) );
NAND2_X1 U1116 ( .A1(n1135), .A2(n1136), .ZN(n1138) );
NAND2_X1 U1117 ( .A1(G217), .A2(n1349), .ZN(n1136) );
NAND2_X1 U1118 ( .A1(G234), .A2(n1204), .ZN(n1349) );
NOR2_X1 U1119 ( .A1(n1191), .A2(G902), .ZN(n1135) );
XOR2_X1 U1120 ( .A(n1412), .B(n1413), .Z(n1191) );
XOR2_X1 U1121 ( .A(n1414), .B(n1415), .Z(n1413) );
XNOR2_X1 U1122 ( .A(G110), .B(G125), .ZN(n1415) );
NAND2_X1 U1123 ( .A1(KEYINPUT47), .A2(G140), .ZN(n1414) );
XOR2_X1 U1124 ( .A(n1360), .B(n1416), .Z(n1412) );
XOR2_X1 U1125 ( .A(n1417), .B(n1418), .Z(n1416) );
NAND3_X1 U1126 ( .A1(G234), .A2(n1089), .A3(G221), .ZN(n1418) );
NAND2_X1 U1127 ( .A1(KEYINPUT34), .A2(G119), .ZN(n1417) );
XNOR2_X1 U1128 ( .A(n1419), .B(n1310), .ZN(n1360) );
XOR2_X1 U1129 ( .A(n1420), .B(n1219), .Z(n1326) );
INV_X1 U1130 ( .A(G472), .ZN(n1219) );
NAND2_X1 U1131 ( .A1(n1421), .A2(n1204), .ZN(n1420) );
INV_X1 U1132 ( .A(G902), .ZN(n1204) );
XOR2_X1 U1133 ( .A(n1422), .B(n1423), .Z(n1421) );
XOR2_X1 U1134 ( .A(n1217), .B(n1216), .Z(n1423) );
AND3_X1 U1135 ( .A1(n1365), .A2(n1089), .A3(G210), .ZN(n1216) );
INV_X1 U1136 ( .A(G953), .ZN(n1089) );
INV_X1 U1137 ( .A(G237), .ZN(n1365) );
XOR2_X1 U1138 ( .A(n1424), .B(n1425), .Z(n1217) );
XOR2_X1 U1139 ( .A(n1377), .B(n1371), .Z(n1425) );
XNOR2_X1 U1140 ( .A(n1426), .B(n1427), .ZN(n1371) );
XOR2_X1 U1141 ( .A(KEYINPUT15), .B(G119), .Z(n1427) );
XNOR2_X1 U1142 ( .A(G116), .B(G113), .ZN(n1426) );
XNOR2_X1 U1143 ( .A(n1428), .B(G143), .ZN(n1377) );
NAND2_X1 U1144 ( .A1(n1429), .A2(n1310), .ZN(n1428) );
INV_X1 U1145 ( .A(G146), .ZN(n1310) );
XNOR2_X1 U1146 ( .A(KEYINPUT40), .B(KEYINPUT37), .ZN(n1429) );
XOR2_X1 U1147 ( .A(n1419), .B(n1163), .Z(n1424) );
XOR2_X1 U1148 ( .A(G131), .B(G134), .Z(n1163) );
XNOR2_X1 U1149 ( .A(G128), .B(n1164), .ZN(n1419) );
XNOR2_X1 U1150 ( .A(n1321), .B(KEYINPUT63), .ZN(n1164) );
INV_X1 U1151 ( .A(G137), .ZN(n1321) );
XNOR2_X1 U1152 ( .A(n1430), .B(n1431), .ZN(n1422) );
INV_X1 U1153 ( .A(G101), .ZN(n1431) );
XNOR2_X1 U1154 ( .A(KEYINPUT59), .B(KEYINPUT32), .ZN(n1430) );
endmodule


