//Key = 0100000000010101111101000110001000101011010111010010011111101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425;

XNOR2_X1 U781 ( .A(G107), .B(n1076), .ZN(G9) );
NOR2_X1 U782 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR4_X1 U783 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
NOR2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U785 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR2_X1 U786 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U787 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR3_X1 U789 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1091) );
NOR2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U791 ( .A(KEYINPUT26), .B(n1098), .ZN(n1097) );
INV_X1 U792 ( .A(n1099), .ZN(n1096) );
NOR2_X1 U793 ( .A1(n1100), .A2(n1101), .ZN(n1093) );
NOR2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR3_X1 U795 ( .A1(n1101), .A2(n1104), .A3(n1098), .ZN(n1089) );
NOR2_X1 U796 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U798 ( .A1(KEYINPUT61), .A2(n1109), .ZN(n1105) );
NOR4_X1 U799 ( .A1(n1110), .A2(n1098), .A3(n1092), .A4(n1101), .ZN(n1085) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U801 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND4_X1 U802 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1079) );
NAND3_X1 U803 ( .A1(n1119), .A2(n1120), .A3(KEYINPUT61), .ZN(n1115) );
OR4_X1 U804 ( .A1(n1084), .A2(n1101), .A3(n1098), .A4(n1109), .ZN(n1120) );
INV_X1 U805 ( .A(n1121), .ZN(n1098) );
NOR3_X1 U806 ( .A1(n1122), .A2(G953), .A3(G952), .ZN(n1077) );
INV_X1 U807 ( .A(n1117), .ZN(n1122) );
NAND3_X1 U808 ( .A1(n1123), .A2(n1114), .A3(n1124), .ZN(n1117) );
NOR3_X1 U809 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
NOR2_X1 U810 ( .A1(KEYINPUT44), .A2(n1128), .ZN(n1127) );
NOR3_X1 U811 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
AND2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
AND2_X1 U813 ( .A1(n1092), .A2(KEYINPUT44), .ZN(n1126) );
XOR2_X1 U814 ( .A(n1134), .B(n1135), .Z(n1125) );
XOR2_X1 U815 ( .A(n1136), .B(KEYINPUT63), .Z(n1123) );
NAND4_X1 U816 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
NOR3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
XOR2_X1 U818 ( .A(n1144), .B(KEYINPUT34), .Z(n1143) );
NOR2_X1 U819 ( .A1(G478), .A2(n1145), .ZN(n1142) );
NAND2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(n1138) );
NAND2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
INV_X1 U823 ( .A(KEYINPUT38), .ZN(n1151) );
INV_X1 U824 ( .A(n1152), .ZN(n1148) );
NAND3_X1 U825 ( .A1(KEYINPUT38), .A2(n1150), .A3(n1153), .ZN(n1137) );
INV_X1 U826 ( .A(n1146), .ZN(n1153) );
XNOR2_X1 U827 ( .A(n1152), .B(KEYINPUT23), .ZN(n1150) );
XOR2_X1 U828 ( .A(n1154), .B(n1155), .Z(G72) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND3_X1 U830 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
XOR2_X1 U831 ( .A(KEYINPUT54), .B(n1161), .Z(n1160) );
NOR2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U833 ( .A(n1164), .B(n1165), .ZN(n1163) );
NAND2_X1 U834 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
OR2_X1 U835 ( .A1(n1118), .A2(G900), .ZN(n1159) );
NAND3_X1 U836 ( .A1(n1168), .A2(n1169), .A3(n1162), .ZN(n1158) );
NAND3_X1 U837 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1162) );
NAND2_X1 U838 ( .A1(KEYINPUT9), .A2(n1173), .ZN(n1171) );
OR2_X1 U839 ( .A1(n1174), .A2(KEYINPUT9), .ZN(n1170) );
OR2_X1 U840 ( .A1(n1166), .A2(n1165), .ZN(n1169) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1166), .ZN(n1168) );
XNOR2_X1 U842 ( .A(n1176), .B(G128), .ZN(n1166) );
XNOR2_X1 U843 ( .A(n1167), .B(n1165), .ZN(n1175) );
INV_X1 U844 ( .A(KEYINPUT42), .ZN(n1167) );
NAND2_X1 U845 ( .A1(n1177), .A2(n1118), .ZN(n1156) );
NAND2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U847 ( .A(n1116), .B(KEYINPUT35), .Z(n1178) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1181), .ZN(n1154) );
AND2_X1 U849 ( .A1(G227), .A2(G900), .ZN(n1180) );
XOR2_X1 U850 ( .A(n1182), .B(n1183), .Z(G69) );
XOR2_X1 U851 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U852 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U853 ( .A1(G953), .A2(n1188), .ZN(n1187) );
NAND2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
NAND2_X1 U855 ( .A1(G898), .A2(G224), .ZN(n1190) );
INV_X1 U856 ( .A(n1181), .ZN(n1189) );
XOR2_X1 U857 ( .A(G953), .B(KEYINPUT55), .Z(n1181) );
NOR2_X1 U858 ( .A1(n1191), .A2(G953), .ZN(n1182) );
NOR3_X1 U859 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(G66) );
NOR4_X1 U860 ( .A1(n1195), .A2(n1196), .A3(KEYINPUT48), .A4(n1152), .ZN(n1194) );
INV_X1 U861 ( .A(n1197), .ZN(n1195) );
NOR2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(n1193) );
NOR3_X1 U863 ( .A1(n1196), .A2(n1199), .A3(n1152), .ZN(n1198) );
AND2_X1 U864 ( .A1(n1200), .A2(KEYINPUT48), .ZN(n1199) );
NOR2_X1 U865 ( .A1(KEYINPUT3), .A2(n1200), .ZN(n1197) );
NOR2_X1 U866 ( .A1(n1192), .A2(n1201), .ZN(G63) );
XOR2_X1 U867 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U868 ( .A1(n1204), .A2(n1196), .ZN(n1202) );
NOR3_X1 U869 ( .A1(n1192), .A2(n1205), .A3(n1206), .ZN(G60) );
NOR3_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
XOR2_X1 U871 ( .A(KEYINPUT43), .B(n1210), .Z(n1209) );
NOR2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1208) );
INV_X1 U873 ( .A(KEYINPUT6), .ZN(n1212) );
NOR2_X1 U874 ( .A1(n1213), .A2(n1214), .ZN(n1205) );
NOR2_X1 U875 ( .A1(KEYINPUT6), .A2(n1211), .ZN(n1214) );
XOR2_X1 U876 ( .A(n1210), .B(KEYINPUT47), .Z(n1211) );
INV_X1 U877 ( .A(n1207), .ZN(n1213) );
NAND2_X1 U878 ( .A1(n1215), .A2(G475), .ZN(n1207) );
XNOR2_X1 U879 ( .A(G104), .B(n1216), .ZN(G6) );
NAND2_X1 U880 ( .A1(n1094), .A2(n1217), .ZN(n1216) );
NOR2_X1 U881 ( .A1(n1192), .A2(n1218), .ZN(G57) );
XOR2_X1 U882 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U883 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NOR2_X1 U884 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
INV_X1 U885 ( .A(n1225), .ZN(n1224) );
XNOR2_X1 U886 ( .A(KEYINPUT40), .B(n1226), .ZN(n1223) );
NOR2_X1 U887 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
NAND2_X1 U888 ( .A1(n1215), .A2(G472), .ZN(n1226) );
INV_X1 U889 ( .A(n1196), .ZN(n1215) );
XNOR2_X1 U890 ( .A(n1227), .B(n1228), .ZN(n1225) );
XOR2_X1 U891 ( .A(n1229), .B(G116), .Z(n1227) );
NAND2_X1 U892 ( .A1(KEYINPUT57), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U893 ( .A(n1231), .B(n1232), .ZN(n1219) );
NOR2_X1 U894 ( .A1(n1192), .A2(n1233), .ZN(G54) );
XOR2_X1 U895 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U896 ( .A(n1236), .B(n1237), .Z(n1235) );
NOR2_X1 U897 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U898 ( .A1(KEYINPUT25), .A2(n1165), .ZN(n1239) );
NOR2_X1 U899 ( .A1(KEYINPUT51), .A2(n1240), .ZN(n1238) );
XNOR2_X1 U900 ( .A(n1241), .B(n1242), .ZN(n1234) );
NOR2_X1 U901 ( .A1(n1129), .A2(n1196), .ZN(n1242) );
NOR2_X1 U902 ( .A1(n1192), .A2(n1243), .ZN(G51) );
XOR2_X1 U903 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U904 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U905 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U906 ( .A(n1173), .B(G116), .ZN(n1249) );
XOR2_X1 U907 ( .A(KEYINPUT5), .B(KEYINPUT41), .Z(n1248) );
XOR2_X1 U908 ( .A(n1250), .B(n1251), .Z(n1246) );
XOR2_X1 U909 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U910 ( .A1(n1135), .A2(n1196), .ZN(n1253) );
NAND2_X1 U911 ( .A1(n1254), .A2(n1255), .ZN(n1196) );
NAND3_X1 U912 ( .A1(n1179), .A2(n1116), .A3(n1191), .ZN(n1255) );
INV_X1 U913 ( .A(n1080), .ZN(n1191) );
NAND4_X1 U914 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1080) );
NOR4_X1 U915 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1259) );
INV_X1 U916 ( .A(n1264), .ZN(n1263) );
NOR2_X1 U917 ( .A1(n1265), .A2(n1266), .ZN(n1258) );
NOR3_X1 U918 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1266) );
NAND3_X1 U919 ( .A1(n1270), .A2(n1109), .A3(n1112), .ZN(n1267) );
INV_X1 U920 ( .A(n1076), .ZN(n1265) );
NAND3_X1 U921 ( .A1(n1121), .A2(n1217), .A3(n1099), .ZN(n1076) );
NAND3_X1 U922 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1257) );
OR2_X1 U923 ( .A1(n1274), .A2(KEYINPUT7), .ZN(n1272) );
NAND2_X1 U924 ( .A1(KEYINPUT7), .A2(n1275), .ZN(n1271) );
NAND3_X1 U925 ( .A1(n1276), .A2(n1270), .A3(n1277), .ZN(n1275) );
NAND2_X1 U926 ( .A1(n1217), .A2(n1278), .ZN(n1256) );
NAND2_X1 U927 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U928 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U929 ( .A(KEYINPUT49), .B(n1103), .Z(n1282) );
NAND2_X1 U930 ( .A1(n1094), .A2(n1269), .ZN(n1279) );
INV_X1 U931 ( .A(KEYINPUT10), .ZN(n1269) );
INV_X1 U932 ( .A(n1268), .ZN(n1094) );
NAND2_X1 U933 ( .A1(n1283), .A2(n1121), .ZN(n1268) );
INV_X1 U934 ( .A(n1082), .ZN(n1179) );
NAND4_X1 U935 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1082) );
NOR4_X1 U936 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(n1287) );
NOR2_X1 U937 ( .A1(n1292), .A2(n1293), .ZN(n1286) );
INV_X1 U938 ( .A(n1294), .ZN(n1292) );
NAND3_X1 U939 ( .A1(n1295), .A2(n1276), .A3(n1296), .ZN(n1285) );
INV_X1 U940 ( .A(KEYINPUT53), .ZN(n1296) );
NAND2_X1 U941 ( .A1(n1297), .A2(KEYINPUT53), .ZN(n1284) );
XNOR2_X1 U942 ( .A(G902), .B(KEYINPUT30), .ZN(n1254) );
XNOR2_X1 U943 ( .A(n1298), .B(n1299), .ZN(n1250) );
NOR2_X1 U944 ( .A1(n1118), .A2(G952), .ZN(n1192) );
XNOR2_X1 U945 ( .A(n1300), .B(n1293), .ZN(G48) );
AND2_X1 U946 ( .A1(n1301), .A2(n1283), .ZN(n1293) );
XNOR2_X1 U947 ( .A(n1302), .B(n1297), .ZN(G45) );
AND2_X1 U948 ( .A1(n1295), .A2(n1112), .ZN(n1297) );
AND4_X1 U949 ( .A1(n1102), .A2(n1303), .A3(n1141), .A4(n1304), .ZN(n1295) );
XNOR2_X1 U950 ( .A(G140), .B(n1294), .ZN(G42) );
NAND3_X1 U951 ( .A1(n1283), .A2(n1305), .A3(n1103), .ZN(n1294) );
XNOR2_X1 U952 ( .A(n1306), .B(n1291), .ZN(G39) );
AND2_X1 U953 ( .A1(n1273), .A2(n1305), .ZN(n1291) );
XOR2_X1 U954 ( .A(n1290), .B(n1307), .Z(G36) );
NOR2_X1 U955 ( .A1(KEYINPUT37), .A2(n1308), .ZN(n1307) );
INV_X1 U956 ( .A(G134), .ZN(n1308) );
AND3_X1 U957 ( .A1(n1305), .A2(n1099), .A3(n1102), .ZN(n1290) );
XNOR2_X1 U958 ( .A(G131), .B(n1116), .ZN(G33) );
NAND3_X1 U959 ( .A1(n1283), .A2(n1305), .A3(n1102), .ZN(n1116) );
AND2_X1 U960 ( .A1(n1303), .A2(n1119), .ZN(n1305) );
INV_X1 U961 ( .A(n1088), .ZN(n1119) );
NAND2_X1 U962 ( .A1(n1309), .A2(n1114), .ZN(n1088) );
INV_X1 U963 ( .A(n1113), .ZN(n1309) );
XOR2_X1 U964 ( .A(G128), .B(n1289), .Z(G30) );
AND2_X1 U965 ( .A1(n1301), .A2(n1099), .ZN(n1289) );
AND4_X1 U966 ( .A1(n1303), .A2(n1112), .A3(n1310), .A4(n1311), .ZN(n1301) );
INV_X1 U967 ( .A(n1276), .ZN(n1112) );
NOR2_X1 U968 ( .A1(n1109), .A2(n1312), .ZN(n1303) );
XNOR2_X1 U969 ( .A(G101), .B(n1264), .ZN(G3) );
NAND3_X1 U970 ( .A1(n1102), .A2(n1217), .A3(n1281), .ZN(n1264) );
XNOR2_X1 U971 ( .A(n1288), .B(n1313), .ZN(G27) );
NAND2_X1 U972 ( .A1(KEYINPUT36), .A2(G125), .ZN(n1313) );
AND4_X1 U973 ( .A1(n1103), .A2(n1277), .A3(n1314), .A4(n1283), .ZN(n1288) );
NOR2_X1 U974 ( .A1(n1312), .A2(n1276), .ZN(n1314) );
AND2_X1 U975 ( .A1(n1315), .A2(n1084), .ZN(n1312) );
NAND4_X1 U976 ( .A1(G902), .A2(G953), .A3(n1316), .A4(n1317), .ZN(n1315) );
XOR2_X1 U977 ( .A(KEYINPUT58), .B(G900), .Z(n1316) );
XOR2_X1 U978 ( .A(G122), .B(n1262), .Z(G24) );
AND4_X1 U979 ( .A1(n1274), .A2(n1121), .A3(n1141), .A4(n1304), .ZN(n1262) );
NOR2_X1 U980 ( .A1(n1311), .A2(n1310), .ZN(n1121) );
XNOR2_X1 U981 ( .A(n1318), .B(n1319), .ZN(G21) );
AND2_X1 U982 ( .A1(n1274), .A2(n1273), .ZN(n1319) );
AND3_X1 U983 ( .A1(n1310), .A2(n1311), .A3(n1281), .ZN(n1273) );
XOR2_X1 U984 ( .A(G116), .B(n1261), .Z(G18) );
AND3_X1 U985 ( .A1(n1102), .A2(n1099), .A3(n1274), .ZN(n1261) );
NOR2_X1 U986 ( .A1(n1141), .A2(n1320), .ZN(n1099) );
XOR2_X1 U987 ( .A(G113), .B(n1260), .Z(G15) );
AND3_X1 U988 ( .A1(n1102), .A2(n1283), .A3(n1274), .ZN(n1260) );
NOR3_X1 U989 ( .A1(n1276), .A2(n1321), .A3(n1092), .ZN(n1274) );
INV_X1 U990 ( .A(n1277), .ZN(n1092) );
NOR2_X1 U991 ( .A1(n1107), .A2(n1130), .ZN(n1277) );
INV_X1 U992 ( .A(n1108), .ZN(n1130) );
AND2_X1 U993 ( .A1(n1320), .A2(n1141), .ZN(n1283) );
INV_X1 U994 ( .A(n1304), .ZN(n1320) );
NOR2_X1 U995 ( .A1(n1310), .A2(n1139), .ZN(n1102) );
XNOR2_X1 U996 ( .A(G110), .B(n1322), .ZN(G12) );
NAND3_X1 U997 ( .A1(n1217), .A2(n1323), .A3(n1103), .ZN(n1322) );
AND2_X1 U998 ( .A1(n1139), .A2(n1310), .ZN(n1103) );
XNOR2_X1 U999 ( .A(n1146), .B(n1152), .ZN(n1310) );
NAND2_X1 U1000 ( .A1(G217), .A2(n1324), .ZN(n1152) );
NOR2_X1 U1001 ( .A1(n1200), .A2(G902), .ZN(n1146) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1200) );
XOR2_X1 U1003 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1004 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1005 ( .A1(G128), .A2(n1318), .ZN(n1330) );
XOR2_X1 U1006 ( .A(KEYINPUT16), .B(n1331), .Z(n1329) );
NOR2_X1 U1007 ( .A1(G128), .A2(n1318), .ZN(n1331) );
NAND2_X1 U1008 ( .A1(KEYINPUT11), .A2(n1306), .ZN(n1327) );
XOR2_X1 U1009 ( .A(n1332), .B(n1333), .Z(n1325) );
NOR2_X1 U1010 ( .A1(KEYINPUT52), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1011 ( .A(G146), .B(n1335), .ZN(n1334) );
NAND2_X1 U1012 ( .A1(n1336), .A2(n1172), .ZN(n1335) );
XOR2_X1 U1013 ( .A(n1174), .B(KEYINPUT2), .Z(n1336) );
XOR2_X1 U1014 ( .A(n1337), .B(G110), .Z(n1332) );
NAND3_X1 U1015 ( .A1(G234), .A2(n1118), .A3(G221), .ZN(n1337) );
INV_X1 U1016 ( .A(n1311), .ZN(n1139) );
XNOR2_X1 U1017 ( .A(n1338), .B(G472), .ZN(n1311) );
NAND2_X1 U1018 ( .A1(n1339), .A2(n1132), .ZN(n1338) );
XOR2_X1 U1019 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1020 ( .A(n1342), .B(n1228), .Z(n1341) );
XOR2_X1 U1021 ( .A(G113), .B(n1343), .Z(n1228) );
XNOR2_X1 U1022 ( .A(KEYINPUT27), .B(n1318), .ZN(n1343) );
XOR2_X1 U1023 ( .A(n1231), .B(n1344), .Z(n1340) );
XNOR2_X1 U1024 ( .A(n1345), .B(KEYINPUT18), .ZN(n1344) );
NAND2_X1 U1025 ( .A1(KEYINPUT17), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1026 ( .A(KEYINPUT29), .B(n1230), .ZN(n1346) );
XNOR2_X1 U1027 ( .A(n1347), .B(n1165), .ZN(n1230) );
NAND3_X1 U1028 ( .A1(n1348), .A2(n1118), .A3(G210), .ZN(n1231) );
XNOR2_X1 U1029 ( .A(KEYINPUT20), .B(n1101), .ZN(n1323) );
INV_X1 U1030 ( .A(n1281), .ZN(n1101) );
NOR2_X1 U1031 ( .A1(n1304), .A2(n1141), .ZN(n1281) );
XNOR2_X1 U1032 ( .A(n1349), .B(G475), .ZN(n1141) );
NAND2_X1 U1033 ( .A1(n1210), .A2(n1132), .ZN(n1349) );
XNOR2_X1 U1034 ( .A(n1350), .B(n1351), .ZN(n1210) );
XNOR2_X1 U1035 ( .A(n1300), .B(n1352), .ZN(n1351) );
NOR2_X1 U1036 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1037 ( .A(n1355), .B(KEYINPUT1), .Z(n1354) );
NAND2_X1 U1038 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NOR2_X1 U1039 ( .A1(n1356), .A2(n1357), .ZN(n1353) );
XNOR2_X1 U1040 ( .A(KEYINPUT39), .B(n1358), .ZN(n1357) );
INV_X1 U1041 ( .A(G131), .ZN(n1358) );
XOR2_X1 U1042 ( .A(n1359), .B(n1360), .Z(n1356) );
NOR2_X1 U1043 ( .A1(G143), .A2(KEYINPUT12), .ZN(n1360) );
NAND3_X1 U1044 ( .A1(n1348), .A2(n1118), .A3(G214), .ZN(n1359) );
XNOR2_X1 U1045 ( .A(n1361), .B(KEYINPUT21), .ZN(n1348) );
XOR2_X1 U1046 ( .A(n1362), .B(n1363), .Z(n1350) );
NAND2_X1 U1047 ( .A1(n1364), .A2(n1174), .ZN(n1362) );
NAND2_X1 U1048 ( .A1(G125), .A2(n1365), .ZN(n1174) );
XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n1172), .ZN(n1364) );
NAND2_X1 U1050 ( .A1(G140), .A2(n1173), .ZN(n1172) );
NAND2_X1 U1051 ( .A1(n1366), .A2(n1144), .ZN(n1304) );
NAND2_X1 U1052 ( .A1(G478), .A2(n1145), .ZN(n1144) );
INV_X1 U1053 ( .A(n1367), .ZN(n1145) );
NAND2_X1 U1054 ( .A1(n1367), .A2(n1204), .ZN(n1366) );
INV_X1 U1055 ( .A(G478), .ZN(n1204) );
NOR2_X1 U1056 ( .A1(n1203), .A2(G902), .ZN(n1367) );
XNOR2_X1 U1057 ( .A(n1368), .B(n1369), .ZN(n1203) );
NOR2_X1 U1058 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1059 ( .A(KEYINPUT31), .B(n1372), .Z(n1371) );
NOR2_X1 U1060 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
AND2_X1 U1061 ( .A1(n1374), .A2(n1373), .ZN(n1370) );
AND2_X1 U1062 ( .A1(n1375), .A2(n1376), .ZN(n1373) );
NAND2_X1 U1063 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
XNOR2_X1 U1064 ( .A(G107), .B(KEYINPUT14), .ZN(n1378) );
XNOR2_X1 U1065 ( .A(G122), .B(G116), .ZN(n1377) );
NAND2_X1 U1066 ( .A1(n1379), .A2(n1380), .ZN(n1375) );
XNOR2_X1 U1067 ( .A(KEYINPUT4), .B(n1381), .ZN(n1380) );
XOR2_X1 U1068 ( .A(G122), .B(G116), .Z(n1379) );
NAND2_X1 U1069 ( .A1(n1382), .A2(n1383), .ZN(n1374) );
NAND2_X1 U1070 ( .A1(G134), .A2(n1384), .ZN(n1383) );
XOR2_X1 U1071 ( .A(KEYINPUT15), .B(n1385), .Z(n1382) );
NOR2_X1 U1072 ( .A1(G134), .A2(n1384), .ZN(n1385) );
NAND2_X1 U1073 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
NAND2_X1 U1074 ( .A1(G128), .A2(n1302), .ZN(n1387) );
XOR2_X1 U1075 ( .A(KEYINPUT56), .B(n1388), .Z(n1386) );
NOR2_X1 U1076 ( .A1(G128), .A2(n1302), .ZN(n1388) );
NAND3_X1 U1077 ( .A1(G217), .A2(n1118), .A3(G234), .ZN(n1368) );
NOR3_X1 U1078 ( .A1(n1276), .A2(n1321), .A3(n1109), .ZN(n1217) );
NAND2_X1 U1079 ( .A1(n1107), .A2(n1108), .ZN(n1109) );
NAND2_X1 U1080 ( .A1(G221), .A2(n1324), .ZN(n1108) );
NAND2_X1 U1081 ( .A1(G234), .A2(n1132), .ZN(n1324) );
XOR2_X1 U1082 ( .A(n1389), .B(n1129), .Z(n1107) );
INV_X1 U1083 ( .A(G469), .ZN(n1129) );
NAND2_X1 U1084 ( .A1(n1133), .A2(n1132), .ZN(n1389) );
XNOR2_X1 U1085 ( .A(n1390), .B(n1391), .ZN(n1133) );
XOR2_X1 U1086 ( .A(KEYINPUT24), .B(n1392), .Z(n1391) );
NOR2_X1 U1087 ( .A1(KEYINPUT32), .A2(n1240), .ZN(n1392) );
INV_X1 U1088 ( .A(n1165), .ZN(n1240) );
XOR2_X1 U1089 ( .A(G131), .B(n1393), .Z(n1165) );
XNOR2_X1 U1090 ( .A(n1306), .B(G134), .ZN(n1393) );
INV_X1 U1091 ( .A(G137), .ZN(n1306) );
XNOR2_X1 U1092 ( .A(n1236), .B(n1394), .ZN(n1390) );
INV_X1 U1093 ( .A(n1241), .ZN(n1394) );
XNOR2_X1 U1094 ( .A(n1395), .B(n1396), .ZN(n1241) );
XNOR2_X1 U1095 ( .A(n1365), .B(G110), .ZN(n1396) );
INV_X1 U1096 ( .A(G140), .ZN(n1365) );
NAND2_X1 U1097 ( .A1(G227), .A2(n1118), .ZN(n1395) );
XOR2_X1 U1098 ( .A(n1298), .B(n1397), .Z(n1236) );
XOR2_X1 U1099 ( .A(n1398), .B(n1176), .Z(n1397) );
XNOR2_X1 U1100 ( .A(KEYINPUT45), .B(n1399), .ZN(n1176) );
NOR2_X1 U1101 ( .A1(KEYINPUT28), .A2(n1299), .ZN(n1399) );
NAND3_X1 U1102 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1398) );
OR2_X1 U1103 ( .A1(n1381), .A2(KEYINPUT19), .ZN(n1402) );
NAND3_X1 U1104 ( .A1(KEYINPUT19), .A2(n1381), .A3(G104), .ZN(n1401) );
NAND2_X1 U1105 ( .A1(n1403), .A2(n1404), .ZN(n1400) );
INV_X1 U1106 ( .A(G104), .ZN(n1404) );
NAND2_X1 U1107 ( .A1(n1405), .A2(KEYINPUT19), .ZN(n1403) );
XNOR2_X1 U1108 ( .A(G107), .B(KEYINPUT46), .ZN(n1405) );
XNOR2_X1 U1109 ( .A(G101), .B(G128), .ZN(n1298) );
INV_X1 U1110 ( .A(n1270), .ZN(n1321) );
NAND2_X1 U1111 ( .A1(n1084), .A2(n1406), .ZN(n1270) );
NAND4_X1 U1112 ( .A1(n1407), .A2(G902), .A3(n1317), .A4(n1188), .ZN(n1406) );
INV_X1 U1113 ( .A(G898), .ZN(n1188) );
XNOR2_X1 U1114 ( .A(G953), .B(KEYINPUT13), .ZN(n1407) );
NAND3_X1 U1115 ( .A1(n1317), .A2(n1118), .A3(G952), .ZN(n1084) );
NAND2_X1 U1116 ( .A1(G237), .A2(G234), .ZN(n1317) );
NAND2_X1 U1117 ( .A1(n1113), .A2(n1114), .ZN(n1276) );
NAND2_X1 U1118 ( .A1(G214), .A2(n1408), .ZN(n1114) );
XNOR2_X1 U1119 ( .A(n1135), .B(n1409), .ZN(n1113) );
NOR2_X1 U1120 ( .A1(KEYINPUT0), .A2(n1134), .ZN(n1409) );
NAND2_X1 U1121 ( .A1(n1410), .A2(n1132), .ZN(n1134) );
XOR2_X1 U1122 ( .A(n1411), .B(n1186), .Z(n1410) );
XOR2_X1 U1123 ( .A(n1244), .B(n1342), .Z(n1186) );
XNOR2_X1 U1124 ( .A(n1232), .B(G116), .ZN(n1342) );
INV_X1 U1125 ( .A(G101), .ZN(n1232) );
XOR2_X1 U1126 ( .A(n1412), .B(n1413), .Z(n1244) );
XNOR2_X1 U1127 ( .A(n1381), .B(n1414), .ZN(n1413) );
XOR2_X1 U1128 ( .A(KEYINPUT33), .B(G110), .Z(n1414) );
INV_X1 U1129 ( .A(G107), .ZN(n1381) );
XNOR2_X1 U1130 ( .A(n1363), .B(n1415), .ZN(n1412) );
NOR2_X1 U1131 ( .A1(KEYINPUT62), .A2(n1416), .ZN(n1415) );
XNOR2_X1 U1132 ( .A(KEYINPUT50), .B(n1318), .ZN(n1416) );
INV_X1 U1133 ( .A(G119), .ZN(n1318) );
XOR2_X1 U1134 ( .A(G104), .B(n1417), .Z(n1363) );
XOR2_X1 U1135 ( .A(G122), .B(G113), .Z(n1417) );
NAND3_X1 U1136 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n1411) );
NAND2_X1 U1137 ( .A1(n1421), .A2(n1422), .ZN(n1420) );
NAND2_X1 U1138 ( .A1(n1252), .A2(n1423), .ZN(n1422) );
XNOR2_X1 U1139 ( .A(n1347), .B(G125), .ZN(n1421) );
OR2_X1 U1140 ( .A1(n1424), .A2(n1252), .ZN(n1419) );
NAND4_X1 U1141 ( .A1(n1424), .A2(n1423), .A3(n1425), .A4(n1252), .ZN(n1418) );
AND2_X1 U1142 ( .A1(G224), .A2(n1118), .ZN(n1252) );
INV_X1 U1143 ( .A(G953), .ZN(n1118) );
XNOR2_X1 U1144 ( .A(n1173), .B(n1347), .ZN(n1425) );
XNOR2_X1 U1145 ( .A(G128), .B(n1299), .ZN(n1347) );
XNOR2_X1 U1146 ( .A(n1302), .B(n1300), .ZN(n1299) );
INV_X1 U1147 ( .A(G146), .ZN(n1300) );
INV_X1 U1148 ( .A(G143), .ZN(n1302) );
INV_X1 U1149 ( .A(G125), .ZN(n1173) );
INV_X1 U1150 ( .A(KEYINPUT59), .ZN(n1423) );
XNOR2_X1 U1151 ( .A(KEYINPUT8), .B(KEYINPUT22), .ZN(n1424) );
NAND2_X1 U1152 ( .A1(G210), .A2(n1408), .ZN(n1135) );
NAND2_X1 U1153 ( .A1(n1361), .A2(n1132), .ZN(n1408) );
INV_X1 U1154 ( .A(G902), .ZN(n1132) );
INV_X1 U1155 ( .A(G237), .ZN(n1361) );
endmodule


