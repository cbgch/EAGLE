//Key = 0100101000110110100100010011001110110011111111110010110111011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405;

XOR2_X1 U768 ( .A(n1073), .B(n1074), .Z(G9) );
NAND2_X1 U769 ( .A1(KEYINPUT6), .A2(n1075), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(G75) );
NOR3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NAND3_X1 U772 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND3_X1 U775 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND2_X1 U777 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
OR2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U779 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
XNOR2_X1 U780 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND3_X1 U781 ( .A1(n1093), .A2(n1101), .A3(n1097), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U783 ( .A1(n1090), .A2(n1104), .ZN(n1103) );
OR2_X1 U784 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U785 ( .A1(n1088), .A2(n1107), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U787 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR3_X1 U788 ( .A1(n1112), .A2(G953), .A3(n1113), .ZN(n1076) );
INV_X1 U789 ( .A(n1081), .ZN(n1113) );
NAND4_X1 U790 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1081) );
NOR4_X1 U791 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1117) );
XOR2_X1 U792 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U793 ( .A(G475), .B(n1124), .ZN(n1120) );
NOR3_X1 U794 ( .A1(n1125), .A2(n1110), .A3(n1099), .ZN(n1116) );
NOR2_X1 U795 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR2_X1 U796 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U797 ( .A1(KEYINPUT53), .A2(n1130), .ZN(n1128) );
NAND3_X1 U798 ( .A1(n1131), .A2(n1132), .A3(KEYINPUT53), .ZN(n1115) );
NAND2_X1 U799 ( .A1(G469), .A2(n1130), .ZN(n1132) );
INV_X1 U800 ( .A(KEYINPUT4), .ZN(n1130) );
NAND2_X1 U801 ( .A1(KEYINPUT4), .A2(n1133), .ZN(n1131) );
NAND2_X1 U802 ( .A1(G469), .A2(n1127), .ZN(n1133) );
XOR2_X1 U803 ( .A(n1134), .B(n1135), .Z(n1114) );
XNOR2_X1 U804 ( .A(G472), .B(KEYINPUT13), .ZN(n1135) );
XNOR2_X1 U805 ( .A(KEYINPUT17), .B(n1079), .ZN(n1112) );
XOR2_X1 U806 ( .A(n1136), .B(n1137), .Z(G72) );
XOR2_X1 U807 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U808 ( .A1(G953), .A2(n1140), .ZN(n1139) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1140) );
NAND2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND2_X1 U811 ( .A1(G953), .A2(n1143), .ZN(n1142) );
XOR2_X1 U812 ( .A(n1144), .B(n1145), .Z(n1141) );
NAND2_X1 U813 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NAND2_X1 U814 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U815 ( .A(n1150), .B(KEYINPUT0), .Z(n1146) );
OR2_X1 U816 ( .A1(n1149), .A2(n1148), .ZN(n1150) );
XOR2_X1 U817 ( .A(n1151), .B(n1152), .Z(n1148) );
NOR2_X1 U818 ( .A1(G137), .A2(KEYINPUT22), .ZN(n1152) );
XNOR2_X1 U819 ( .A(G131), .B(G134), .ZN(n1151) );
AND2_X1 U820 ( .A1(n1153), .A2(n1082), .ZN(n1136) );
NAND3_X1 U821 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(G69) );
NAND2_X1 U822 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
OR2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U826 ( .A1(KEYINPUT7), .A2(n1164), .ZN(n1163) );
NAND2_X1 U827 ( .A1(n1159), .A2(n1165), .ZN(n1164) );
NAND3_X1 U828 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1162) );
INV_X1 U829 ( .A(KEYINPUT7), .ZN(n1168) );
NAND2_X1 U830 ( .A1(n1157), .A2(n1159), .ZN(n1166) );
XNOR2_X1 U831 ( .A(n1167), .B(KEYINPUT47), .ZN(n1159) );
NAND2_X1 U832 ( .A1(n1169), .A2(G953), .ZN(n1167) );
XOR2_X1 U833 ( .A(n1170), .B(KEYINPUT37), .Z(n1169) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1170) );
INV_X1 U835 ( .A(n1165), .ZN(n1157) );
NAND2_X1 U836 ( .A1(n1082), .A2(n1171), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1158), .A2(n1172), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1082), .A2(G898), .ZN(n1172) );
XNOR2_X1 U839 ( .A(n1173), .B(n1174), .ZN(n1158) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR3_X1 U841 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(G66) );
NOR3_X1 U842 ( .A1(n1180), .A2(n1082), .A3(n1079), .ZN(n1179) );
INV_X1 U843 ( .A(G952), .ZN(n1079) );
AND2_X1 U844 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
INV_X1 U845 ( .A(KEYINPUT5), .ZN(n1180) );
XNOR2_X1 U846 ( .A(n1182), .B(n1183), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1186), .ZN(G63) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U850 ( .A1(n1189), .A2(n1185), .ZN(n1188) );
NAND2_X1 U851 ( .A1(KEYINPUT52), .A2(n1190), .ZN(n1187) );
NOR2_X1 U852 ( .A1(n1181), .A2(n1191), .ZN(G60) );
NOR3_X1 U853 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NOR3_X1 U854 ( .A1(n1195), .A2(n1196), .A3(n1185), .ZN(n1194) );
NOR2_X1 U855 ( .A1(n1197), .A2(n1198), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1199), .A2(n1196), .ZN(n1197) );
XNOR2_X1 U857 ( .A(n1200), .B(n1201), .ZN(G6) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U859 ( .A1(KEYINPUT62), .A2(n1204), .ZN(n1203) );
INV_X1 U860 ( .A(n1205), .ZN(n1204) );
NOR2_X1 U861 ( .A1(KEYINPUT26), .A2(n1205), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1206), .A2(n1207), .ZN(G57) );
XOR2_X1 U863 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U864 ( .A(n1210), .B(n1211), .ZN(n1209) );
NOR2_X1 U865 ( .A1(KEYINPUT36), .A2(n1212), .ZN(n1210) );
NOR3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
NOR2_X1 U867 ( .A1(KEYINPUT35), .A2(n1216), .ZN(n1215) );
NOR2_X1 U868 ( .A1(n1199), .A2(G902), .ZN(n1216) );
AND2_X1 U869 ( .A1(n1185), .A2(KEYINPUT35), .ZN(n1214) );
INV_X1 U870 ( .A(G472), .ZN(n1213) );
XNOR2_X1 U871 ( .A(n1217), .B(n1218), .ZN(n1208) );
NOR2_X1 U872 ( .A1(n1219), .A2(n1082), .ZN(n1206) );
XNOR2_X1 U873 ( .A(G952), .B(KEYINPUT43), .ZN(n1219) );
NOR2_X1 U874 ( .A1(n1181), .A2(n1220), .ZN(G54) );
XOR2_X1 U875 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U876 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U877 ( .A(n1225), .B(n1226), .Z(n1221) );
NOR2_X1 U878 ( .A1(n1129), .A2(n1185), .ZN(n1226) );
XNOR2_X1 U879 ( .A(KEYINPUT48), .B(n1227), .ZN(n1225) );
NOR2_X1 U880 ( .A1(KEYINPUT25), .A2(n1228), .ZN(n1227) );
NOR2_X1 U881 ( .A1(n1181), .A2(n1229), .ZN(G51) );
XOR2_X1 U882 ( .A(n1230), .B(n1231), .Z(n1229) );
XOR2_X1 U883 ( .A(n1232), .B(n1233), .Z(n1230) );
NOR2_X1 U884 ( .A1(n1123), .A2(n1185), .ZN(n1233) );
NAND2_X1 U885 ( .A1(G902), .A2(n1080), .ZN(n1185) );
INV_X1 U886 ( .A(n1199), .ZN(n1080) );
NOR2_X1 U887 ( .A1(n1153), .A2(n1171), .ZN(n1199) );
NAND4_X1 U888 ( .A1(n1205), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1171) );
NOR4_X1 U889 ( .A1(n1237), .A2(n1238), .A3(n1074), .A4(n1239), .ZN(n1236) );
INV_X1 U890 ( .A(n1240), .ZN(n1239) );
AND3_X1 U891 ( .A1(n1095), .A2(n1088), .A3(n1241), .ZN(n1074) );
NAND2_X1 U892 ( .A1(n1242), .A2(n1243), .ZN(n1235) );
NAND2_X1 U893 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NAND4_X1 U894 ( .A1(n1105), .A2(n1093), .A3(n1095), .A4(n1246), .ZN(n1245) );
XNOR2_X1 U895 ( .A(KEYINPUT27), .B(n1247), .ZN(n1246) );
NAND3_X1 U896 ( .A1(n1241), .A2(n1088), .A3(n1096), .ZN(n1205) );
NAND4_X1 U897 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1153) );
AND4_X1 U898 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1251) );
NAND2_X1 U899 ( .A1(n1256), .A2(n1257), .ZN(n1250) );
NAND2_X1 U900 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U901 ( .A1(n1097), .A2(n1090), .ZN(n1259) );
NAND2_X1 U902 ( .A1(n1095), .A2(n1242), .ZN(n1258) );
NAND2_X1 U903 ( .A1(KEYINPUT31), .A2(n1260), .ZN(n1232) );
INV_X1 U904 ( .A(n1261), .ZN(n1260) );
NOR2_X1 U905 ( .A1(n1082), .A2(G952), .ZN(n1181) );
XNOR2_X1 U906 ( .A(G146), .B(n1248), .ZN(G48) );
NAND2_X1 U907 ( .A1(n1256), .A2(n1262), .ZN(n1248) );
XNOR2_X1 U908 ( .A(G143), .B(n1249), .ZN(G45) );
NAND4_X1 U909 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1242), .ZN(n1249) );
XNOR2_X1 U910 ( .A(G140), .B(n1255), .ZN(G42) );
NAND4_X1 U911 ( .A1(n1090), .A2(n1266), .A3(n1106), .A4(n1096), .ZN(n1255) );
NAND2_X1 U912 ( .A1(n1267), .A2(n1268), .ZN(G39) );
NAND2_X1 U913 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U914 ( .A(KEYINPUT50), .B(n1271), .Z(n1267) );
NOR2_X1 U915 ( .A1(n1269), .A2(n1270), .ZN(n1271) );
NAND2_X1 U916 ( .A1(n1090), .A2(n1272), .ZN(n1270) );
XOR2_X1 U917 ( .A(KEYINPUT18), .B(n1273), .Z(n1272) );
NOR3_X1 U918 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NOR2_X1 U919 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U920 ( .A(KEYINPUT21), .ZN(n1278) );
NOR2_X1 U921 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
NOR2_X1 U922 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NOR2_X1 U923 ( .A1(KEYINPUT21), .A2(n1256), .ZN(n1275) );
INV_X1 U924 ( .A(n1097), .ZN(n1274) );
XNOR2_X1 U925 ( .A(KEYINPUT16), .B(G137), .ZN(n1269) );
XNOR2_X1 U926 ( .A(G134), .B(n1254), .ZN(G36) );
NAND3_X1 U927 ( .A1(n1264), .A2(n1095), .A3(n1090), .ZN(n1254) );
XNOR2_X1 U928 ( .A(G131), .B(n1253), .ZN(G33) );
NAND3_X1 U929 ( .A1(n1264), .A2(n1096), .A3(n1090), .ZN(n1253) );
AND2_X1 U930 ( .A1(n1111), .A2(n1283), .ZN(n1090) );
AND2_X1 U931 ( .A1(n1105), .A2(n1266), .ZN(n1264) );
INV_X1 U932 ( .A(n1280), .ZN(n1266) );
XNOR2_X1 U933 ( .A(G128), .B(n1284), .ZN(G30) );
NAND3_X1 U934 ( .A1(n1256), .A2(n1095), .A3(n1285), .ZN(n1284) );
XNOR2_X1 U935 ( .A(n1242), .B(KEYINPUT44), .ZN(n1285) );
NOR3_X1 U936 ( .A1(n1282), .A2(n1281), .A3(n1280), .ZN(n1256) );
NAND3_X1 U937 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1280) );
XNOR2_X1 U938 ( .A(G101), .B(n1234), .ZN(G3) );
NAND3_X1 U939 ( .A1(n1105), .A2(n1241), .A3(n1097), .ZN(n1234) );
XNOR2_X1 U940 ( .A(G125), .B(n1252), .ZN(G27) );
NAND4_X1 U941 ( .A1(n1093), .A2(n1262), .A3(n1106), .A4(n1286), .ZN(n1252) );
NAND2_X1 U942 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
NAND2_X1 U943 ( .A1(n1291), .A2(n1143), .ZN(n1290) );
INV_X1 U944 ( .A(G900), .ZN(n1143) );
NAND2_X1 U945 ( .A1(n1292), .A2(n1293), .ZN(G24) );
NAND2_X1 U946 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U947 ( .A(KEYINPUT32), .B(n1296), .Z(n1292) );
NOR2_X1 U948 ( .A1(n1294), .A2(n1295), .ZN(n1296) );
INV_X1 U949 ( .A(G122), .ZN(n1295) );
AND2_X1 U950 ( .A1(n1242), .A2(n1297), .ZN(n1294) );
XNOR2_X1 U951 ( .A(KEYINPUT51), .B(n1244), .ZN(n1297) );
NAND4_X1 U952 ( .A1(n1265), .A2(n1247), .A3(n1088), .A4(n1298), .ZN(n1244) );
AND2_X1 U953 ( .A1(n1093), .A2(n1263), .ZN(n1298) );
NOR2_X1 U954 ( .A1(n1299), .A2(n1118), .ZN(n1088) );
XOR2_X1 U955 ( .A(G119), .B(n1238), .Z(G21) );
AND4_X1 U956 ( .A1(n1093), .A2(n1242), .A3(n1097), .A4(n1300), .ZN(n1238) );
NOR3_X1 U957 ( .A1(n1282), .A2(n1301), .A3(n1281), .ZN(n1300) );
XNOR2_X1 U958 ( .A(G116), .B(n1302), .ZN(G18) );
NAND3_X1 U959 ( .A1(KEYINPUT1), .A2(n1242), .A3(n1303), .ZN(n1302) );
XOR2_X1 U960 ( .A(n1304), .B(KEYINPUT10), .Z(n1303) );
NAND2_X1 U961 ( .A1(n1305), .A2(n1095), .ZN(n1304) );
AND2_X1 U962 ( .A1(n1306), .A2(n1307), .ZN(n1095) );
XOR2_X1 U963 ( .A(n1265), .B(KEYINPUT8), .Z(n1306) );
XNOR2_X1 U964 ( .A(n1119), .B(KEYINPUT34), .ZN(n1265) );
XNOR2_X1 U965 ( .A(G113), .B(n1240), .ZN(G15) );
NAND2_X1 U966 ( .A1(n1305), .A2(n1262), .ZN(n1240) );
AND2_X1 U967 ( .A1(n1096), .A2(n1242), .ZN(n1262) );
NOR2_X1 U968 ( .A1(n1307), .A2(n1119), .ZN(n1096) );
AND3_X1 U969 ( .A1(n1093), .A2(n1247), .A3(n1105), .ZN(n1305) );
NOR2_X1 U970 ( .A1(n1118), .A2(n1281), .ZN(n1105) );
INV_X1 U971 ( .A(n1299), .ZN(n1281) );
NOR2_X1 U972 ( .A1(n1288), .A2(n1099), .ZN(n1093) );
XOR2_X1 U973 ( .A(n1237), .B(n1308), .Z(G12) );
XOR2_X1 U974 ( .A(KEYINPUT3), .B(G110), .Z(n1308) );
AND3_X1 U975 ( .A1(n1106), .A2(n1241), .A3(n1097), .ZN(n1237) );
NOR2_X1 U976 ( .A1(n1119), .A2(n1263), .ZN(n1097) );
INV_X1 U977 ( .A(n1307), .ZN(n1263) );
XOR2_X1 U978 ( .A(n1309), .B(n1124), .Z(n1307) );
INV_X1 U979 ( .A(n1192), .ZN(n1124) );
NOR2_X1 U980 ( .A1(n1198), .A2(G902), .ZN(n1192) );
INV_X1 U981 ( .A(n1195), .ZN(n1198) );
XNOR2_X1 U982 ( .A(n1310), .B(n1311), .ZN(n1195) );
XOR2_X1 U983 ( .A(n1145), .B(n1312), .Z(n1311) );
XNOR2_X1 U984 ( .A(n1313), .B(n1314), .ZN(n1312) );
NOR2_X1 U985 ( .A1(G143), .A2(KEYINPUT2), .ZN(n1314) );
NAND2_X1 U986 ( .A1(KEYINPUT42), .A2(n1315), .ZN(n1313) );
INV_X1 U987 ( .A(G131), .ZN(n1315) );
XOR2_X1 U988 ( .A(G140), .B(G125), .Z(n1145) );
XOR2_X1 U989 ( .A(n1316), .B(n1317), .Z(n1310) );
AND3_X1 U990 ( .A1(G214), .A2(n1082), .A3(n1318), .ZN(n1317) );
XNOR2_X1 U991 ( .A(G146), .B(n1319), .ZN(n1316) );
NOR2_X1 U992 ( .A1(KEYINPUT24), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U993 ( .A(n1321), .B(n1322), .ZN(n1320) );
XNOR2_X1 U994 ( .A(n1323), .B(n1324), .ZN(n1322) );
NOR2_X1 U995 ( .A1(G104), .A2(KEYINPUT15), .ZN(n1324) );
NAND2_X1 U996 ( .A1(KEYINPUT57), .A2(n1196), .ZN(n1309) );
INV_X1 U997 ( .A(G475), .ZN(n1196) );
XOR2_X1 U998 ( .A(n1325), .B(n1189), .Z(n1119) );
INV_X1 U999 ( .A(G478), .ZN(n1189) );
NAND2_X1 U1000 ( .A1(n1326), .A2(n1190), .ZN(n1325) );
NAND2_X1 U1001 ( .A1(n1327), .A2(n1328), .ZN(n1190) );
NAND2_X1 U1002 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1003 ( .A(KEYINPUT19), .B(n1331), .Z(n1327) );
NOR2_X1 U1004 ( .A1(n1329), .A2(n1330), .ZN(n1331) );
NAND3_X1 U1005 ( .A1(G234), .A2(n1082), .A3(G217), .ZN(n1330) );
XNOR2_X1 U1006 ( .A(n1332), .B(n1333), .ZN(n1329) );
XNOR2_X1 U1007 ( .A(n1334), .B(n1321), .ZN(n1333) );
NAND2_X1 U1008 ( .A1(KEYINPUT30), .A2(G134), .ZN(n1334) );
XOR2_X1 U1009 ( .A(n1335), .B(n1336), .Z(n1332) );
XNOR2_X1 U1010 ( .A(G116), .B(n1075), .ZN(n1336) );
INV_X1 U1011 ( .A(G107), .ZN(n1075) );
NAND2_X1 U1012 ( .A1(n1337), .A2(n1338), .ZN(n1335) );
NAND2_X1 U1013 ( .A1(G143), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1014 ( .A(KEYINPUT60), .B(n1340), .Z(n1337) );
NOR2_X1 U1015 ( .A1(G143), .A2(n1339), .ZN(n1340) );
XNOR2_X1 U1016 ( .A(KEYINPUT55), .B(n1341), .ZN(n1326) );
NOR4_X1 U1017 ( .A1(n1108), .A2(n1100), .A3(n1301), .A4(n1099), .ZN(n1241) );
INV_X1 U1018 ( .A(n1287), .ZN(n1099) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1342), .ZN(n1287) );
XOR2_X1 U1020 ( .A(KEYINPUT23), .B(n1343), .Z(n1342) );
INV_X1 U1021 ( .A(n1247), .ZN(n1301) );
NAND2_X1 U1022 ( .A1(n1289), .A2(n1344), .ZN(n1247) );
NAND2_X1 U1023 ( .A1(n1291), .A2(n1345), .ZN(n1344) );
INV_X1 U1024 ( .A(G898), .ZN(n1345) );
AND3_X1 U1025 ( .A1(G902), .A2(n1085), .A3(G953), .ZN(n1291) );
NAND3_X1 U1026 ( .A1(n1085), .A2(n1082), .A3(G952), .ZN(n1289) );
NAND2_X1 U1027 ( .A1(n1346), .A2(G237), .ZN(n1085) );
INV_X1 U1028 ( .A(n1288), .ZN(n1100) );
XOR2_X1 U1029 ( .A(n1127), .B(n1129), .Z(n1288) );
INV_X1 U1030 ( .A(G469), .ZN(n1129) );
NAND2_X1 U1031 ( .A1(n1347), .A2(n1341), .ZN(n1127) );
XNOR2_X1 U1032 ( .A(n1348), .B(n1224), .ZN(n1347) );
XOR2_X1 U1033 ( .A(n1349), .B(n1350), .Z(n1224) );
XNOR2_X1 U1034 ( .A(n1200), .B(n1351), .ZN(n1350) );
XNOR2_X1 U1035 ( .A(n1149), .B(n1352), .ZN(n1349) );
XOR2_X1 U1036 ( .A(G143), .B(n1353), .Z(n1149) );
NOR2_X1 U1037 ( .A1(KEYINPUT12), .A2(n1354), .ZN(n1348) );
XNOR2_X1 U1038 ( .A(n1228), .B(n1355), .ZN(n1354) );
NAND2_X1 U1039 ( .A1(G227), .A2(n1082), .ZN(n1228) );
INV_X1 U1040 ( .A(n1242), .ZN(n1108) );
NOR2_X1 U1041 ( .A1(n1111), .A2(n1110), .ZN(n1242) );
INV_X1 U1042 ( .A(n1283), .ZN(n1110) );
NAND2_X1 U1043 ( .A1(G214), .A2(n1356), .ZN(n1283) );
XOR2_X1 U1044 ( .A(n1357), .B(n1122), .Z(n1111) );
NAND2_X1 U1045 ( .A1(n1358), .A2(n1341), .ZN(n1122) );
XOR2_X1 U1046 ( .A(n1359), .B(n1231), .Z(n1358) );
XNOR2_X1 U1047 ( .A(n1360), .B(n1361), .ZN(n1231) );
XNOR2_X1 U1048 ( .A(n1362), .B(n1174), .ZN(n1361) );
XNOR2_X1 U1049 ( .A(n1363), .B(G110), .ZN(n1174) );
NAND2_X1 U1050 ( .A1(KEYINPUT39), .A2(n1321), .ZN(n1363) );
XOR2_X1 U1051 ( .A(G122), .B(KEYINPUT38), .Z(n1321) );
NAND2_X1 U1052 ( .A1(G224), .A2(n1082), .ZN(n1362) );
XOR2_X1 U1053 ( .A(n1364), .B(n1365), .Z(n1360) );
NOR2_X1 U1054 ( .A1(KEYINPUT54), .A2(n1366), .ZN(n1365) );
XNOR2_X1 U1055 ( .A(n1367), .B(n1176), .ZN(n1366) );
XOR2_X1 U1056 ( .A(n1368), .B(n1369), .Z(n1176) );
NOR2_X1 U1057 ( .A1(KEYINPUT20), .A2(n1323), .ZN(n1369) );
NAND2_X1 U1058 ( .A1(KEYINPUT45), .A2(n1175), .ZN(n1367) );
XOR2_X1 U1059 ( .A(n1370), .B(n1352), .Z(n1175) );
XOR2_X1 U1060 ( .A(G101), .B(G107), .Z(n1352) );
NAND2_X1 U1061 ( .A1(KEYINPUT46), .A2(n1200), .ZN(n1370) );
INV_X1 U1062 ( .A(G104), .ZN(n1200) );
XNOR2_X1 U1063 ( .A(G125), .B(KEYINPUT61), .ZN(n1364) );
NOR2_X1 U1064 ( .A1(KEYINPUT9), .A2(n1261), .ZN(n1359) );
NAND2_X1 U1065 ( .A1(KEYINPUT56), .A2(n1123), .ZN(n1357) );
NAND2_X1 U1066 ( .A1(G210), .A2(n1356), .ZN(n1123) );
NAND2_X1 U1067 ( .A1(n1318), .A2(n1341), .ZN(n1356) );
NOR2_X1 U1068 ( .A1(n1299), .A2(n1282), .ZN(n1106) );
INV_X1 U1069 ( .A(n1118), .ZN(n1282) );
XNOR2_X1 U1070 ( .A(n1371), .B(n1372), .ZN(n1118) );
NOR2_X1 U1071 ( .A1(n1343), .A2(n1184), .ZN(n1372) );
INV_X1 U1072 ( .A(G217), .ZN(n1184) );
AND2_X1 U1073 ( .A1(n1346), .A2(n1341), .ZN(n1343) );
XNOR2_X1 U1074 ( .A(KEYINPUT14), .B(G234), .ZN(n1346) );
NAND2_X1 U1075 ( .A1(n1373), .A2(n1341), .ZN(n1371) );
XNOR2_X1 U1076 ( .A(KEYINPUT33), .B(n1374), .ZN(n1373) );
INV_X1 U1077 ( .A(n1182), .ZN(n1374) );
XNOR2_X1 U1078 ( .A(n1375), .B(n1376), .ZN(n1182) );
XOR2_X1 U1079 ( .A(G119), .B(n1377), .Z(n1376) );
XOR2_X1 U1080 ( .A(G137), .B(G125), .Z(n1377) );
XNOR2_X1 U1081 ( .A(n1223), .B(n1378), .ZN(n1375) );
XOR2_X1 U1082 ( .A(n1379), .B(n1353), .Z(n1378) );
XNOR2_X1 U1083 ( .A(n1339), .B(G146), .ZN(n1353) );
INV_X1 U1084 ( .A(G128), .ZN(n1339) );
AND3_X1 U1085 ( .A1(G221), .A2(n1082), .A3(G234), .ZN(n1379) );
INV_X1 U1086 ( .A(n1355), .ZN(n1223) );
XNOR2_X1 U1087 ( .A(G110), .B(G140), .ZN(n1355) );
XOR2_X1 U1088 ( .A(n1380), .B(n1134), .Z(n1299) );
NAND3_X1 U1089 ( .A1(n1381), .A2(n1341), .A3(n1382), .ZN(n1134) );
NAND3_X1 U1090 ( .A1(n1211), .A2(n1383), .A3(n1384), .ZN(n1382) );
XOR2_X1 U1091 ( .A(n1385), .B(n1386), .Z(n1384) );
NOR2_X1 U1092 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
INV_X1 U1093 ( .A(n1217), .ZN(n1387) );
INV_X1 U1094 ( .A(G902), .ZN(n1341) );
NAND2_X1 U1095 ( .A1(n1389), .A2(n1390), .ZN(n1381) );
NAND2_X1 U1096 ( .A1(n1211), .A2(n1383), .ZN(n1390) );
INV_X1 U1097 ( .A(KEYINPUT29), .ZN(n1383) );
XNOR2_X1 U1098 ( .A(n1351), .B(n1261), .ZN(n1211) );
XOR2_X1 U1099 ( .A(G128), .B(n1391), .Z(n1261) );
NOR2_X1 U1100 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
AND3_X1 U1101 ( .A1(n1394), .A2(n1395), .A3(G143), .ZN(n1393) );
NOR2_X1 U1102 ( .A1(n1396), .A2(n1394), .ZN(n1392) );
INV_X1 U1103 ( .A(KEYINPUT40), .ZN(n1394) );
XNOR2_X1 U1104 ( .A(n1395), .B(G143), .ZN(n1396) );
INV_X1 U1105 ( .A(G146), .ZN(n1395) );
AND2_X1 U1106 ( .A1(n1397), .A2(n1398), .ZN(n1351) );
NAND2_X1 U1107 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
XOR2_X1 U1108 ( .A(KEYINPUT11), .B(n1401), .Z(n1397) );
NOR2_X1 U1109 ( .A1(n1399), .A2(n1400), .ZN(n1401) );
XNOR2_X1 U1110 ( .A(G134), .B(n1402), .ZN(n1400) );
XOR2_X1 U1111 ( .A(KEYINPUT58), .B(G137), .Z(n1402) );
XNOR2_X1 U1112 ( .A(G131), .B(KEYINPUT49), .ZN(n1399) );
XOR2_X1 U1113 ( .A(n1403), .B(n1386), .Z(n1389) );
XOR2_X1 U1114 ( .A(n1218), .B(KEYINPUT28), .Z(n1386) );
XOR2_X1 U1115 ( .A(G101), .B(n1404), .Z(n1218) );
AND3_X1 U1116 ( .A1(G210), .A2(n1082), .A3(n1318), .ZN(n1404) );
INV_X1 U1117 ( .A(G237), .ZN(n1318) );
INV_X1 U1118 ( .A(G953), .ZN(n1082) );
NOR2_X1 U1119 ( .A1(n1217), .A2(n1388), .ZN(n1403) );
INV_X1 U1120 ( .A(KEYINPUT41), .ZN(n1388) );
XNOR2_X1 U1121 ( .A(n1405), .B(n1368), .ZN(n1217) );
XOR2_X1 U1122 ( .A(G116), .B(G119), .Z(n1368) );
NAND2_X1 U1123 ( .A1(KEYINPUT63), .A2(n1323), .ZN(n1405) );
INV_X1 U1124 ( .A(G113), .ZN(n1323) );
NAND2_X1 U1125 ( .A1(KEYINPUT59), .A2(G472), .ZN(n1380) );
endmodule


