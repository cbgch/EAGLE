//Key = 0011000101001110010111011010110001100010001000011100110000111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327;

XOR2_X1 U724 ( .A(n1003), .B(n1004), .Z(G9) );
NAND4_X1 U725 ( .A1(KEYINPUT48), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
INV_X1 U727 ( .A(n1010), .ZN(n1009) );
XOR2_X1 U728 ( .A(n1011), .B(KEYINPUT43), .Z(n1008) );
NOR2_X1 U729 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR3_X1 U730 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U731 ( .A1(KEYINPUT58), .A2(n1017), .ZN(n1015) );
NOR4_X1 U732 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NAND2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NAND3_X1 U734 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1014) );
NAND2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U737 ( .A1(n1022), .A2(n1031), .A3(n1032), .ZN(n1030) );
NAND2_X1 U738 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U740 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U742 ( .A1(KEYINPUT58), .A2(n1023), .ZN(n1037) );
NAND2_X1 U743 ( .A1(n1007), .A2(n1041), .ZN(n1033) );
NAND2_X1 U744 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U745 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U746 ( .A1(n1007), .A2(n1046), .A3(n1035), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U748 ( .A1(n1022), .A2(n1049), .ZN(n1048) );
OR2_X1 U749 ( .A1(n1050), .A2(n1005), .ZN(n1049) );
NAND2_X1 U750 ( .A1(n1032), .A2(n1051), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1011), .A2(n1052), .ZN(n1051) );
NAND2_X1 U752 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U753 ( .A(n1021), .ZN(n1027) );
NOR3_X1 U754 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1012) );
INV_X1 U755 ( .A(n1024), .ZN(n1055) );
NAND4_X1 U756 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1024) );
NOR4_X1 U757 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
XOR2_X1 U758 ( .A(n1064), .B(n1065), .Z(n1063) );
XNOR2_X1 U759 ( .A(G469), .B(KEYINPUT4), .ZN(n1065) );
XOR2_X1 U760 ( .A(n1066), .B(n1067), .Z(n1062) );
XOR2_X1 U761 ( .A(KEYINPUT3), .B(G475), .Z(n1067) );
NOR2_X1 U762 ( .A1(n1068), .A2(KEYINPUT39), .ZN(n1066) );
NOR3_X1 U763 ( .A1(n1069), .A2(n1070), .A3(n1044), .ZN(n1058) );
XOR2_X1 U764 ( .A(n1071), .B(n1072), .Z(n1056) );
NAND2_X1 U765 ( .A1(KEYINPUT20), .A2(n1073), .ZN(n1072) );
XOR2_X1 U766 ( .A(n1074), .B(n1075), .Z(G72) );
NOR2_X1 U767 ( .A1(n1076), .A2(n1025), .ZN(n1075) );
NOR2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NAND2_X1 U770 ( .A1(n1081), .A2(n1025), .ZN(n1080) );
XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
XOR2_X1 U773 ( .A(KEYINPUT2), .B(n1086), .Z(n1085) );
INV_X1 U774 ( .A(n1087), .ZN(n1084) );
OR3_X1 U775 ( .A1(n1078), .A2(n1083), .A3(n1025), .ZN(n1079) );
XNOR2_X1 U776 ( .A(n1088), .B(n1089), .ZN(n1083) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U779 ( .A(n1094), .B(KEYINPUT53), .Z(n1093) );
NAND2_X1 U780 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U781 ( .A(KEYINPUT40), .B(G140), .Z(n1095) );
NOR2_X1 U782 ( .A1(G140), .A2(n1096), .ZN(n1092) );
NOR2_X1 U783 ( .A1(KEYINPUT0), .A2(n1097), .ZN(n1090) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(n1088) );
XOR2_X1 U786 ( .A(G131), .B(G128), .Z(n1101) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U788 ( .A1(n1104), .A2(G953), .ZN(n1103) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U790 ( .A(n1107), .B(n1108), .Z(n1102) );
NOR2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U793 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U794 ( .A1(KEYINPUT18), .A2(n1115), .ZN(n1113) );
NAND3_X1 U795 ( .A1(n1116), .A2(n1117), .A3(KEYINPUT47), .ZN(n1107) );
NAND2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
INV_X1 U797 ( .A(KEYINPUT55), .ZN(n1119) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
OR2_X1 U799 ( .A1(n1025), .A2(G224), .ZN(n1121) );
INV_X1 U800 ( .A(n1109), .ZN(n1120) );
NAND3_X1 U801 ( .A1(n1122), .A2(n1025), .A3(KEYINPUT55), .ZN(n1116) );
NAND2_X1 U802 ( .A1(G898), .A2(G224), .ZN(n1122) );
NOR2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U804 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NOR2_X1 U806 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XNOR2_X1 U807 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND2_X1 U808 ( .A1(n1127), .A2(G478), .ZN(n1130) );
NOR2_X1 U809 ( .A1(n1123), .A2(n1132), .ZN(G60) );
NOR3_X1 U810 ( .A1(n1068), .A2(n1133), .A3(n1134), .ZN(n1132) );
AND3_X1 U811 ( .A1(n1135), .A2(G475), .A3(n1127), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1136), .A2(n1135), .ZN(n1133) );
AND2_X1 U813 ( .A1(n1016), .A2(G475), .ZN(n1136) );
XNOR2_X1 U814 ( .A(G104), .B(n1137), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1123), .A2(n1138), .ZN(G57) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR3_X1 U818 ( .A1(n1143), .A2(KEYINPUT30), .A3(n1144), .ZN(n1142) );
INV_X1 U819 ( .A(G472), .ZN(n1144) );
NOR2_X1 U820 ( .A1(n1123), .A2(n1145), .ZN(G54) );
XOR2_X1 U821 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U824 ( .A1(n1127), .A2(G469), .ZN(n1151) );
NAND2_X1 U825 ( .A1(KEYINPUT60), .A2(n1152), .ZN(n1150) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1146) );
XOR2_X1 U827 ( .A(n1155), .B(G128), .Z(n1153) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U829 ( .A(KEYINPUT21), .B(KEYINPUT15), .Z(n1157) );
XOR2_X1 U830 ( .A(n1098), .B(n1158), .Z(n1156) );
NOR2_X1 U831 ( .A1(n1123), .A2(n1159), .ZN(G51) );
XOR2_X1 U832 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U833 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U834 ( .A1(n1127), .A2(n1164), .ZN(n1162) );
INV_X1 U835 ( .A(n1143), .ZN(n1127) );
NAND2_X1 U836 ( .A1(G902), .A2(n1016), .ZN(n1143) );
NAND4_X1 U837 ( .A1(n1086), .A2(n1087), .A3(n1165), .A4(n1166), .ZN(n1016) );
XNOR2_X1 U838 ( .A(KEYINPUT16), .B(n1105), .ZN(n1166) );
NAND3_X1 U839 ( .A1(n1167), .A2(n1137), .A3(n1168), .ZN(n1105) );
OR2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND4_X1 U841 ( .A1(n1050), .A2(n1007), .A3(n1010), .A4(n1171), .ZN(n1137) );
NAND2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
NAND2_X1 U843 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND3_X1 U844 ( .A1(n1007), .A2(n1010), .A3(n1005), .ZN(n1174) );
NAND2_X1 U845 ( .A1(n1032), .A2(n1175), .ZN(n1173) );
NAND2_X1 U846 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND4_X1 U847 ( .A1(n1178), .A2(n1023), .A3(n1179), .A4(n1169), .ZN(n1177) );
INV_X1 U848 ( .A(KEYINPUT12), .ZN(n1169) );
INV_X1 U849 ( .A(n1106), .ZN(n1165) );
NAND4_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1106) );
NAND3_X1 U851 ( .A1(n1022), .A2(n1005), .A3(n1184), .ZN(n1181) );
NAND2_X1 U852 ( .A1(n1185), .A2(n1179), .ZN(n1180) );
NOR3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1087) );
AND2_X1 U854 ( .A1(n1035), .A2(n1189), .ZN(n1186) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1192), .A2(n1171), .ZN(n1191) );
NAND2_X1 U857 ( .A1(n1032), .A2(n1193), .ZN(n1190) );
AND4_X1 U858 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1086) );
NOR2_X1 U859 ( .A1(n1025), .A2(G952), .ZN(n1123) );
XOR2_X1 U860 ( .A(G146), .B(n1187), .Z(G48) );
NOR3_X1 U861 ( .A1(n1198), .A2(n1042), .A3(n1199), .ZN(n1187) );
XOR2_X1 U862 ( .A(n1200), .B(n1201), .Z(G45) );
NAND2_X1 U863 ( .A1(KEYINPUT23), .A2(n1188), .ZN(n1201) );
AND4_X1 U864 ( .A1(n1202), .A2(n1179), .A3(n1203), .A4(n1204), .ZN(n1188) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(G42) );
NAND2_X1 U866 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1206) );
NAND3_X1 U867 ( .A1(n1171), .A2(n1207), .A3(n1192), .ZN(n1205) );
XOR2_X1 U868 ( .A(KEYINPUT1), .B(n1035), .Z(n1207) );
XOR2_X1 U869 ( .A(n1208), .B(n1209), .Z(G39) );
NOR2_X1 U870 ( .A1(KEYINPUT41), .A2(n1098), .ZN(n1209) );
INV_X1 U871 ( .A(G137), .ZN(n1098) );
NOR3_X1 U872 ( .A1(n1210), .A2(n1199), .A3(n1020), .ZN(n1208) );
XOR2_X1 U873 ( .A(KEYINPUT52), .B(n1035), .Z(n1210) );
XNOR2_X1 U874 ( .A(G134), .B(n1194), .ZN(G36) );
NAND3_X1 U875 ( .A1(n1035), .A2(n1005), .A3(n1202), .ZN(n1194) );
XOR2_X1 U876 ( .A(n1195), .B(n1211), .Z(G33) );
NAND2_X1 U877 ( .A1(KEYINPUT61), .A2(G131), .ZN(n1211) );
NAND3_X1 U878 ( .A1(n1035), .A2(n1050), .A3(n1202), .ZN(n1195) );
AND4_X1 U879 ( .A1(n1039), .A2(n1171), .A3(n1040), .A4(n1212), .ZN(n1202) );
INV_X1 U880 ( .A(n1018), .ZN(n1035) );
NAND2_X1 U881 ( .A1(n1045), .A2(n1213), .ZN(n1018) );
XNOR2_X1 U882 ( .A(G128), .B(n1196), .ZN(G30) );
NAND3_X1 U883 ( .A1(n1005), .A2(n1179), .A3(n1193), .ZN(n1196) );
INV_X1 U884 ( .A(n1199), .ZN(n1193) );
NAND4_X1 U885 ( .A1(n1039), .A2(n1171), .A3(n1061), .A4(n1212), .ZN(n1199) );
XOR2_X1 U886 ( .A(G101), .B(n1214), .Z(G3) );
NOR4_X1 U887 ( .A1(KEYINPUT8), .A2(n1011), .A3(n1020), .A4(n1176), .ZN(n1214) );
INV_X1 U888 ( .A(n1032), .ZN(n1020) );
XOR2_X1 U889 ( .A(n1096), .B(n1197), .Z(G27) );
NAND3_X1 U890 ( .A1(n1192), .A2(n1179), .A3(n1022), .ZN(n1197) );
AND3_X1 U891 ( .A1(n1050), .A2(n1212), .A3(n1023), .ZN(n1192) );
NAND2_X1 U892 ( .A1(n1021), .A2(n1215), .ZN(n1212) );
NAND4_X1 U893 ( .A1(G902), .A2(G953), .A3(n1216), .A4(n1078), .ZN(n1215) );
INV_X1 U894 ( .A(G900), .ZN(n1078) );
XOR2_X1 U895 ( .A(G122), .B(n1217), .Z(G24) );
NOR2_X1 U896 ( .A1(n1042), .A2(n1218), .ZN(n1217) );
XOR2_X1 U897 ( .A(KEYINPUT38), .B(n1185), .Z(n1218) );
AND4_X1 U898 ( .A1(n1022), .A2(n1007), .A3(n1219), .A4(n1203), .ZN(n1185) );
NOR2_X1 U899 ( .A1(n1220), .A2(n1178), .ZN(n1219) );
NOR2_X1 U900 ( .A1(n1061), .A2(n1221), .ZN(n1007) );
XOR2_X1 U901 ( .A(n1222), .B(n1182), .Z(G21) );
NAND4_X1 U902 ( .A1(n1010), .A2(n1061), .A3(n1022), .A4(n1223), .ZN(n1182) );
AND2_X1 U903 ( .A1(n1032), .A2(n1039), .ZN(n1223) );
INV_X1 U904 ( .A(n1040), .ZN(n1061) );
XNOR2_X1 U905 ( .A(G116), .B(n1224), .ZN(G18) );
NAND4_X1 U906 ( .A1(KEYINPUT9), .A2(n1184), .A3(n1022), .A4(n1005), .ZN(n1224) );
NOR2_X1 U907 ( .A1(n1203), .A2(n1220), .ZN(n1005) );
XNOR2_X1 U908 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U909 ( .A1(n1022), .A2(n1050), .A3(n1184), .ZN(n1183) );
INV_X1 U910 ( .A(n1176), .ZN(n1184) );
NAND3_X1 U911 ( .A1(n1040), .A2(n1010), .A3(n1039), .ZN(n1176) );
XOR2_X1 U912 ( .A(n1221), .B(KEYINPUT32), .Z(n1039) );
INV_X1 U913 ( .A(n1198), .ZN(n1050) );
NAND2_X1 U914 ( .A1(n1220), .A2(n1203), .ZN(n1198) );
NOR2_X1 U915 ( .A1(n1225), .A2(n1053), .ZN(n1022) );
INV_X1 U916 ( .A(n1057), .ZN(n1053) );
XOR2_X1 U917 ( .A(n1226), .B(n1170), .Z(G12) );
NAND4_X1 U918 ( .A1(n1032), .A2(n1023), .A3(n1010), .A4(n1171), .ZN(n1170) );
INV_X1 U919 ( .A(n1011), .ZN(n1171) );
NAND2_X1 U920 ( .A1(n1225), .A2(n1057), .ZN(n1011) );
NAND2_X1 U921 ( .A1(n1227), .A2(G221), .ZN(n1057) );
XOR2_X1 U922 ( .A(n1228), .B(KEYINPUT50), .Z(n1227) );
INV_X1 U923 ( .A(n1054), .ZN(n1225) );
XNOR2_X1 U924 ( .A(G469), .B(n1229), .ZN(n1054) );
NOR2_X1 U925 ( .A1(KEYINPUT11), .A2(n1064), .ZN(n1229) );
NAND3_X1 U926 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1064) );
NAND2_X1 U927 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
XOR2_X1 U928 ( .A(n1235), .B(n1236), .Z(n1233) );
OR3_X1 U929 ( .A1(n1235), .A2(n1236), .A3(n1234), .ZN(n1230) );
INV_X1 U930 ( .A(KEYINPUT10), .ZN(n1234) );
XOR2_X1 U931 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U932 ( .A(KEYINPUT35), .B(n1239), .Z(n1238) );
XOR2_X1 U933 ( .A(n1148), .B(n1158), .Z(n1237) );
XOR2_X1 U934 ( .A(n1240), .B(n1100), .Z(n1148) );
NAND2_X1 U935 ( .A1(KEYINPUT59), .A2(n1241), .ZN(n1100) );
NAND3_X1 U936 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1235) );
NAND2_X1 U937 ( .A1(KEYINPUT27), .A2(n1245), .ZN(n1244) );
OR2_X1 U938 ( .A1(n1246), .A2(n1154), .ZN(n1245) );
OR3_X1 U939 ( .A1(n1247), .A2(KEYINPUT27), .A3(n1246), .ZN(n1243) );
AND2_X1 U940 ( .A1(KEYINPUT42), .A2(n1154), .ZN(n1247) );
NAND3_X1 U941 ( .A1(KEYINPUT42), .A2(n1154), .A3(n1246), .ZN(n1242) );
XNOR2_X1 U942 ( .A(n1226), .B(n1248), .ZN(n1246) );
NOR2_X1 U943 ( .A1(G140), .A2(KEYINPUT57), .ZN(n1248) );
NOR2_X1 U944 ( .A1(n1077), .A2(G953), .ZN(n1154) );
INV_X1 U945 ( .A(G227), .ZN(n1077) );
NOR2_X1 U946 ( .A1(n1042), .A2(n1178), .ZN(n1010) );
AND2_X1 U947 ( .A1(n1021), .A2(n1249), .ZN(n1178) );
NAND3_X1 U948 ( .A1(n1109), .A2(n1216), .A3(G902), .ZN(n1249) );
NOR2_X1 U949 ( .A1(n1025), .A2(G898), .ZN(n1109) );
NAND3_X1 U950 ( .A1(n1216), .A2(n1025), .A3(G952), .ZN(n1021) );
NAND2_X1 U951 ( .A1(G237), .A2(G234), .ZN(n1216) );
INV_X1 U952 ( .A(n1179), .ZN(n1042) );
NOR2_X1 U953 ( .A1(n1045), .A2(n1044), .ZN(n1179) );
INV_X1 U954 ( .A(n1213), .ZN(n1044) );
NAND2_X1 U955 ( .A1(G214), .A2(n1250), .ZN(n1213) );
XOR2_X1 U956 ( .A(n1073), .B(n1164), .Z(n1045) );
INV_X1 U957 ( .A(n1071), .ZN(n1164) );
NAND2_X1 U958 ( .A1(G210), .A2(n1250), .ZN(n1071) );
NAND2_X1 U959 ( .A1(n1232), .A2(n1251), .ZN(n1250) );
INV_X1 U960 ( .A(G237), .ZN(n1251) );
NAND2_X1 U961 ( .A1(n1252), .A2(n1232), .ZN(n1073) );
XOR2_X1 U962 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U963 ( .A(n1255), .B(n1256), .Z(n1254) );
INV_X1 U964 ( .A(n1163), .ZN(n1256) );
XOR2_X1 U965 ( .A(n1257), .B(n1258), .Z(n1163) );
XOR2_X1 U966 ( .A(G128), .B(G125), .Z(n1258) );
XOR2_X1 U967 ( .A(n1259), .B(n1260), .Z(n1257) );
NAND2_X1 U968 ( .A1(G224), .A2(n1025), .ZN(n1259) );
NAND2_X1 U969 ( .A1(KEYINPUT34), .A2(n1261), .ZN(n1255) );
XOR2_X1 U970 ( .A(KEYINPUT19), .B(n1160), .Z(n1261) );
XOR2_X1 U971 ( .A(n1114), .B(n1262), .Z(n1160) );
NOR2_X1 U972 ( .A1(KEYINPUT36), .A2(n1263), .ZN(n1262) );
NOR3_X1 U973 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
NOR2_X1 U974 ( .A1(n1267), .A2(n1111), .ZN(n1266) );
NOR2_X1 U975 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U976 ( .A(KEYINPUT33), .B(n1240), .Z(n1269) );
INV_X1 U977 ( .A(KEYINPUT26), .ZN(n1268) );
AND3_X1 U978 ( .A1(n1111), .A2(n1240), .A3(KEYINPUT26), .ZN(n1265) );
XOR2_X1 U979 ( .A(G113), .B(n1270), .Z(n1111) );
NOR2_X1 U980 ( .A1(KEYINPUT44), .A2(n1271), .ZN(n1270) );
XOR2_X1 U981 ( .A(n1222), .B(n1272), .Z(n1271) );
INV_X1 U982 ( .A(G119), .ZN(n1222) );
NOR2_X1 U983 ( .A1(KEYINPUT26), .A2(n1240), .ZN(n1264) );
INV_X1 U984 ( .A(n1115), .ZN(n1240) );
XNOR2_X1 U985 ( .A(G101), .B(n1273), .ZN(n1115) );
XOR2_X1 U986 ( .A(G107), .B(G104), .Z(n1273) );
XOR2_X1 U987 ( .A(n1226), .B(n1274), .Z(n1114) );
XNOR2_X1 U988 ( .A(KEYINPUT6), .B(KEYINPUT56), .ZN(n1253) );
NOR2_X1 U989 ( .A1(n1221), .A2(n1040), .ZN(n1023) );
XOR2_X1 U990 ( .A(n1275), .B(n1128), .Z(n1040) );
AND2_X1 U991 ( .A1(G217), .A2(n1228), .ZN(n1128) );
NAND2_X1 U992 ( .A1(G234), .A2(n1232), .ZN(n1228) );
NAND2_X1 U993 ( .A1(n1276), .A2(n1232), .ZN(n1275) );
XOR2_X1 U994 ( .A(n1126), .B(KEYINPUT51), .Z(n1276) );
XOR2_X1 U995 ( .A(n1277), .B(n1278), .Z(n1126) );
XOR2_X1 U996 ( .A(n1279), .B(n1152), .Z(n1278) );
XOR2_X1 U997 ( .A(G110), .B(G140), .Z(n1152) );
XOR2_X1 U998 ( .A(n1280), .B(n1281), .Z(n1277) );
XOR2_X1 U999 ( .A(n1282), .B(KEYINPUT17), .Z(n1280) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1001 ( .A(n1060), .B(KEYINPUT7), .ZN(n1221) );
XNOR2_X1 U1002 ( .A(n1284), .B(G472), .ZN(n1060) );
NAND2_X1 U1003 ( .A1(n1285), .A2(n1232), .ZN(n1284) );
INV_X1 U1004 ( .A(G902), .ZN(n1232) );
XOR2_X1 U1005 ( .A(n1286), .B(n1287), .Z(n1285) );
INV_X1 U1006 ( .A(n1139), .ZN(n1287) );
XOR2_X1 U1007 ( .A(n1288), .B(G101), .Z(n1139) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1009 ( .A(n1141), .B(KEYINPUT5), .Z(n1286) );
XOR2_X1 U1010 ( .A(n1290), .B(n1291), .Z(n1141) );
XOR2_X1 U1011 ( .A(n1281), .B(n1260), .Z(n1291) );
AND2_X1 U1012 ( .A1(n1292), .A2(n1293), .ZN(n1260) );
NAND2_X1 U1013 ( .A1(n1241), .A2(n1294), .ZN(n1293) );
INV_X1 U1014 ( .A(KEYINPUT45), .ZN(n1294) );
XOR2_X1 U1015 ( .A(n1200), .B(G146), .Z(n1241) );
NAND3_X1 U1016 ( .A1(G143), .A2(n1295), .A3(KEYINPUT45), .ZN(n1292) );
XOR2_X1 U1017 ( .A(G119), .B(n1239), .Z(n1281) );
XOR2_X1 U1018 ( .A(G137), .B(G128), .Z(n1239) );
XOR2_X1 U1019 ( .A(n1296), .B(n1272), .Z(n1290) );
XNOR2_X1 U1020 ( .A(G113), .B(n1158), .ZN(n1296) );
XOR2_X1 U1021 ( .A(n1297), .B(n1099), .Z(n1158) );
XNOR2_X1 U1022 ( .A(G131), .B(KEYINPUT62), .ZN(n1297) );
NOR2_X1 U1023 ( .A1(n1204), .A2(n1203), .ZN(n1032) );
XOR2_X1 U1024 ( .A(n1068), .B(G475), .Z(n1203) );
NOR2_X1 U1025 ( .A1(n1135), .A2(G902), .ZN(n1068) );
XOR2_X1 U1026 ( .A(n1298), .B(n1299), .Z(n1135) );
XOR2_X1 U1027 ( .A(n1300), .B(n1301), .Z(n1299) );
NAND3_X1 U1028 ( .A1(G214), .A2(n1289), .A3(KEYINPUT28), .ZN(n1301) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1289) );
NAND2_X1 U1030 ( .A1(n1302), .A2(KEYINPUT29), .ZN(n1300) );
XOR2_X1 U1031 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1032 ( .A(KEYINPUT46), .B(G122), .Z(n1304) );
XNOR2_X1 U1033 ( .A(G104), .B(G113), .ZN(n1303) );
XOR2_X1 U1034 ( .A(n1305), .B(n1306), .Z(n1298) );
NOR2_X1 U1035 ( .A1(KEYINPUT25), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1036 ( .A(n1279), .B(n1308), .ZN(n1307) );
NOR2_X1 U1037 ( .A1(G140), .A2(KEYINPUT63), .ZN(n1308) );
XOR2_X1 U1038 ( .A(n1096), .B(n1295), .Z(n1279) );
INV_X1 U1039 ( .A(G146), .ZN(n1295) );
INV_X1 U1040 ( .A(G125), .ZN(n1096) );
XOR2_X1 U1041 ( .A(G131), .B(n1200), .Z(n1305) );
INV_X1 U1042 ( .A(G143), .ZN(n1200) );
INV_X1 U1043 ( .A(n1220), .ZN(n1204) );
NOR2_X1 U1044 ( .A1(n1309), .A2(n1069), .ZN(n1220) );
NOR3_X1 U1045 ( .A1(G478), .A2(G902), .A3(n1131), .ZN(n1069) );
XNOR2_X1 U1046 ( .A(KEYINPUT24), .B(n1070), .ZN(n1309) );
AND2_X1 U1047 ( .A1(G478), .A2(n1310), .ZN(n1070) );
OR2_X1 U1048 ( .A1(n1131), .A2(G902), .ZN(n1310) );
XNOR2_X1 U1049 ( .A(n1311), .B(n1312), .ZN(n1131) );
NOR2_X1 U1050 ( .A1(KEYINPUT22), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1051 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1052 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND2_X1 U1053 ( .A1(KEYINPUT13), .A2(n1099), .ZN(n1317) );
XNOR2_X1 U1054 ( .A(G134), .B(KEYINPUT14), .ZN(n1099) );
NAND3_X1 U1055 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1316) );
NAND2_X1 U1056 ( .A1(G107), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1057 ( .A1(KEYINPUT54), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1058 ( .A1(n1323), .A2(n1003), .ZN(n1322) );
INV_X1 U1059 ( .A(G107), .ZN(n1003) );
XNOR2_X1 U1060 ( .A(n1321), .B(KEYINPUT31), .ZN(n1323) );
NAND2_X1 U1061 ( .A1(n1324), .A2(n1325), .ZN(n1318) );
INV_X1 U1062 ( .A(KEYINPUT54), .ZN(n1325) );
NAND2_X1 U1063 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
OR3_X1 U1064 ( .A1(n1321), .A2(G107), .A3(KEYINPUT31), .ZN(n1327) );
NAND2_X1 U1065 ( .A1(KEYINPUT31), .A2(n1321), .ZN(n1326) );
XNOR2_X1 U1066 ( .A(n1274), .B(n1272), .ZN(n1321) );
XOR2_X1 U1067 ( .A(G116), .B(KEYINPUT37), .Z(n1272) );
INV_X1 U1068 ( .A(G122), .ZN(n1274) );
XOR2_X1 U1069 ( .A(G143), .B(G128), .Z(n1314) );
NAND2_X1 U1070 ( .A1(G217), .A2(n1283), .ZN(n1311) );
AND2_X1 U1071 ( .A1(G234), .A2(n1025), .ZN(n1283) );
INV_X1 U1072 ( .A(G953), .ZN(n1025) );
INV_X1 U1073 ( .A(G110), .ZN(n1226) );
endmodule


