//Key = 0010110100010101111101111011000001101110111010111101110110111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399;

XNOR2_X1 U765 ( .A(G107), .B(n1072), .ZN(G9) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U768 ( .A1(n1077), .A2(n1078), .A3(G953), .A4(n1079), .ZN(n1076) );
NAND3_X1 U769 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
NAND3_X1 U770 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
INV_X1 U771 ( .A(n1086), .ZN(n1085) );
NOR3_X1 U772 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1084) );
NOR2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U774 ( .A(n1092), .ZN(n1088) );
AND3_X1 U775 ( .A1(KEYINPUT52), .A2(n1093), .A3(n1094), .ZN(n1083) );
NAND4_X1 U776 ( .A1(n1095), .A2(n1092), .A3(KEYINPUT52), .A4(n1086), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U778 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U780 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
INV_X1 U781 ( .A(KEYINPUT17), .ZN(n1103) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1105), .ZN(n1100) );
NAND2_X1 U783 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U784 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1102), .ZN(n1096) );
NAND3_X1 U786 ( .A1(n1110), .A2(n1111), .A3(n1093), .ZN(n1102) );
NAND2_X1 U787 ( .A1(n1094), .A2(n1112), .ZN(n1111) );
NAND2_X1 U788 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1115), .ZN(n1110) );
NAND2_X1 U790 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U791 ( .A1(KEYINPUT17), .A2(n1104), .ZN(n1117) );
NOR3_X1 U792 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1075) );
AND4_X1 U793 ( .A1(n1093), .A2(n1086), .A3(n1118), .A4(n1119), .ZN(n1079) );
NOR3_X1 U794 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
XOR2_X1 U795 ( .A(n1123), .B(n1124), .Z(n1121) );
NOR2_X1 U796 ( .A1(G472), .A2(KEYINPUT35), .ZN(n1124) );
XOR2_X1 U797 ( .A(n1125), .B(n1126), .Z(n1118) );
NOR2_X1 U798 ( .A1(KEYINPUT10), .A2(n1127), .ZN(n1126) );
XOR2_X1 U799 ( .A(KEYINPUT2), .B(G475), .Z(n1127) );
XOR2_X1 U800 ( .A(n1128), .B(n1129), .Z(G72) );
NOR2_X1 U801 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR3_X1 U802 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U803 ( .A1(G953), .A2(n1135), .ZN(n1130) );
XNOR2_X1 U804 ( .A(n1136), .B(n1134), .ZN(n1135) );
NAND2_X1 U805 ( .A1(n1137), .A2(KEYINPUT26), .ZN(n1134) );
XOR2_X1 U806 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U807 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U808 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U809 ( .A1(G125), .A2(KEYINPUT12), .ZN(n1143) );
NAND2_X1 U810 ( .A1(KEYINPUT21), .A2(n1144), .ZN(n1142) );
XOR2_X1 U811 ( .A(KEYINPUT7), .B(G140), .Z(n1140) );
XOR2_X1 U812 ( .A(n1145), .B(n1146), .Z(n1138) );
XNOR2_X1 U813 ( .A(n1147), .B(n1148), .ZN(n1145) );
NOR2_X1 U814 ( .A1(KEYINPUT9), .A2(n1149), .ZN(n1128) );
NOR2_X1 U815 ( .A1(n1150), .A2(n1132), .ZN(n1149) );
AND2_X1 U816 ( .A1(G227), .A2(G900), .ZN(n1150) );
NAND3_X1 U817 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(G69) );
NAND2_X1 U818 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U819 ( .A1(KEYINPUT24), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U820 ( .A(n1157), .B(n1082), .ZN(n1156) );
NAND2_X1 U821 ( .A1(G953), .A2(n1158), .ZN(n1154) );
NAND4_X1 U822 ( .A1(G953), .A2(n1158), .A3(KEYINPUT24), .A4(n1157), .ZN(n1152) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1158) );
OR2_X1 U824 ( .A1(n1157), .A2(KEYINPUT24), .ZN(n1151) );
NAND2_X1 U825 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U826 ( .A1(G953), .A2(n1161), .ZN(n1160) );
NOR3_X1 U827 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(G66) );
AND3_X1 U828 ( .A1(KEYINPUT61), .A2(G953), .A3(G952), .ZN(n1164) );
NOR2_X1 U829 ( .A1(KEYINPUT61), .A2(n1165), .ZN(n1163) );
INV_X1 U830 ( .A(n1166), .ZN(n1165) );
XOR2_X1 U831 ( .A(n1167), .B(n1168), .Z(n1162) );
NOR2_X1 U832 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1171), .ZN(G63) );
XNOR2_X1 U834 ( .A(n1172), .B(n1173), .ZN(n1171) );
AND2_X1 U835 ( .A1(G478), .A2(n1174), .ZN(n1173) );
NOR2_X1 U836 ( .A1(n1166), .A2(n1175), .ZN(G60) );
XOR2_X1 U837 ( .A(n1176), .B(KEYINPUT25), .Z(n1175) );
NAND2_X1 U838 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U840 ( .A1(KEYINPUT5), .A2(n1181), .ZN(n1179) );
OR2_X1 U841 ( .A1(n1182), .A2(KEYINPUT14), .ZN(n1181) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1177) );
NAND2_X1 U843 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U844 ( .A1(n1186), .A2(KEYINPUT5), .ZN(n1185) );
INV_X1 U845 ( .A(n1180), .ZN(n1186) );
NAND2_X1 U846 ( .A1(n1174), .A2(G475), .ZN(n1180) );
INV_X1 U847 ( .A(KEYINPUT14), .ZN(n1184) );
XOR2_X1 U848 ( .A(n1187), .B(G104), .Z(G6) );
NAND2_X1 U849 ( .A1(KEYINPUT13), .A2(n1188), .ZN(n1187) );
NOR3_X1 U850 ( .A1(n1189), .A2(n1166), .A3(n1190), .ZN(G57) );
NOR3_X1 U851 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1191) );
NOR2_X1 U853 ( .A1(n1196), .A2(KEYINPUT0), .ZN(n1194) );
NOR2_X1 U854 ( .A1(n1197), .A2(n1198), .ZN(n1189) );
XNOR2_X1 U855 ( .A(n1199), .B(n1195), .ZN(n1198) );
XOR2_X1 U856 ( .A(n1200), .B(n1201), .Z(n1195) );
NAND2_X1 U857 ( .A1(KEYINPUT18), .A2(n1202), .ZN(n1200) );
NAND2_X1 U858 ( .A1(n1196), .A2(n1203), .ZN(n1199) );
INV_X1 U859 ( .A(KEYINPUT0), .ZN(n1203) );
AND2_X1 U860 ( .A1(n1174), .A2(G472), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1193), .A2(n1192), .ZN(n1197) );
INV_X1 U862 ( .A(KEYINPUT53), .ZN(n1192) );
XNOR2_X1 U863 ( .A(G113), .B(n1204), .ZN(n1193) );
NOR2_X1 U864 ( .A1(n1166), .A2(n1205), .ZN(G54) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U866 ( .A(n1208), .B(n1209), .Z(n1207) );
AND2_X1 U867 ( .A1(G469), .A2(n1174), .ZN(n1209) );
INV_X1 U868 ( .A(n1170), .ZN(n1174) );
NAND3_X1 U869 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1208) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR3_X1 U871 ( .A1(n1214), .A2(n1213), .A3(KEYINPUT45), .ZN(n1211) );
NAND2_X1 U872 ( .A1(KEYINPUT27), .A2(n1215), .ZN(n1214) );
NAND2_X1 U873 ( .A1(n1216), .A2(KEYINPUT45), .ZN(n1210) );
INV_X1 U874 ( .A(n1215), .ZN(n1216) );
XOR2_X1 U875 ( .A(n1217), .B(n1147), .Z(n1215) );
NAND2_X1 U876 ( .A1(KEYINPUT36), .A2(n1218), .ZN(n1217) );
NOR3_X1 U877 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(G51) );
AND2_X1 U878 ( .A1(n1166), .A2(KEYINPUT34), .ZN(n1221) );
NOR2_X1 U879 ( .A1(n1132), .A2(G952), .ZN(n1166) );
NOR3_X1 U880 ( .A1(KEYINPUT34), .A2(G953), .A3(G952), .ZN(n1220) );
XOR2_X1 U881 ( .A(n1222), .B(n1223), .Z(n1219) );
NOR2_X1 U882 ( .A1(n1224), .A2(n1170), .ZN(n1223) );
NAND2_X1 U883 ( .A1(n1225), .A2(n1226), .ZN(n1170) );
NAND2_X1 U884 ( .A1(n1082), .A2(n1136), .ZN(n1226) );
INV_X1 U885 ( .A(n1078), .ZN(n1136) );
NAND4_X1 U886 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1078) );
AND4_X1 U887 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1230) );
NOR2_X1 U888 ( .A1(n1235), .A2(n1236), .ZN(n1229) );
NOR3_X1 U889 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
NOR2_X1 U890 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
INV_X1 U891 ( .A(KEYINPUT30), .ZN(n1241) );
NOR4_X1 U892 ( .A1(n1242), .A2(n1090), .A3(n1243), .A4(n1244), .ZN(n1240) );
INV_X1 U893 ( .A(n1245), .ZN(n1090) );
NOR2_X1 U894 ( .A1(KEYINPUT30), .A2(n1246), .ZN(n1238) );
INV_X1 U895 ( .A(n1247), .ZN(n1237) );
NAND3_X1 U896 ( .A1(n1246), .A2(n1094), .A3(n1248), .ZN(n1228) );
XNOR2_X1 U897 ( .A(KEYINPUT22), .B(n1249), .ZN(n1248) );
NAND2_X1 U898 ( .A1(n1250), .A2(n1251), .ZN(n1227) );
XOR2_X1 U899 ( .A(n1252), .B(KEYINPUT15), .Z(n1250) );
AND2_X1 U900 ( .A1(n1253), .A2(n1254), .ZN(n1082) );
AND4_X1 U901 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
INV_X1 U902 ( .A(n1259), .ZN(n1257) );
NOR4_X1 U903 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1253) );
NOR3_X1 U904 ( .A1(n1116), .A2(n1264), .A3(n1265), .ZN(n1263) );
XNOR2_X1 U905 ( .A(n1098), .B(KEYINPUT1), .ZN(n1264) );
INV_X1 U906 ( .A(n1188), .ZN(n1262) );
NAND2_X1 U907 ( .A1(n1104), .A2(n1074), .ZN(n1188) );
NOR2_X1 U908 ( .A1(n1087), .A2(n1265), .ZN(n1074) );
INV_X1 U909 ( .A(n1098), .ZN(n1087) );
XNOR2_X1 U910 ( .A(KEYINPUT3), .B(n1266), .ZN(n1225) );
NAND2_X1 U911 ( .A1(KEYINPUT37), .A2(n1267), .ZN(n1222) );
XOR2_X1 U912 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U913 ( .A(G125), .B(n1270), .Z(n1269) );
XNOR2_X1 U914 ( .A(n1159), .B(n1271), .ZN(n1268) );
XNOR2_X1 U915 ( .A(n1272), .B(n1273), .ZN(G48) );
NOR2_X1 U916 ( .A1(n1106), .A2(n1252), .ZN(n1273) );
NAND3_X1 U917 ( .A1(n1104), .A2(n1249), .A3(n1274), .ZN(n1252) );
XOR2_X1 U918 ( .A(G143), .B(n1235), .Z(G45) );
AND3_X1 U919 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1235) );
NOR3_X1 U920 ( .A1(n1106), .A2(n1277), .A3(n1278), .ZN(n1276) );
INV_X1 U921 ( .A(n1251), .ZN(n1106) );
XOR2_X1 U922 ( .A(n1234), .B(n1279), .Z(G42) );
NAND2_X1 U923 ( .A1(KEYINPUT47), .A2(G140), .ZN(n1279) );
NAND3_X1 U924 ( .A1(n1104), .A2(n1280), .A3(n1246), .ZN(n1234) );
XNOR2_X1 U925 ( .A(G137), .B(n1281), .ZN(G39) );
NAND3_X1 U926 ( .A1(n1094), .A2(n1249), .A3(n1246), .ZN(n1281) );
XNOR2_X1 U927 ( .A(G134), .B(n1282), .ZN(G36) );
NAND2_X1 U928 ( .A1(n1246), .A2(n1247), .ZN(n1282) );
XNOR2_X1 U929 ( .A(G131), .B(n1233), .ZN(G33) );
NAND3_X1 U930 ( .A1(n1104), .A2(n1275), .A3(n1246), .ZN(n1233) );
AND2_X1 U931 ( .A1(n1274), .A2(n1093), .ZN(n1246) );
INV_X1 U932 ( .A(n1243), .ZN(n1093) );
NAND2_X1 U933 ( .A1(n1109), .A2(n1283), .ZN(n1243) );
XNOR2_X1 U934 ( .A(G128), .B(n1232), .ZN(G30) );
NAND4_X1 U935 ( .A1(n1274), .A2(n1073), .A3(n1251), .A4(n1249), .ZN(n1232) );
INV_X1 U936 ( .A(n1116), .ZN(n1073) );
AND3_X1 U937 ( .A1(n1244), .A2(n1091), .A3(n1245), .ZN(n1274) );
XNOR2_X1 U938 ( .A(n1201), .B(n1259), .ZN(G3) );
NOR3_X1 U939 ( .A1(n1114), .A2(n1265), .A3(n1284), .ZN(n1259) );
XNOR2_X1 U940 ( .A(G125), .B(n1231), .ZN(G27) );
NAND4_X1 U941 ( .A1(n1280), .A2(n1244), .A3(n1251), .A4(n1285), .ZN(n1231) );
AND2_X1 U942 ( .A1(n1086), .A2(n1104), .ZN(n1285) );
NAND2_X1 U943 ( .A1(n1286), .A2(n1287), .ZN(n1244) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1092), .A4(n1133), .ZN(n1287) );
INV_X1 U945 ( .A(G900), .ZN(n1133) );
XNOR2_X1 U946 ( .A(G122), .B(n1256), .ZN(G24) );
NAND4_X1 U947 ( .A1(n1288), .A2(n1098), .A3(n1289), .A4(n1120), .ZN(n1256) );
XNOR2_X1 U948 ( .A(G119), .B(n1255), .ZN(G21) );
NAND3_X1 U949 ( .A1(n1288), .A2(n1249), .A3(n1094), .ZN(n1255) );
INV_X1 U950 ( .A(n1284), .ZN(n1094) );
NAND2_X1 U951 ( .A1(n1290), .A2(n1291), .ZN(n1249) );
NAND2_X1 U952 ( .A1(n1275), .A2(n1292), .ZN(n1291) );
NAND3_X1 U953 ( .A1(n1293), .A2(n1122), .A3(KEYINPUT23), .ZN(n1290) );
XOR2_X1 U954 ( .A(n1261), .B(n1294), .Z(G18) );
XOR2_X1 U955 ( .A(KEYINPUT6), .B(G116), .Z(n1294) );
AND2_X1 U956 ( .A1(n1247), .A2(n1288), .ZN(n1261) );
NOR2_X1 U957 ( .A1(n1114), .A2(n1116), .ZN(n1247) );
NAND2_X1 U958 ( .A1(n1295), .A2(n1120), .ZN(n1116) );
XOR2_X1 U959 ( .A(G113), .B(n1260), .Z(G15) );
AND3_X1 U960 ( .A1(n1288), .A2(n1275), .A3(n1104), .ZN(n1260) );
NOR2_X1 U961 ( .A1(n1120), .A2(n1278), .ZN(n1104) );
INV_X1 U962 ( .A(n1289), .ZN(n1278) );
XNOR2_X1 U963 ( .A(n1295), .B(KEYINPUT39), .ZN(n1289) );
INV_X1 U964 ( .A(n1114), .ZN(n1275) );
NAND2_X1 U965 ( .A1(n1296), .A2(n1293), .ZN(n1114) );
AND3_X1 U966 ( .A1(n1251), .A2(n1297), .A3(n1086), .ZN(n1288) );
NOR2_X1 U967 ( .A1(n1245), .A2(n1242), .ZN(n1086) );
INV_X1 U968 ( .A(n1091), .ZN(n1242) );
NAND2_X1 U969 ( .A1(n1298), .A2(n1299), .ZN(G12) );
NAND2_X1 U970 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U971 ( .A(n1302), .B(KEYINPUT32), .Z(n1298) );
NAND2_X1 U972 ( .A1(G110), .A2(n1258), .ZN(n1302) );
INV_X1 U973 ( .A(n1300), .ZN(n1258) );
NOR3_X1 U974 ( .A1(n1265), .A2(n1113), .A3(n1284), .ZN(n1300) );
NAND2_X1 U975 ( .A1(n1277), .A2(n1295), .ZN(n1284) );
XOR2_X1 U976 ( .A(n1125), .B(G475), .Z(n1295) );
NAND2_X1 U977 ( .A1(n1182), .A2(n1266), .ZN(n1125) );
XOR2_X1 U978 ( .A(n1303), .B(n1304), .Z(n1182) );
NOR2_X1 U979 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U980 ( .A(KEYINPUT28), .B(n1307), .Z(n1306) );
NOR2_X1 U981 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
AND2_X1 U982 ( .A1(n1309), .A2(n1308), .ZN(n1305) );
XOR2_X1 U983 ( .A(n1310), .B(n1148), .Z(n1308) );
XOR2_X1 U984 ( .A(n1311), .B(G143), .Z(n1310) );
NAND2_X1 U985 ( .A1(G214), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U986 ( .A(n1313), .B(n1314), .ZN(n1309) );
XNOR2_X1 U987 ( .A(n1272), .B(G125), .ZN(n1314) );
NAND2_X1 U988 ( .A1(KEYINPUT59), .A2(n1315), .ZN(n1313) );
XOR2_X1 U989 ( .A(KEYINPUT46), .B(G140), .Z(n1315) );
NAND3_X1 U990 ( .A1(n1316), .A2(n1317), .A3(KEYINPUT33), .ZN(n1303) );
OR3_X1 U991 ( .A1(n1318), .A2(G104), .A3(KEYINPUT11), .ZN(n1317) );
NAND2_X1 U992 ( .A1(n1319), .A2(KEYINPUT11), .ZN(n1316) );
XNOR2_X1 U993 ( .A(G104), .B(n1320), .ZN(n1319) );
NAND2_X1 U994 ( .A1(KEYINPUT44), .A2(n1318), .ZN(n1320) );
XNOR2_X1 U995 ( .A(G113), .B(n1321), .ZN(n1318) );
INV_X1 U996 ( .A(n1120), .ZN(n1277) );
XNOR2_X1 U997 ( .A(n1322), .B(G478), .ZN(n1120) );
NAND2_X1 U998 ( .A1(n1172), .A2(n1266), .ZN(n1322) );
XNOR2_X1 U999 ( .A(n1323), .B(n1324), .ZN(n1172) );
XOR2_X1 U1000 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1001 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1002 ( .A1(G217), .A2(n1329), .ZN(n1328) );
NAND2_X1 U1003 ( .A1(KEYINPUT41), .A2(n1330), .ZN(n1327) );
XOR2_X1 U1004 ( .A(n1331), .B(n1332), .Z(n1323) );
XNOR2_X1 U1005 ( .A(KEYINPUT62), .B(n1333), .ZN(n1332) );
NAND2_X1 U1006 ( .A1(n1334), .A2(n1335), .ZN(n1331) );
NAND2_X1 U1007 ( .A1(n1336), .A2(n1321), .ZN(n1335) );
XOR2_X1 U1008 ( .A(KEYINPUT60), .B(n1337), .Z(n1334) );
NOR2_X1 U1009 ( .A1(n1338), .A2(n1321), .ZN(n1337) );
XNOR2_X1 U1010 ( .A(n1336), .B(KEYINPUT48), .ZN(n1338) );
XOR2_X1 U1011 ( .A(G116), .B(KEYINPUT31), .Z(n1336) );
INV_X1 U1012 ( .A(n1280), .ZN(n1113) );
NAND2_X1 U1013 ( .A1(n1339), .A2(n1340), .ZN(n1280) );
NAND2_X1 U1014 ( .A1(n1098), .A2(n1292), .ZN(n1340) );
NOR2_X1 U1015 ( .A1(n1122), .A2(n1293), .ZN(n1098) );
OR3_X1 U1016 ( .A1(n1296), .A2(n1293), .A3(n1292), .ZN(n1339) );
INV_X1 U1017 ( .A(KEYINPUT23), .ZN(n1292) );
XNOR2_X1 U1018 ( .A(n1123), .B(n1341), .ZN(n1293) );
XOR2_X1 U1019 ( .A(KEYINPUT54), .B(G472), .Z(n1341) );
NAND2_X1 U1020 ( .A1(n1342), .A2(n1266), .ZN(n1123) );
XOR2_X1 U1021 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1022 ( .A(KEYINPUT43), .B(n1202), .ZN(n1344) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1312), .ZN(n1202) );
NOR2_X1 U1024 ( .A1(G953), .A2(G237), .ZN(n1312) );
XOR2_X1 U1025 ( .A(n1345), .B(n1204), .Z(n1343) );
XNOR2_X1 U1026 ( .A(n1346), .B(n1347), .ZN(n1204) );
XNOR2_X1 U1027 ( .A(n1213), .B(n1348), .ZN(n1347) );
INV_X1 U1028 ( .A(n1271), .ZN(n1348) );
INV_X1 U1029 ( .A(n1122), .ZN(n1296) );
XOR2_X1 U1030 ( .A(n1349), .B(n1169), .Z(n1122) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1350), .ZN(n1169) );
OR2_X1 U1032 ( .A1(n1168), .A2(G902), .ZN(n1349) );
XNOR2_X1 U1033 ( .A(n1351), .B(n1352), .ZN(n1168) );
XOR2_X1 U1034 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1035 ( .A(n1355), .B(n1356), .ZN(n1354) );
NOR2_X1 U1036 ( .A1(KEYINPUT50), .A2(n1357), .ZN(n1356) );
XOR2_X1 U1037 ( .A(G140), .B(G125), .Z(n1357) );
NOR2_X1 U1038 ( .A1(KEYINPUT8), .A2(n1358), .ZN(n1355) );
XNOR2_X1 U1039 ( .A(G128), .B(n1359), .ZN(n1358) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1329), .ZN(n1353) );
AND2_X1 U1041 ( .A1(G234), .A2(n1132), .ZN(n1329) );
XNOR2_X1 U1042 ( .A(G110), .B(n1360), .ZN(n1351) );
XNOR2_X1 U1043 ( .A(n1272), .B(G137), .ZN(n1360) );
NAND4_X1 U1044 ( .A1(n1251), .A2(n1245), .A3(n1297), .A4(n1091), .ZN(n1265) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1350), .ZN(n1091) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1266), .ZN(n1350) );
NAND2_X1 U1047 ( .A1(n1286), .A2(n1361), .ZN(n1297) );
NAND4_X1 U1048 ( .A1(G953), .A2(G902), .A3(n1092), .A4(n1161), .ZN(n1361) );
INV_X1 U1049 ( .A(G898), .ZN(n1161) );
NAND3_X1 U1050 ( .A1(n1092), .A2(n1132), .A3(G952), .ZN(n1286) );
NAND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1092) );
XNOR2_X1 U1052 ( .A(n1362), .B(G469), .ZN(n1245) );
NAND2_X1 U1053 ( .A1(n1363), .A2(n1266), .ZN(n1362) );
XOR2_X1 U1054 ( .A(n1364), .B(n1365), .Z(n1363) );
XNOR2_X1 U1055 ( .A(n1213), .B(n1206), .ZN(n1365) );
XOR2_X1 U1056 ( .A(n1366), .B(n1367), .Z(n1206) );
XNOR2_X1 U1057 ( .A(G140), .B(n1301), .ZN(n1367) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1132), .ZN(n1366) );
XNOR2_X1 U1059 ( .A(n1368), .B(n1148), .ZN(n1213) );
XOR2_X1 U1060 ( .A(G131), .B(KEYINPUT29), .Z(n1148) );
NAND2_X1 U1061 ( .A1(KEYINPUT49), .A2(n1369), .ZN(n1368) );
XNOR2_X1 U1062 ( .A(n1144), .B(n1146), .ZN(n1369) );
XNOR2_X1 U1063 ( .A(n1330), .B(KEYINPUT55), .ZN(n1146) );
INV_X1 U1064 ( .A(G134), .ZN(n1330) );
INV_X1 U1065 ( .A(G137), .ZN(n1144) );
XOR2_X1 U1066 ( .A(n1370), .B(n1218), .Z(n1364) );
AND2_X1 U1067 ( .A1(n1371), .A2(n1372), .ZN(n1218) );
NAND2_X1 U1068 ( .A1(n1373), .A2(n1201), .ZN(n1372) );
XOR2_X1 U1069 ( .A(KEYINPUT51), .B(n1374), .Z(n1371) );
NOR2_X1 U1070 ( .A1(n1373), .A2(n1201), .ZN(n1374) );
INV_X1 U1071 ( .A(G101), .ZN(n1201) );
XNOR2_X1 U1072 ( .A(G104), .B(G107), .ZN(n1373) );
NAND2_X1 U1073 ( .A1(KEYINPUT42), .A2(n1147), .ZN(n1370) );
XOR2_X1 U1074 ( .A(G146), .B(n1325), .Z(n1147) );
XOR2_X1 U1075 ( .A(G128), .B(G143), .Z(n1325) );
NOR2_X1 U1076 ( .A1(n1109), .A2(n1108), .ZN(n1251) );
INV_X1 U1077 ( .A(n1283), .ZN(n1108) );
NAND2_X1 U1078 ( .A1(n1375), .A2(n1376), .ZN(n1283) );
XNOR2_X1 U1079 ( .A(G214), .B(KEYINPUT58), .ZN(n1375) );
XNOR2_X1 U1080 ( .A(n1377), .B(n1224), .ZN(n1109) );
NAND2_X1 U1081 ( .A1(G210), .A2(n1376), .ZN(n1224) );
NAND2_X1 U1082 ( .A1(n1378), .A2(n1266), .ZN(n1376) );
INV_X1 U1083 ( .A(G237), .ZN(n1378) );
NAND2_X1 U1084 ( .A1(n1379), .A2(n1266), .ZN(n1377) );
INV_X1 U1085 ( .A(G902), .ZN(n1266) );
XNOR2_X1 U1086 ( .A(n1159), .B(n1380), .ZN(n1379) );
NOR2_X1 U1087 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
NOR2_X1 U1088 ( .A1(KEYINPUT40), .A2(n1383), .ZN(n1382) );
AND2_X1 U1089 ( .A1(KEYINPUT38), .A2(n1383), .ZN(n1381) );
AND2_X1 U1090 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
OR2_X1 U1091 ( .A1(n1386), .A2(n1270), .ZN(n1385) );
XOR2_X1 U1092 ( .A(n1387), .B(KEYINPUT63), .Z(n1384) );
NAND2_X1 U1093 ( .A1(n1270), .A2(n1386), .ZN(n1387) );
XOR2_X1 U1094 ( .A(n1271), .B(n1388), .Z(n1386) );
NOR2_X1 U1095 ( .A1(KEYINPUT20), .A2(G125), .ZN(n1388) );
XOR2_X1 U1096 ( .A(G128), .B(n1389), .Z(n1271) );
NOR2_X1 U1097 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
AND3_X1 U1098 ( .A1(n1392), .A2(n1272), .A3(G143), .ZN(n1391) );
NOR2_X1 U1099 ( .A1(n1393), .A2(n1392), .ZN(n1390) );
INV_X1 U1100 ( .A(KEYINPUT16), .ZN(n1392) );
XNOR2_X1 U1101 ( .A(n1272), .B(G143), .ZN(n1393) );
INV_X1 U1102 ( .A(G146), .ZN(n1272) );
AND2_X1 U1103 ( .A1(G224), .A2(n1132), .ZN(n1270) );
INV_X1 U1104 ( .A(G953), .ZN(n1132) );
XNOR2_X1 U1105 ( .A(n1394), .B(n1395), .ZN(n1159) );
XOR2_X1 U1106 ( .A(n1345), .B(n1396), .Z(n1395) );
XOR2_X1 U1107 ( .A(n1397), .B(n1321), .Z(n1396) );
XOR2_X1 U1108 ( .A(G122), .B(KEYINPUT19), .Z(n1321) );
NAND2_X1 U1109 ( .A1(KEYINPUT56), .A2(n1333), .ZN(n1397) );
INV_X1 U1110 ( .A(G107), .ZN(n1333) );
XNOR2_X1 U1111 ( .A(G101), .B(G113), .ZN(n1345) );
XOR2_X1 U1112 ( .A(n1398), .B(n1399), .Z(n1394) );
XNOR2_X1 U1113 ( .A(n1301), .B(G104), .ZN(n1399) );
INV_X1 U1114 ( .A(G110), .ZN(n1301) );
NAND2_X1 U1115 ( .A1(KEYINPUT4), .A2(n1346), .ZN(n1398) );
XNOR2_X1 U1116 ( .A(G116), .B(n1359), .ZN(n1346) );
XOR2_X1 U1117 ( .A(G119), .B(KEYINPUT57), .Z(n1359) );
endmodule


