//Key = 0000100000110101010001110110011110101100011100110000001001001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353;

XNOR2_X1 U754 ( .A(G107), .B(n1027), .ZN(G9) );
NAND3_X1 U755 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(G75) );
NAND2_X1 U756 ( .A1(G952), .A2(n1031), .ZN(n1030) );
NAND3_X1 U757 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR3_X1 U758 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U759 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U760 ( .A(n1040), .B(KEYINPUT49), .Z(n1038) );
NOR3_X1 U761 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1036) );
OR2_X1 U762 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
NOR2_X1 U763 ( .A1(n1045), .A2(n1046), .ZN(n1035) );
INV_X1 U764 ( .A(n1047), .ZN(n1046) );
NOR3_X1 U765 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1045) );
NOR2_X1 U766 ( .A1(n1051), .A2(n1043), .ZN(n1050) );
NOR3_X1 U767 ( .A1(n1044), .A2(n1052), .A3(n1053), .ZN(n1049) );
NOR2_X1 U768 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U769 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U770 ( .A(n1058), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
XOR2_X1 U772 ( .A(KEYINPUT18), .B(n1061), .Z(n1048) );
NOR3_X1 U773 ( .A1(n1062), .A2(n1043), .A3(n1063), .ZN(n1061) );
NAND3_X1 U774 ( .A1(n1058), .A2(n1064), .A3(n1065), .ZN(n1043) );
INV_X1 U775 ( .A(n1053), .ZN(n1064) );
XOR2_X1 U776 ( .A(n1066), .B(KEYINPUT15), .Z(n1053) );
NAND4_X1 U777 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1028) );
NOR4_X1 U778 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
XOR2_X1 U779 ( .A(n1075), .B(KEYINPUT4), .Z(n1071) );
AND2_X1 U780 ( .A1(n1062), .A2(n1041), .ZN(n1069) );
XOR2_X1 U781 ( .A(n1076), .B(n1077), .Z(n1068) );
NOR2_X1 U782 ( .A1(G478), .A2(KEYINPUT7), .ZN(n1077) );
XOR2_X1 U783 ( .A(n1078), .B(n1079), .Z(n1067) );
NOR2_X1 U784 ( .A1(n1080), .A2(KEYINPUT2), .ZN(n1078) );
XOR2_X1 U785 ( .A(n1081), .B(n1082), .Z(G72) );
XOR2_X1 U786 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U787 ( .A1(G953), .A2(n1085), .ZN(n1084) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1085) );
NAND3_X1 U789 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1083) );
XOR2_X1 U790 ( .A(n1089), .B(KEYINPUT58), .Z(n1088) );
NAND2_X1 U791 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U792 ( .A(n1092), .ZN(n1091) );
XOR2_X1 U793 ( .A(KEYINPUT25), .B(n1093), .Z(n1090) );
NAND2_X1 U794 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
XNOR2_X1 U795 ( .A(n1094), .B(n1095), .ZN(n1093) );
XOR2_X1 U796 ( .A(KEYINPUT1), .B(n1096), .Z(n1095) );
XOR2_X1 U797 ( .A(KEYINPUT43), .B(KEYINPUT28), .Z(n1096) );
XOR2_X1 U798 ( .A(n1097), .B(n1098), .Z(n1094) );
XOR2_X1 U799 ( .A(n1099), .B(G137), .Z(n1097) );
XOR2_X1 U800 ( .A(n1100), .B(n1101), .Z(n1092) );
NOR2_X1 U801 ( .A1(G140), .A2(KEYINPUT59), .ZN(n1101) );
NAND2_X1 U802 ( .A1(G953), .A2(n1102), .ZN(n1086) );
NOR2_X1 U803 ( .A1(n1033), .A2(G953), .ZN(n1081) );
XOR2_X1 U804 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U805 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U806 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U808 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U809 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U810 ( .A(n1111), .B(n1112), .Z(n1108) );
XOR2_X1 U811 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U812 ( .A1(KEYINPUT44), .A2(n1115), .ZN(n1114) );
XOR2_X1 U813 ( .A(G122), .B(G110), .Z(n1115) );
NAND2_X1 U814 ( .A1(KEYINPUT13), .A2(n1116), .ZN(n1111) );
XNOR2_X1 U815 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U816 ( .A1(n1032), .A2(G953), .ZN(n1103) );
NOR2_X1 U817 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XNOR2_X1 U818 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U819 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U820 ( .A1(n1119), .A2(n1125), .ZN(G63) );
NOR3_X1 U821 ( .A1(n1076), .A2(n1126), .A3(n1127), .ZN(n1125) );
NOR3_X1 U822 ( .A1(n1128), .A2(n1129), .A3(n1124), .ZN(n1127) );
INV_X1 U823 ( .A(n1130), .ZN(n1128) );
NOR2_X1 U824 ( .A1(n1131), .A2(n1130), .ZN(n1126) );
NOR2_X1 U825 ( .A1(n1132), .A2(n1129), .ZN(n1131) );
NOR2_X1 U826 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR3_X1 U827 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(G60) );
NOR3_X1 U828 ( .A1(n1138), .A2(n1029), .A3(n1139), .ZN(n1137) );
AND2_X1 U829 ( .A1(n1138), .A2(n1119), .ZN(n1136) );
INV_X1 U830 ( .A(KEYINPUT9), .ZN(n1138) );
XOR2_X1 U831 ( .A(n1140), .B(n1141), .Z(n1135) );
NOR2_X1 U832 ( .A1(n1142), .A2(n1124), .ZN(n1140) );
XNOR2_X1 U833 ( .A(G475), .B(KEYINPUT27), .ZN(n1142) );
XNOR2_X1 U834 ( .A(G104), .B(n1143), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1119), .A2(n1144), .ZN(G57) );
XOR2_X1 U836 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U837 ( .A1(n1147), .A2(n1124), .ZN(n1146) );
INV_X1 U838 ( .A(G472), .ZN(n1147) );
NOR2_X1 U839 ( .A1(n1119), .A2(n1148), .ZN(G54) );
XOR2_X1 U840 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U841 ( .A1(n1151), .A2(n1124), .ZN(n1150) );
INV_X1 U842 ( .A(G469), .ZN(n1151) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
XOR2_X1 U844 ( .A(KEYINPUT56), .B(n1154), .Z(n1153) );
NOR2_X1 U845 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
INV_X1 U846 ( .A(n1157), .ZN(n1156) );
NOR2_X1 U847 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
XNOR2_X1 U848 ( .A(n1155), .B(KEYINPUT53), .ZN(n1158) );
XOR2_X1 U849 ( .A(n1159), .B(n1160), .Z(n1155) );
XOR2_X1 U850 ( .A(n1099), .B(n1161), .Z(n1159) );
XNOR2_X1 U851 ( .A(n1162), .B(n1163), .ZN(n1157) );
XOR2_X1 U852 ( .A(n1164), .B(KEYINPUT52), .Z(n1162) );
NAND2_X1 U853 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U854 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U855 ( .A(n1169), .B(KEYINPUT33), .Z(n1165) );
NAND2_X1 U856 ( .A1(n1170), .A2(G110), .ZN(n1169) );
XOR2_X1 U857 ( .A(n1167), .B(KEYINPUT29), .Z(n1170) );
XNOR2_X1 U858 ( .A(G140), .B(KEYINPUT11), .ZN(n1167) );
NOR2_X1 U859 ( .A1(n1119), .A2(n1171), .ZN(G51) );
XOR2_X1 U860 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND3_X1 U861 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1172) );
NAND2_X1 U862 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
INV_X1 U863 ( .A(n1179), .ZN(n1178) );
NAND3_X1 U864 ( .A1(n1179), .A2(n1180), .A3(G125), .ZN(n1175) );
NAND2_X1 U865 ( .A1(n1181), .A2(n1100), .ZN(n1174) );
XOR2_X1 U866 ( .A(n1179), .B(n1180), .Z(n1181) );
NOR2_X1 U867 ( .A1(n1124), .A2(n1182), .ZN(n1179) );
NAND2_X1 U868 ( .A1(G902), .A2(n1183), .ZN(n1124) );
NAND2_X1 U869 ( .A1(n1032), .A2(n1033), .ZN(n1183) );
INV_X1 U870 ( .A(n1133), .ZN(n1033) );
NAND4_X1 U871 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1133) );
AND4_X1 U872 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U873 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
NOR2_X1 U874 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U875 ( .A1(n1196), .A2(n1197), .ZN(n1192) );
NOR2_X1 U876 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
XOR2_X1 U877 ( .A(KEYINPUT35), .B(n1200), .Z(n1199) );
NAND3_X1 U878 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1185) );
INV_X1 U879 ( .A(KEYINPUT31), .ZN(n1203) );
NAND2_X1 U880 ( .A1(n1204), .A2(KEYINPUT31), .ZN(n1184) );
INV_X1 U881 ( .A(n1134), .ZN(n1032) );
NAND4_X1 U882 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1134) );
AND3_X1 U883 ( .A1(n1209), .A2(n1143), .A3(n1027), .ZN(n1208) );
NAND3_X1 U884 ( .A1(n1058), .A2(n1210), .A3(n1060), .ZN(n1027) );
NAND3_X1 U885 ( .A1(n1058), .A2(n1210), .A3(n1059), .ZN(n1143) );
NAND2_X1 U886 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
NAND2_X1 U887 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U888 ( .A1(n1215), .A2(n1058), .ZN(n1214) );
XNOR2_X1 U889 ( .A(n1216), .B(KEYINPUT57), .ZN(n1215) );
NAND2_X1 U890 ( .A1(n1217), .A2(n1200), .ZN(n1213) );
XOR2_X1 U891 ( .A(n1218), .B(KEYINPUT62), .Z(n1217) );
NAND2_X1 U892 ( .A1(n1054), .A2(n1210), .ZN(n1205) );
AND2_X1 U893 ( .A1(n1065), .A2(n1219), .ZN(n1054) );
NAND2_X1 U894 ( .A1(n1194), .A2(n1220), .ZN(n1219) );
NOR2_X1 U895 ( .A1(n1029), .A2(G952), .ZN(n1119) );
XOR2_X1 U896 ( .A(n1221), .B(n1191), .Z(G48) );
NAND3_X1 U897 ( .A1(n1059), .A2(n1222), .A3(n1223), .ZN(n1191) );
XOR2_X1 U898 ( .A(G143), .B(n1224), .Z(G45) );
NOR2_X1 U899 ( .A1(n1195), .A2(n1225), .ZN(n1224) );
XOR2_X1 U900 ( .A(KEYINPUT30), .B(n1200), .Z(n1225) );
NAND3_X1 U901 ( .A1(n1216), .A2(n1222), .A3(n1226), .ZN(n1195) );
XOR2_X1 U902 ( .A(G140), .B(n1227), .Z(G42) );
NOR2_X1 U903 ( .A1(n1197), .A2(n1220), .ZN(n1227) );
XOR2_X1 U904 ( .A(n1228), .B(n1190), .Z(G39) );
NAND3_X1 U905 ( .A1(n1223), .A2(n1065), .A3(n1047), .ZN(n1190) );
XOR2_X1 U906 ( .A(n1229), .B(n1189), .Z(G36) );
NAND4_X1 U907 ( .A1(n1047), .A2(n1226), .A3(n1200), .A4(n1060), .ZN(n1189) );
XOR2_X1 U908 ( .A(G131), .B(n1230), .Z(G33) );
NOR2_X1 U909 ( .A1(n1194), .A2(n1197), .ZN(n1230) );
NAND3_X1 U910 ( .A1(n1226), .A2(n1059), .A3(n1047), .ZN(n1197) );
NOR2_X1 U911 ( .A1(n1042), .A2(n1231), .ZN(n1047) );
XOR2_X1 U912 ( .A(KEYINPUT21), .B(n1041), .Z(n1231) );
INV_X1 U913 ( .A(n1218), .ZN(n1059) );
INV_X1 U914 ( .A(n1200), .ZN(n1194) );
XNOR2_X1 U915 ( .A(G128), .B(n1188), .ZN(G30) );
NAND3_X1 U916 ( .A1(n1060), .A2(n1222), .A3(n1223), .ZN(n1188) );
AND3_X1 U917 ( .A1(n1074), .A2(n1232), .A3(n1226), .ZN(n1223) );
NOR2_X1 U918 ( .A1(n1202), .A2(n1051), .ZN(n1226) );
XOR2_X1 U919 ( .A(n1233), .B(n1234), .Z(G3) );
NAND3_X1 U920 ( .A1(n1210), .A2(n1235), .A3(n1200), .ZN(n1234) );
XOR2_X1 U921 ( .A(KEYINPUT19), .B(n1065), .Z(n1235) );
NOR2_X1 U922 ( .A1(n1051), .A2(n1236), .ZN(n1210) );
XOR2_X1 U923 ( .A(G125), .B(n1204), .Z(G27) );
NOR2_X1 U924 ( .A1(n1237), .A2(n1202), .ZN(n1204) );
NAND3_X1 U925 ( .A1(n1238), .A2(n1239), .A3(n1066), .ZN(n1202) );
NAND2_X1 U926 ( .A1(G953), .A2(n1240), .ZN(n1238) );
NAND2_X1 U927 ( .A1(G902), .A2(n1102), .ZN(n1240) );
INV_X1 U928 ( .A(G900), .ZN(n1102) );
INV_X1 U929 ( .A(n1201), .ZN(n1237) );
NOR4_X1 U930 ( .A1(n1220), .A2(n1044), .A3(n1218), .A4(n1039), .ZN(n1201) );
XOR2_X1 U931 ( .A(n1241), .B(n1242), .Z(G24) );
NAND3_X1 U932 ( .A1(n1211), .A2(n1058), .A3(n1216), .ZN(n1242) );
AND2_X1 U933 ( .A1(n1072), .A2(n1243), .ZN(n1216) );
NOR2_X1 U934 ( .A1(n1232), .A2(n1074), .ZN(n1058) );
XOR2_X1 U935 ( .A(n1244), .B(n1206), .Z(G21) );
NAND4_X1 U936 ( .A1(n1065), .A2(n1211), .A3(n1074), .A4(n1232), .ZN(n1206) );
INV_X1 U937 ( .A(n1075), .ZN(n1232) );
XNOR2_X1 U938 ( .A(n1245), .B(n1209), .ZN(G18) );
NAND2_X1 U939 ( .A1(n1246), .A2(n1060), .ZN(n1209) );
NOR2_X1 U940 ( .A1(n1072), .A2(n1247), .ZN(n1060) );
INV_X1 U941 ( .A(n1248), .ZN(n1246) );
XOR2_X1 U942 ( .A(n1249), .B(KEYINPUT23), .Z(n1245) );
XOR2_X1 U943 ( .A(G113), .B(n1250), .Z(G15) );
NOR2_X1 U944 ( .A1(n1218), .A2(n1248), .ZN(n1250) );
NAND2_X1 U945 ( .A1(n1211), .A2(n1200), .ZN(n1248) );
NOR2_X1 U946 ( .A1(n1074), .A2(n1075), .ZN(n1200) );
NOR2_X1 U947 ( .A1(n1044), .A2(n1236), .ZN(n1211) );
NAND2_X1 U948 ( .A1(n1251), .A2(n1062), .ZN(n1044) );
NAND2_X1 U949 ( .A1(n1247), .A2(n1072), .ZN(n1218) );
INV_X1 U950 ( .A(n1243), .ZN(n1247) );
XOR2_X1 U951 ( .A(n1252), .B(n1253), .Z(G12) );
NAND2_X1 U952 ( .A1(KEYINPUT36), .A2(G110), .ZN(n1253) );
NAND4_X1 U953 ( .A1(n1254), .A2(n1198), .A3(n1065), .A4(n1255), .ZN(n1252) );
INV_X1 U954 ( .A(n1236), .ZN(n1255) );
NAND4_X1 U955 ( .A1(n1222), .A2(n1066), .A3(n1256), .A4(n1239), .ZN(n1236) );
NAND2_X1 U956 ( .A1(n1139), .A2(n1029), .ZN(n1239) );
INV_X1 U957 ( .A(G952), .ZN(n1139) );
NAND2_X1 U958 ( .A1(G953), .A2(n1257), .ZN(n1256) );
NAND2_X1 U959 ( .A1(G902), .A2(n1110), .ZN(n1257) );
INV_X1 U960 ( .A(G898), .ZN(n1110) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1066) );
INV_X1 U962 ( .A(n1039), .ZN(n1222) );
NAND2_X1 U963 ( .A1(n1042), .A2(n1041), .ZN(n1039) );
NAND2_X1 U964 ( .A1(n1258), .A2(G214), .ZN(n1041) );
XOR2_X1 U965 ( .A(n1259), .B(KEYINPUT8), .Z(n1258) );
XOR2_X1 U966 ( .A(n1073), .B(KEYINPUT0), .Z(n1042) );
XOR2_X1 U967 ( .A(n1260), .B(n1182), .Z(n1073) );
NAND2_X1 U968 ( .A1(G210), .A2(n1259), .ZN(n1182) );
NAND2_X1 U969 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
INV_X1 U970 ( .A(G237), .ZN(n1262) );
NAND2_X1 U971 ( .A1(n1263), .A2(n1261), .ZN(n1260) );
XOR2_X1 U972 ( .A(n1173), .B(n1264), .Z(n1263) );
NOR2_X1 U973 ( .A1(n1177), .A2(n1265), .ZN(n1264) );
XOR2_X1 U974 ( .A(n1266), .B(KEYINPUT26), .Z(n1265) );
NAND2_X1 U975 ( .A1(n1267), .A2(n1100), .ZN(n1266) );
XOR2_X1 U976 ( .A(KEYINPUT55), .B(n1180), .Z(n1267) );
NOR2_X1 U977 ( .A1(n1180), .A2(n1100), .ZN(n1177) );
XOR2_X1 U978 ( .A(n1268), .B(n1269), .Z(n1173) );
XOR2_X1 U979 ( .A(n1117), .B(n1270), .Z(n1269) );
NAND3_X1 U980 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1117) );
NAND2_X1 U981 ( .A1(KEYINPUT48), .A2(G119), .ZN(n1273) );
NAND3_X1 U982 ( .A1(n1244), .A2(n1274), .A3(G116), .ZN(n1272) );
NAND2_X1 U983 ( .A1(n1275), .A2(n1249), .ZN(n1271) );
NAND2_X1 U984 ( .A1(n1276), .A2(n1274), .ZN(n1275) );
INV_X1 U985 ( .A(KEYINPUT48), .ZN(n1274) );
XOR2_X1 U986 ( .A(n1244), .B(KEYINPUT12), .Z(n1276) );
XOR2_X1 U987 ( .A(n1277), .B(n1278), .Z(n1268) );
NOR2_X1 U988 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U989 ( .A(G224), .B(KEYINPUT14), .ZN(n1280) );
XOR2_X1 U990 ( .A(n1113), .B(G110), .Z(n1277) );
NAND3_X1 U991 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1113) );
NAND2_X1 U992 ( .A1(KEYINPUT3), .A2(n1284), .ZN(n1283) );
OR3_X1 U993 ( .A1(n1285), .A2(KEYINPUT3), .A3(G101), .ZN(n1282) );
NAND2_X1 U994 ( .A1(G101), .A2(n1285), .ZN(n1281) );
NAND2_X1 U995 ( .A1(KEYINPUT37), .A2(n1286), .ZN(n1285) );
NOR2_X1 U996 ( .A1(n1243), .A2(n1072), .ZN(n1065) );
XNOR2_X1 U997 ( .A(n1287), .B(G475), .ZN(n1072) );
OR2_X1 U998 ( .A1(n1141), .A2(G902), .ZN(n1287) );
XNOR2_X1 U999 ( .A(n1288), .B(n1289), .ZN(n1141) );
XOR2_X1 U1000 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1001 ( .A(n1270), .B(n1292), .Z(n1291) );
NOR2_X1 U1002 ( .A1(KEYINPUT40), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1003 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1004 ( .A1(KEYINPUT16), .A2(G143), .ZN(n1295) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1296), .ZN(n1294) );
XOR2_X1 U1006 ( .A(n1241), .B(n1118), .Z(n1270) );
INV_X1 U1007 ( .A(G122), .ZN(n1241) );
XNOR2_X1 U1008 ( .A(G104), .B(n1297), .ZN(n1288) );
XOR2_X1 U1009 ( .A(G146), .B(G131), .Z(n1297) );
NAND2_X1 U1010 ( .A1(n1298), .A2(n1299), .ZN(n1243) );
NAND2_X1 U1011 ( .A1(n1076), .A2(n1129), .ZN(n1299) );
XOR2_X1 U1012 ( .A(KEYINPUT17), .B(n1300), .Z(n1298) );
NOR2_X1 U1013 ( .A1(n1076), .A2(n1129), .ZN(n1300) );
INV_X1 U1014 ( .A(G478), .ZN(n1129) );
NOR2_X1 U1015 ( .A1(n1130), .A2(G902), .ZN(n1076) );
XOR2_X1 U1016 ( .A(n1301), .B(n1302), .Z(n1130) );
NOR2_X1 U1017 ( .A1(KEYINPUT24), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1018 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U1019 ( .A(G107), .B(n1306), .Z(n1305) );
NOR2_X1 U1020 ( .A1(KEYINPUT6), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1021 ( .A(G134), .B(n1308), .Z(n1307) );
XOR2_X1 U1022 ( .A(G122), .B(G116), .Z(n1304) );
NAND3_X1 U1023 ( .A1(G217), .A2(n1309), .A3(G234), .ZN(n1301) );
INV_X1 U1024 ( .A(n1220), .ZN(n1198) );
NAND2_X1 U1025 ( .A1(n1075), .A2(n1074), .ZN(n1220) );
XOR2_X1 U1026 ( .A(n1310), .B(n1123), .Z(n1074) );
NAND2_X1 U1027 ( .A1(G217), .A2(n1311), .ZN(n1123) );
NAND2_X1 U1028 ( .A1(n1121), .A2(n1261), .ZN(n1310) );
XNOR2_X1 U1029 ( .A(n1312), .B(n1313), .ZN(n1121) );
XOR2_X1 U1030 ( .A(G137), .B(n1314), .Z(n1313) );
NOR2_X1 U1031 ( .A1(KEYINPUT5), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1032 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U1033 ( .A(n1318), .B(n1290), .Z(n1317) );
XOR2_X1 U1034 ( .A(G140), .B(n1100), .Z(n1290) );
INV_X1 U1035 ( .A(G125), .ZN(n1100) );
NAND2_X1 U1036 ( .A1(n1319), .A2(KEYINPUT41), .ZN(n1318) );
XOR2_X1 U1037 ( .A(n1221), .B(KEYINPUT61), .Z(n1319) );
XOR2_X1 U1038 ( .A(G110), .B(n1320), .Z(n1316) );
XOR2_X1 U1039 ( .A(G128), .B(G119), .Z(n1320) );
NAND3_X1 U1040 ( .A1(G234), .A2(n1321), .A3(G221), .ZN(n1312) );
XOR2_X1 U1041 ( .A(KEYINPUT50), .B(n1309), .Z(n1321) );
XOR2_X1 U1042 ( .A(n1322), .B(G472), .Z(n1075) );
NAND2_X1 U1043 ( .A1(n1323), .A2(n1261), .ZN(n1322) );
XOR2_X1 U1044 ( .A(n1145), .B(KEYINPUT10), .Z(n1323) );
XOR2_X1 U1045 ( .A(n1324), .B(n1325), .Z(n1145) );
XNOR2_X1 U1046 ( .A(n1180), .B(n1160), .ZN(n1325) );
XNOR2_X1 U1047 ( .A(n1221), .B(n1308), .ZN(n1180) );
XOR2_X1 U1048 ( .A(G128), .B(G143), .Z(n1308) );
XOR2_X1 U1049 ( .A(n1326), .B(n1327), .Z(n1324) );
AND2_X1 U1050 ( .A1(n1296), .A2(G210), .ZN(n1327) );
NOR2_X1 U1051 ( .A1(n1279), .A2(G237), .ZN(n1296) );
XOR2_X1 U1052 ( .A(n1328), .B(G101), .Z(n1326) );
NAND3_X1 U1053 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
OR2_X1 U1054 ( .A1(n1332), .A2(KEYINPUT32), .ZN(n1331) );
OR3_X1 U1055 ( .A1(n1333), .A2(n1334), .A3(n1118), .ZN(n1330) );
INV_X1 U1056 ( .A(KEYINPUT32), .ZN(n1333) );
NAND2_X1 U1057 ( .A1(n1118), .A2(n1334), .ZN(n1329) );
NAND2_X1 U1058 ( .A1(KEYINPUT47), .A2(n1332), .ZN(n1334) );
XOR2_X1 U1059 ( .A(n1249), .B(n1244), .Z(n1332) );
INV_X1 U1060 ( .A(G119), .ZN(n1244) );
INV_X1 U1061 ( .A(G116), .ZN(n1249) );
XOR2_X1 U1062 ( .A(G113), .B(KEYINPUT51), .Z(n1118) );
XOR2_X1 U1063 ( .A(n1051), .B(KEYINPUT42), .Z(n1254) );
NAND2_X1 U1064 ( .A1(n1063), .A2(n1062), .ZN(n1051) );
NAND2_X1 U1065 ( .A1(G221), .A2(n1311), .ZN(n1062) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1261), .ZN(n1311) );
INV_X1 U1067 ( .A(n1251), .ZN(n1063) );
XNOR2_X1 U1068 ( .A(n1080), .B(n1079), .ZN(n1251) );
XOR2_X1 U1069 ( .A(G469), .B(KEYINPUT45), .Z(n1079) );
AND2_X1 U1070 ( .A1(n1335), .A2(n1261), .ZN(n1080) );
INV_X1 U1071 ( .A(G902), .ZN(n1261) );
XOR2_X1 U1072 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1073 ( .A(n1163), .B(n1160), .Z(n1337) );
XOR2_X1 U1074 ( .A(n1338), .B(n1098), .Z(n1160) );
XNOR2_X1 U1075 ( .A(G131), .B(n1229), .ZN(n1098) );
INV_X1 U1076 ( .A(G134), .ZN(n1229) );
NAND2_X1 U1077 ( .A1(KEYINPUT46), .A2(n1228), .ZN(n1338) );
INV_X1 U1078 ( .A(G137), .ZN(n1228) );
NAND2_X1 U1079 ( .A1(G227), .A2(n1309), .ZN(n1163) );
INV_X1 U1080 ( .A(n1279), .ZN(n1309) );
XOR2_X1 U1081 ( .A(n1029), .B(KEYINPUT54), .Z(n1279) );
INV_X1 U1082 ( .A(G953), .ZN(n1029) );
XOR2_X1 U1083 ( .A(n1339), .B(n1340), .Z(n1336) );
XOR2_X1 U1084 ( .A(G140), .B(n1168), .Z(n1340) );
INV_X1 U1085 ( .A(G110), .ZN(n1168) );
NAND2_X1 U1086 ( .A1(KEYINPUT22), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1087 ( .A(n1161), .B(n1342), .Z(n1341) );
NOR2_X1 U1088 ( .A1(KEYINPUT39), .A2(n1099), .ZN(n1342) );
XNOR2_X1 U1089 ( .A(G128), .B(n1343), .ZN(n1099) );
NOR2_X1 U1090 ( .A1(n1344), .A2(KEYINPUT20), .ZN(n1343) );
NOR2_X1 U1091 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1092 ( .A(n1347), .B(KEYINPUT63), .Z(n1346) );
NAND2_X1 U1093 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1094 ( .A(n1221), .B(KEYINPUT34), .Z(n1348) );
INV_X1 U1095 ( .A(G146), .ZN(n1221) );
NOR2_X1 U1096 ( .A1(G146), .A2(n1349), .ZN(n1345) );
INV_X1 U1097 ( .A(G143), .ZN(n1349) );
AND3_X1 U1098 ( .A1(n1350), .A2(n1351), .A3(n1352), .ZN(n1161) );
NAND2_X1 U1099 ( .A1(KEYINPUT38), .A2(n1286), .ZN(n1352) );
OR3_X1 U1100 ( .A1(n1353), .A2(KEYINPUT38), .A3(n1233), .ZN(n1351) );
NAND2_X1 U1101 ( .A1(n1353), .A2(n1233), .ZN(n1350) );
INV_X1 U1102 ( .A(G101), .ZN(n1233) );
NAND2_X1 U1103 ( .A1(KEYINPUT60), .A2(n1284), .ZN(n1353) );
INV_X1 U1104 ( .A(n1286), .ZN(n1284) );
XOR2_X1 U1105 ( .A(G104), .B(G107), .Z(n1286) );
endmodule


