//Key = 1101111001010101111001001111000001111000001011011001001111100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337;

XOR2_X1 U750 ( .A(G107), .B(n1023), .Z(G9) );
NOR2_X1 U751 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR4_X1 U753 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1027) );
NOR4_X1 U754 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1030) );
NOR2_X1 U755 ( .A1(KEYINPUT41), .A2(n1037), .ZN(n1036) );
NOR2_X1 U756 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
NOR2_X1 U757 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U758 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
AND2_X1 U759 ( .A1(n1044), .A2(n1045), .ZN(n1034) );
NOR2_X1 U760 ( .A1(n1046), .A2(n1047), .ZN(n1029) );
NOR2_X1 U761 ( .A1(n1037), .A2(n1048), .ZN(n1047) );
INV_X1 U762 ( .A(KEYINPUT41), .ZN(n1048) );
NAND3_X1 U763 ( .A1(n1049), .A2(n1050), .A3(n1045), .ZN(n1037) );
NAND3_X1 U764 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1026) );
NAND4_X1 U765 ( .A1(n1046), .A2(n1045), .A3(n1054), .A4(n1055), .ZN(n1053) );
NAND4_X1 U766 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
NAND3_X1 U767 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
XOR2_X1 U768 ( .A(n1032), .B(KEYINPUT34), .Z(n1062) );
NAND2_X1 U769 ( .A1(n1063), .A2(n1064), .ZN(n1058) );
XOR2_X1 U770 ( .A(KEYINPUT20), .B(n1065), .Z(n1064) );
NAND2_X1 U771 ( .A1(n1065), .A2(n1066), .ZN(n1057) );
NAND2_X1 U772 ( .A1(n1067), .A2(n1068), .ZN(n1056) );
INV_X1 U773 ( .A(n1033), .ZN(n1046) );
NOR3_X1 U774 ( .A1(n1069), .A2(G953), .A3(G952), .ZN(n1024) );
INV_X1 U775 ( .A(n1051), .ZN(n1069) );
NAND4_X1 U776 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1051) );
NOR4_X1 U777 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U779 ( .A(KEYINPUT60), .B(n1080), .Z(n1076) );
NOR3_X1 U780 ( .A1(n1081), .A2(n1061), .A3(n1082), .ZN(n1072) );
AND2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XOR2_X1 U782 ( .A(n1085), .B(n1086), .Z(n1071) );
NAND2_X1 U783 ( .A1(KEYINPUT21), .A2(n1087), .ZN(n1086) );
XOR2_X1 U784 ( .A(KEYINPUT15), .B(n1088), .Z(n1070) );
NOR2_X1 U785 ( .A1(n1084), .A2(n1083), .ZN(n1088) );
XNOR2_X1 U786 ( .A(n1089), .B(KEYINPUT61), .ZN(n1083) );
XOR2_X1 U787 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND3_X1 U789 ( .A1(KEYINPUT18), .A2(n1094), .A3(G953), .ZN(n1093) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1094) );
NOR3_X1 U791 ( .A1(G953), .A2(KEYINPUT8), .A3(n1095), .ZN(n1092) );
NOR2_X1 U792 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(n1090) );
NAND2_X1 U794 ( .A1(G953), .A2(n1100), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(n1098) );
XOR2_X1 U796 ( .A(KEYINPUT3), .B(KEYINPUT19), .Z(n1102) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(n1101) );
NAND2_X1 U798 ( .A1(n1105), .A2(KEYINPUT24), .ZN(n1103) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U800 ( .A(G131), .B(n1108), .Z(n1107) );
NAND2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND3_X1 U802 ( .A1(G953), .A2(n1111), .A3(n1112), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
NAND2_X1 U804 ( .A1(G953), .A2(n1111), .ZN(n1114) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1111) );
XOR2_X1 U806 ( .A(n1112), .B(n1115), .Z(n1113) );
NOR2_X1 U807 ( .A1(n1023), .A2(n1116), .ZN(n1115) );
INV_X1 U808 ( .A(n1117), .ZN(n1023) );
AND2_X1 U809 ( .A1(KEYINPUT48), .A2(n1118), .ZN(n1112) );
NAND2_X1 U810 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U811 ( .A1(G953), .A2(n1121), .ZN(n1120) );
XOR2_X1 U812 ( .A(n1122), .B(n1123), .Z(n1119) );
XNOR2_X1 U813 ( .A(n1124), .B(n1125), .ZN(n1122) );
NOR2_X1 U814 ( .A1(KEYINPUT30), .A2(n1126), .ZN(n1125) );
NOR2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U818 ( .A1(n1127), .A2(n1133), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1084), .A2(n1134), .A3(n1135), .ZN(n1133) );
NOR3_X1 U820 ( .A1(n1136), .A2(n1089), .A3(n1132), .ZN(n1135) );
NOR2_X1 U821 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1089), .ZN(n1138) );
INV_X1 U823 ( .A(G478), .ZN(n1089) );
NOR2_X1 U824 ( .A1(n1127), .A2(n1140), .ZN(G60) );
XOR2_X1 U825 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1132), .ZN(n1141) );
INV_X1 U827 ( .A(G475), .ZN(n1143) );
XOR2_X1 U828 ( .A(G104), .B(n1144), .Z(G6) );
NOR2_X1 U829 ( .A1(n1127), .A2(n1145), .ZN(G57) );
XOR2_X1 U830 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U831 ( .A(n1148), .B(n1149), .ZN(n1147) );
NOR2_X1 U832 ( .A1(n1078), .A2(n1132), .ZN(n1148) );
INV_X1 U833 ( .A(G472), .ZN(n1078) );
XOR2_X1 U834 ( .A(n1150), .B(n1151), .Z(n1146) );
NOR2_X1 U835 ( .A1(KEYINPUT40), .A2(n1152), .ZN(n1151) );
NOR3_X1 U836 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1150) );
NOR2_X1 U837 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR3_X1 U838 ( .A1(n1158), .A2(KEYINPUT10), .A3(n1159), .ZN(n1154) );
INV_X1 U839 ( .A(n1157), .ZN(n1159) );
NOR2_X1 U840 ( .A1(KEYINPUT2), .A2(n1160), .ZN(n1157) );
AND2_X1 U841 ( .A1(n1160), .A2(KEYINPUT10), .ZN(n1153) );
INV_X1 U842 ( .A(n1161), .ZN(n1160) );
NOR2_X1 U843 ( .A1(n1127), .A2(n1162), .ZN(G54) );
XOR2_X1 U844 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U845 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U846 ( .A1(n1132), .A2(n1087), .ZN(n1165) );
INV_X1 U847 ( .A(G469), .ZN(n1087) );
XNOR2_X1 U848 ( .A(KEYINPUT36), .B(n1167), .ZN(n1163) );
NOR2_X1 U849 ( .A1(KEYINPUT50), .A2(n1168), .ZN(n1167) );
NOR3_X1 U850 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1168) );
NOR2_X1 U851 ( .A1(n1158), .A2(n1172), .ZN(n1171) );
NOR3_X1 U852 ( .A1(n1156), .A2(n1173), .A3(n1174), .ZN(n1170) );
INV_X1 U853 ( .A(n1172), .ZN(n1174) );
NAND2_X1 U854 ( .A1(n1106), .A2(n1175), .ZN(n1172) );
XOR2_X1 U855 ( .A(KEYINPUT57), .B(n1176), .Z(n1175) );
INV_X1 U856 ( .A(n1177), .ZN(n1169) );
NOR2_X1 U857 ( .A1(n1178), .A2(n1179), .ZN(G51) );
XNOR2_X1 U858 ( .A(n1127), .B(KEYINPUT4), .ZN(n1179) );
AND2_X1 U859 ( .A1(G953), .A2(n1180), .ZN(n1127) );
XOR2_X1 U860 ( .A(KEYINPUT51), .B(G952), .Z(n1180) );
XNOR2_X1 U861 ( .A(n1181), .B(n1182), .ZN(n1178) );
NOR2_X1 U862 ( .A1(n1183), .A2(n1132), .ZN(n1182) );
NAND2_X1 U863 ( .A1(G902), .A2(n1028), .ZN(n1132) );
INV_X1 U864 ( .A(n1139), .ZN(n1028) );
NOR4_X1 U865 ( .A1(n1097), .A2(n1116), .A3(n1184), .A4(n1185), .ZN(n1139) );
XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n1096), .ZN(n1185) );
NOR3_X1 U867 ( .A1(n1186), .A2(n1187), .A3(n1031), .ZN(n1096) );
INV_X1 U868 ( .A(n1065), .ZN(n1031) );
XOR2_X1 U869 ( .A(KEYINPUT44), .B(n1117), .Z(n1184) );
NAND3_X1 U870 ( .A1(n1188), .A2(n1054), .A3(n1066), .ZN(n1117) );
NAND4_X1 U871 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1116) );
NOR4_X1 U872 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1144), .ZN(n1192) );
NOR3_X1 U873 ( .A1(n1196), .A2(n1039), .A3(n1187), .ZN(n1144) );
INV_X1 U874 ( .A(n1054), .ZN(n1039) );
OR2_X1 U875 ( .A1(n1197), .A2(n1198), .ZN(n1191) );
NAND3_X1 U876 ( .A1(n1067), .A2(n1188), .A3(n1199), .ZN(n1189) );
XNOR2_X1 U877 ( .A(n1044), .B(KEYINPUT56), .ZN(n1199) );
NAND4_X1 U878 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1097) );
AND4_X1 U879 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
XNOR2_X1 U880 ( .A(n1202), .B(n1208), .ZN(G48) );
NOR2_X1 U881 ( .A1(KEYINPUT37), .A2(n1209), .ZN(n1208) );
NAND3_X1 U882 ( .A1(n1063), .A2(n1068), .A3(n1210), .ZN(n1202) );
XNOR2_X1 U883 ( .A(G143), .B(n1200), .ZN(G45) );
OR4_X1 U884 ( .A1(n1186), .A2(n1198), .A3(n1211), .A4(n1212), .ZN(n1200) );
XNOR2_X1 U885 ( .A(n1201), .B(n1213), .ZN(G42) );
NOR2_X1 U886 ( .A1(KEYINPUT39), .A2(n1214), .ZN(n1213) );
NAND3_X1 U887 ( .A1(n1215), .A2(n1041), .A3(n1065), .ZN(n1201) );
XOR2_X1 U888 ( .A(n1207), .B(n1216), .Z(G39) );
NOR2_X1 U889 ( .A1(G137), .A2(KEYINPUT52), .ZN(n1216) );
NAND3_X1 U890 ( .A1(n1065), .A2(n1210), .A3(n1067), .ZN(n1207) );
XNOR2_X1 U891 ( .A(G134), .B(n1206), .ZN(G36) );
NAND3_X1 U892 ( .A1(n1217), .A2(n1066), .A3(n1065), .ZN(n1206) );
INV_X1 U893 ( .A(n1186), .ZN(n1217) );
XOR2_X1 U894 ( .A(n1218), .B(n1219), .Z(G33) );
NAND2_X1 U895 ( .A1(n1065), .A2(n1220), .ZN(n1219) );
XOR2_X1 U896 ( .A(KEYINPUT53), .B(n1221), .Z(n1220) );
NOR2_X1 U897 ( .A1(n1187), .A2(n1186), .ZN(n1221) );
NAND4_X1 U898 ( .A1(n1049), .A2(n1041), .A3(n1222), .A4(n1050), .ZN(n1186) );
NOR2_X1 U899 ( .A1(n1080), .A2(n1061), .ZN(n1065) );
INV_X1 U900 ( .A(n1060), .ZN(n1080) );
XOR2_X1 U901 ( .A(n1205), .B(n1223), .Z(G30) );
NAND2_X1 U902 ( .A1(n1224), .A2(KEYINPUT11), .ZN(n1223) );
XNOR2_X1 U903 ( .A(G128), .B(KEYINPUT1), .ZN(n1224) );
NAND3_X1 U904 ( .A1(n1066), .A2(n1068), .A3(n1210), .ZN(n1205) );
AND4_X1 U905 ( .A1(n1041), .A2(n1074), .A3(n1222), .A4(n1050), .ZN(n1210) );
XOR2_X1 U906 ( .A(n1225), .B(n1190), .Z(G3) );
NAND4_X1 U907 ( .A1(n1067), .A2(n1188), .A3(n1049), .A4(n1050), .ZN(n1190) );
INV_X1 U908 ( .A(n1196), .ZN(n1188) );
XNOR2_X1 U909 ( .A(G125), .B(n1204), .ZN(G27) );
NAND3_X1 U910 ( .A1(n1215), .A2(n1068), .A3(n1045), .ZN(n1204) );
AND3_X1 U911 ( .A1(n1063), .A2(n1222), .A3(n1044), .ZN(n1215) );
NAND2_X1 U912 ( .A1(n1033), .A2(n1226), .ZN(n1222) );
NAND4_X1 U913 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1100), .ZN(n1226) );
INV_X1 U914 ( .A(G900), .ZN(n1100) );
XOR2_X1 U915 ( .A(G122), .B(n1228), .Z(G24) );
NOR2_X1 U916 ( .A1(n1197), .A2(n1229), .ZN(n1228) );
XOR2_X1 U917 ( .A(KEYINPUT16), .B(n1068), .Z(n1229) );
NAND3_X1 U918 ( .A1(n1045), .A2(n1054), .A3(n1230), .ZN(n1197) );
NOR3_X1 U919 ( .A1(n1211), .A2(n1231), .A3(n1212), .ZN(n1230) );
INV_X1 U920 ( .A(n1232), .ZN(n1231) );
NOR2_X1 U921 ( .A1(n1050), .A2(n1074), .ZN(n1054) );
XOR2_X1 U922 ( .A(G119), .B(n1195), .Z(G21) );
AND3_X1 U923 ( .A1(n1067), .A2(n1074), .A3(n1233), .ZN(n1195) );
INV_X1 U924 ( .A(n1049), .ZN(n1074) );
XOR2_X1 U925 ( .A(G116), .B(n1194), .Z(G18) );
AND3_X1 U926 ( .A1(n1049), .A2(n1066), .A3(n1233), .ZN(n1194) );
NOR2_X1 U927 ( .A1(n1211), .A2(n1075), .ZN(n1066) );
XOR2_X1 U928 ( .A(G113), .B(n1193), .Z(G15) );
AND3_X1 U929 ( .A1(n1049), .A2(n1063), .A3(n1233), .ZN(n1193) );
AND4_X1 U930 ( .A1(n1045), .A2(n1068), .A3(n1050), .A4(n1232), .ZN(n1233) );
NOR2_X1 U931 ( .A1(n1042), .A2(n1082), .ZN(n1045) );
INV_X1 U932 ( .A(n1043), .ZN(n1082) );
XNOR2_X1 U933 ( .A(n1234), .B(KEYINPUT9), .ZN(n1042) );
INV_X1 U934 ( .A(n1187), .ZN(n1063) );
NAND2_X1 U935 ( .A1(n1235), .A2(n1236), .ZN(n1187) );
XOR2_X1 U936 ( .A(KEYINPUT29), .B(n1075), .Z(n1236) );
INV_X1 U937 ( .A(n1212), .ZN(n1075) );
XNOR2_X1 U938 ( .A(G110), .B(n1237), .ZN(G12) );
NAND4_X1 U939 ( .A1(n1067), .A2(n1044), .A3(n1238), .A4(n1239), .ZN(n1237) );
NAND2_X1 U940 ( .A1(KEYINPUT54), .A2(n1196), .ZN(n1239) );
NAND2_X1 U941 ( .A1(n1068), .A2(n1240), .ZN(n1196) );
NAND2_X1 U942 ( .A1(n1241), .A2(n1242), .ZN(n1238) );
INV_X1 U943 ( .A(KEYINPUT54), .ZN(n1242) );
NAND2_X1 U944 ( .A1(n1240), .A2(n1198), .ZN(n1241) );
INV_X1 U945 ( .A(n1068), .ZN(n1198) );
NOR2_X1 U946 ( .A1(n1060), .A2(n1061), .ZN(n1068) );
AND2_X1 U947 ( .A1(G214), .A2(n1243), .ZN(n1061) );
XNOR2_X1 U948 ( .A(n1244), .B(n1183), .ZN(n1060) );
NAND2_X1 U949 ( .A1(G210), .A2(n1243), .ZN(n1183) );
NAND2_X1 U950 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
XNOR2_X1 U951 ( .A(G237), .B(KEYINPUT43), .ZN(n1245) );
NAND2_X1 U952 ( .A1(n1181), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U953 ( .A(n1247), .B(n1248), .ZN(n1181) );
XOR2_X1 U954 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U955 ( .A(G125), .B(n1251), .Z(n1250) );
NOR2_X1 U956 ( .A1(KEYINPUT38), .A2(n1252), .ZN(n1251) );
XOR2_X1 U957 ( .A(n1176), .B(n1124), .Z(n1252) );
XOR2_X1 U958 ( .A(G116), .B(n1253), .Z(n1124) );
INV_X1 U959 ( .A(n1126), .ZN(n1176) );
AND2_X1 U960 ( .A1(n1052), .A2(G224), .ZN(n1249) );
XOR2_X1 U961 ( .A(n1161), .B(n1123), .Z(n1247) );
XOR2_X1 U962 ( .A(G110), .B(n1254), .Z(n1123) );
XOR2_X1 U963 ( .A(KEYINPUT23), .B(G122), .Z(n1254) );
AND2_X1 U964 ( .A1(n1041), .A2(n1232), .ZN(n1240) );
NAND2_X1 U965 ( .A1(n1033), .A2(n1255), .ZN(n1232) );
NAND4_X1 U966 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1121), .ZN(n1255) );
INV_X1 U967 ( .A(G898), .ZN(n1121) );
NAND3_X1 U968 ( .A1(n1227), .A2(n1052), .A3(n1256), .ZN(n1033) );
XOR2_X1 U969 ( .A(KEYINPUT46), .B(G952), .Z(n1256) );
NAND2_X1 U970 ( .A1(G237), .A2(G234), .ZN(n1227) );
AND2_X1 U971 ( .A1(n1234), .A2(n1043), .ZN(n1041) );
NAND2_X1 U972 ( .A1(G221), .A2(n1257), .ZN(n1043) );
XOR2_X1 U973 ( .A(n1085), .B(n1258), .Z(n1234) );
NOR2_X1 U974 ( .A1(G469), .A2(KEYINPUT62), .ZN(n1258) );
NAND2_X1 U975 ( .A1(n1259), .A2(n1246), .ZN(n1085) );
XNOR2_X1 U976 ( .A(n1260), .B(n1166), .ZN(n1259) );
XNOR2_X1 U977 ( .A(n1261), .B(n1262), .ZN(n1166) );
XOR2_X1 U978 ( .A(G110), .B(n1263), .Z(n1262) );
AND2_X1 U979 ( .A1(n1052), .A2(G227), .ZN(n1263) );
XOR2_X1 U980 ( .A(n1214), .B(KEYINPUT14), .Z(n1261) );
INV_X1 U981 ( .A(G140), .ZN(n1214) );
NAND3_X1 U982 ( .A1(n1264), .A2(n1265), .A3(n1177), .ZN(n1260) );
NAND2_X1 U983 ( .A1(n1156), .A2(n1173), .ZN(n1177) );
NOR2_X1 U984 ( .A1(n1106), .A2(n1126), .ZN(n1173) );
NAND2_X1 U985 ( .A1(n1266), .A2(n1158), .ZN(n1265) );
XOR2_X1 U986 ( .A(n1126), .B(n1106), .Z(n1266) );
NAND3_X1 U987 ( .A1(n1106), .A2(n1126), .A3(n1156), .ZN(n1264) );
INV_X1 U988 ( .A(n1158), .ZN(n1156) );
XOR2_X1 U989 ( .A(n1225), .B(n1267), .Z(n1126) );
XOR2_X1 U990 ( .A(G107), .B(G104), .Z(n1267) );
XOR2_X1 U991 ( .A(n1268), .B(KEYINPUT49), .Z(n1106) );
NOR2_X1 U992 ( .A1(n1050), .A2(n1049), .ZN(n1044) );
XNOR2_X1 U993 ( .A(n1269), .B(n1131), .ZN(n1049) );
NAND2_X1 U994 ( .A1(G217), .A2(n1257), .ZN(n1131) );
NAND2_X1 U995 ( .A1(G234), .A2(n1246), .ZN(n1257) );
OR2_X1 U996 ( .A1(n1130), .A2(G902), .ZN(n1269) );
XNOR2_X1 U997 ( .A(n1270), .B(n1271), .ZN(n1130) );
XNOR2_X1 U998 ( .A(G137), .B(n1272), .ZN(n1271) );
NAND3_X1 U999 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1272) );
NAND2_X1 U1000 ( .A1(KEYINPUT31), .A2(n1276), .ZN(n1275) );
OR3_X1 U1001 ( .A1(n1276), .A2(KEYINPUT31), .A3(n1277), .ZN(n1274) );
NAND2_X1 U1002 ( .A1(n1277), .A2(n1278), .ZN(n1273) );
NAND2_X1 U1003 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U1004 ( .A(KEYINPUT31), .ZN(n1280) );
XNOR2_X1 U1005 ( .A(KEYINPUT59), .B(n1276), .ZN(n1279) );
XNOR2_X1 U1006 ( .A(n1281), .B(n1282), .ZN(n1276) );
NAND2_X1 U1007 ( .A1(KEYINPUT5), .A2(n1209), .ZN(n1281) );
XOR2_X1 U1008 ( .A(n1283), .B(n1284), .Z(n1277) );
XOR2_X1 U1009 ( .A(G119), .B(G110), .Z(n1284) );
XOR2_X1 U1010 ( .A(n1285), .B(G128), .Z(n1283) );
XNOR2_X1 U1011 ( .A(KEYINPUT27), .B(KEYINPUT17), .ZN(n1285) );
NAND3_X1 U1012 ( .A1(G221), .A2(n1286), .A3(KEYINPUT33), .ZN(n1270) );
NAND2_X1 U1013 ( .A1(n1287), .A2(n1288), .ZN(n1050) );
NAND2_X1 U1014 ( .A1(G472), .A2(n1079), .ZN(n1288) );
XOR2_X1 U1015 ( .A(n1289), .B(KEYINPUT28), .Z(n1287) );
OR2_X1 U1016 ( .A1(n1079), .A2(G472), .ZN(n1289) );
NAND2_X1 U1017 ( .A1(n1290), .A2(n1246), .ZN(n1079) );
INV_X1 U1018 ( .A(G902), .ZN(n1246) );
XNOR2_X1 U1019 ( .A(n1291), .B(n1152), .ZN(n1290) );
AND2_X1 U1020 ( .A1(n1292), .A2(n1293), .ZN(n1152) );
NAND2_X1 U1021 ( .A1(n1294), .A2(n1225), .ZN(n1293) );
INV_X1 U1022 ( .A(G101), .ZN(n1225) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1295), .ZN(n1294) );
NAND3_X1 U1024 ( .A1(G210), .A2(n1295), .A3(G101), .ZN(n1292) );
NAND2_X1 U1025 ( .A1(n1296), .A2(n1297), .ZN(n1291) );
NAND2_X1 U1026 ( .A1(n1149), .A2(n1298), .ZN(n1297) );
XOR2_X1 U1027 ( .A(KEYINPUT42), .B(n1299), .Z(n1296) );
NOR2_X1 U1028 ( .A1(n1149), .A2(n1298), .ZN(n1299) );
XOR2_X1 U1029 ( .A(n1158), .B(n1161), .Z(n1298) );
XOR2_X1 U1030 ( .A(n1268), .B(KEYINPUT26), .Z(n1161) );
XOR2_X1 U1031 ( .A(n1209), .B(n1300), .Z(n1268) );
NAND3_X1 U1032 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1158) );
OR2_X1 U1033 ( .A1(n1108), .A2(KEYINPUT13), .ZN(n1303) );
NAND3_X1 U1034 ( .A1(KEYINPUT13), .A2(n1304), .A3(n1218), .ZN(n1302) );
INV_X1 U1035 ( .A(G131), .ZN(n1218) );
INV_X1 U1036 ( .A(n1305), .ZN(n1304) );
NAND2_X1 U1037 ( .A1(G131), .A2(n1305), .ZN(n1301) );
NAND2_X1 U1038 ( .A1(KEYINPUT55), .A2(n1108), .ZN(n1305) );
XOR2_X1 U1039 ( .A(G134), .B(G137), .Z(n1108) );
XNOR2_X1 U1040 ( .A(n1253), .B(n1306), .ZN(n1149) );
NOR2_X1 U1041 ( .A1(G116), .A2(KEYINPUT22), .ZN(n1306) );
XOR2_X1 U1042 ( .A(G113), .B(G119), .Z(n1253) );
INV_X1 U1043 ( .A(n1032), .ZN(n1067) );
NAND2_X1 U1044 ( .A1(n1235), .A2(n1212), .ZN(n1032) );
XOR2_X1 U1045 ( .A(n1307), .B(G475), .Z(n1212) );
OR2_X1 U1046 ( .A1(n1142), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1047 ( .A(n1308), .B(n1309), .ZN(n1142) );
XOR2_X1 U1048 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1049 ( .A(G122), .B(G104), .Z(n1311) );
XOR2_X1 U1050 ( .A(G143), .B(G131), .Z(n1310) );
XOR2_X1 U1051 ( .A(n1312), .B(n1313), .Z(n1308) );
XOR2_X1 U1052 ( .A(n1314), .B(n1315), .Z(n1313) );
AND2_X1 U1053 ( .A1(n1295), .A2(G214), .ZN(n1315) );
NOR2_X1 U1054 ( .A1(G953), .A2(G237), .ZN(n1295) );
NOR2_X1 U1055 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
XOR2_X1 U1056 ( .A(KEYINPUT32), .B(n1318), .Z(n1317) );
NOR2_X1 U1057 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
AND2_X1 U1058 ( .A1(n1320), .A2(n1319), .ZN(n1316) );
XNOR2_X1 U1059 ( .A(n1282), .B(KEYINPUT63), .ZN(n1319) );
INV_X1 U1060 ( .A(n1104), .ZN(n1282) );
XOR2_X1 U1061 ( .A(G125), .B(G140), .Z(n1104) );
XNOR2_X1 U1062 ( .A(n1209), .B(KEYINPUT45), .ZN(n1320) );
INV_X1 U1063 ( .A(G146), .ZN(n1209) );
NAND2_X1 U1064 ( .A1(KEYINPUT58), .A2(n1321), .ZN(n1312) );
INV_X1 U1065 ( .A(G113), .ZN(n1321) );
XNOR2_X1 U1066 ( .A(n1211), .B(KEYINPUT0), .ZN(n1235) );
XOR2_X1 U1067 ( .A(n1084), .B(n1322), .Z(n1211) );
XOR2_X1 U1068 ( .A(KEYINPUT6), .B(G478), .Z(n1322) );
NOR2_X1 U1069 ( .A1(G902), .A2(n1137), .ZN(n1084) );
INV_X1 U1070 ( .A(n1136), .ZN(n1137) );
NAND2_X1 U1071 ( .A1(n1323), .A2(n1324), .ZN(n1136) );
NAND2_X1 U1072 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1073 ( .A(n1327), .B(n1328), .Z(n1323) );
NOR2_X1 U1074 ( .A1(n1325), .A2(n1326), .ZN(n1328) );
INV_X1 U1075 ( .A(KEYINPUT25), .ZN(n1326) );
XOR2_X1 U1076 ( .A(n1329), .B(n1330), .Z(n1325) );
XOR2_X1 U1077 ( .A(n1331), .B(n1300), .Z(n1330) );
XOR2_X1 U1078 ( .A(G128), .B(G143), .Z(n1300) );
NOR4_X1 U1079 ( .A1(n1332), .A2(n1333), .A3(KEYINPUT7), .A4(n1334), .ZN(n1331) );
AND2_X1 U1080 ( .A1(n1335), .A2(G116), .ZN(n1334) );
NOR2_X1 U1081 ( .A1(n1336), .A2(n1337), .ZN(n1333) );
INV_X1 U1082 ( .A(G122), .ZN(n1337) );
NOR2_X1 U1083 ( .A1(G116), .A2(KEYINPUT12), .ZN(n1336) );
NOR4_X1 U1084 ( .A1(G122), .A2(n1335), .A3(KEYINPUT12), .A4(G116), .ZN(n1332) );
INV_X1 U1085 ( .A(KEYINPUT47), .ZN(n1335) );
XNOR2_X1 U1086 ( .A(G107), .B(G134), .ZN(n1329) );
NAND2_X1 U1087 ( .A1(G217), .A2(n1286), .ZN(n1327) );
AND2_X1 U1088 ( .A1(G234), .A2(n1052), .ZN(n1286) );
INV_X1 U1089 ( .A(G953), .ZN(n1052) );
endmodule


