//Key = 1011110000111001010101001110011110101101000100100000100101000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368;

XNOR2_X1 U750 ( .A(G107), .B(n1048), .ZN(G9) );
NAND3_X1 U751 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
XNOR2_X1 U752 ( .A(n1052), .B(KEYINPUT36), .ZN(n1051) );
NAND4_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(G75) );
NAND3_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR3_X1 U755 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
XNOR2_X1 U756 ( .A(n1063), .B(n1064), .ZN(n1062) );
XNOR2_X1 U757 ( .A(KEYINPUT2), .B(n1065), .ZN(n1064) );
NOR2_X1 U758 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
NOR2_X1 U759 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U760 ( .A1(KEYINPUT28), .A2(n1070), .ZN(n1068) );
NOR2_X1 U761 ( .A1(KEYINPUT35), .A2(n1071), .ZN(n1070) );
NOR2_X1 U762 ( .A1(G472), .A2(n1072), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1073), .A2(KEYINPUT35), .ZN(n1072) );
NOR2_X1 U764 ( .A1(KEYINPUT28), .A2(n1074), .ZN(n1073) );
XOR2_X1 U765 ( .A(n1075), .B(n1076), .Z(n1060) );
NOR2_X1 U766 ( .A1(n1077), .A2(KEYINPUT27), .ZN(n1076) );
INV_X1 U767 ( .A(n1078), .ZN(n1077) );
XNOR2_X1 U768 ( .A(n1079), .B(n1080), .ZN(n1058) );
NOR2_X1 U769 ( .A1(KEYINPUT22), .A2(n1081), .ZN(n1080) );
XNOR2_X1 U770 ( .A(KEYINPUT42), .B(n1082), .ZN(n1081) );
XNOR2_X1 U771 ( .A(n1083), .B(KEYINPUT21), .ZN(n1057) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1054) );
NAND2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U774 ( .A1(n1052), .A2(n1088), .A3(n1089), .ZN(n1087) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NAND3_X1 U776 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND3_X1 U778 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1092) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
NAND2_X1 U780 ( .A1(n1102), .A2(n1103), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1104), .ZN(n1086) );
NAND3_X1 U782 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
INV_X1 U783 ( .A(n1108), .ZN(n1107) );
NAND2_X1 U784 ( .A1(n1109), .A2(n1052), .ZN(n1106) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1110), .ZN(n1105) );
NOR3_X1 U786 ( .A1(n1096), .A2(n1095), .A3(n1111), .ZN(n1083) );
INV_X1 U787 ( .A(n1112), .ZN(n1084) );
XOR2_X1 U788 ( .A(n1113), .B(n1114), .Z(G72) );
XOR2_X1 U789 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U790 ( .A1(n1117), .A2(KEYINPUT13), .ZN(n1116) );
NOR2_X1 U791 ( .A1(n1118), .A2(G953), .ZN(n1117) );
NOR2_X1 U792 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U793 ( .A(n1121), .B(KEYINPUT34), .ZN(n1119) );
NAND2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
NAND2_X1 U795 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U796 ( .A(n1125), .B(n1126), .Z(n1122) );
XOR2_X1 U797 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U798 ( .A(KEYINPUT16), .B(n1129), .ZN(n1125) );
NOR3_X1 U799 ( .A1(n1130), .A2(KEYINPUT50), .A3(n1131), .ZN(n1129) );
XOR2_X1 U800 ( .A(KEYINPUT60), .B(n1132), .Z(n1130) );
NOR2_X1 U801 ( .A1(G140), .A2(n1133), .ZN(n1132) );
NAND2_X1 U802 ( .A1(KEYINPUT3), .A2(n1134), .ZN(n1113) );
NAND2_X1 U803 ( .A1(G953), .A2(n1135), .ZN(n1134) );
NAND2_X1 U804 ( .A1(n1136), .A2(G900), .ZN(n1135) );
XNOR2_X1 U805 ( .A(G227), .B(KEYINPUT25), .ZN(n1136) );
NAND2_X1 U806 ( .A1(n1137), .A2(n1138), .ZN(G69) );
NAND2_X1 U807 ( .A1(n1139), .A2(G953), .ZN(n1138) );
XOR2_X1 U808 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U809 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U810 ( .A1(n1144), .A2(n1056), .ZN(n1137) );
NAND2_X1 U811 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U812 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
OR2_X1 U813 ( .A1(n1140), .A2(n1148), .ZN(n1145) );
XOR2_X1 U814 ( .A(n1147), .B(KEYINPUT44), .Z(n1140) );
NAND3_X1 U815 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1147) );
NAND2_X1 U816 ( .A1(G953), .A2(n1143), .ZN(n1151) );
NAND2_X1 U817 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
XOR2_X1 U818 ( .A(n1154), .B(KEYINPUT8), .Z(n1152) );
NOR2_X1 U819 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XNOR2_X1 U820 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U821 ( .A1(n1078), .A2(n1159), .ZN(n1157) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1160), .ZN(G63) );
NOR3_X1 U823 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
NOR3_X1 U824 ( .A1(n1164), .A2(n1079), .A3(n1159), .ZN(n1163) );
NOR2_X1 U825 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
NOR2_X1 U826 ( .A1(n1053), .A2(n1079), .ZN(n1165) );
INV_X1 U827 ( .A(G478), .ZN(n1079) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1167), .ZN(G60) );
NOR3_X1 U829 ( .A1(n1063), .A2(n1168), .A3(n1169), .ZN(n1167) );
NOR3_X1 U830 ( .A1(n1170), .A2(n1065), .A3(n1159), .ZN(n1169) );
INV_X1 U831 ( .A(n1171), .ZN(n1170) );
NOR2_X1 U832 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1053), .A2(n1065), .ZN(n1172) );
XNOR2_X1 U834 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1174), .ZN(G57) );
XOR2_X1 U836 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U837 ( .A(n1177), .B(n1178), .ZN(n1176) );
XNOR2_X1 U838 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U839 ( .A1(KEYINPUT47), .A2(n1181), .ZN(n1180) );
INV_X1 U840 ( .A(n1182), .ZN(n1181) );
NAND2_X1 U841 ( .A1(KEYINPUT17), .A2(n1183), .ZN(n1179) );
XOR2_X1 U842 ( .A(n1184), .B(n1185), .Z(n1175) );
NOR2_X1 U843 ( .A1(n1071), .A2(n1159), .ZN(n1185) );
XOR2_X1 U844 ( .A(n1186), .B(KEYINPUT48), .Z(n1184) );
NOR2_X1 U845 ( .A1(n1155), .A2(n1187), .ZN(G54) );
XOR2_X1 U846 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U847 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U848 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U849 ( .A(n1194), .B(KEYINPUT39), .Z(n1193) );
NAND2_X1 U850 ( .A1(n1195), .A2(n1182), .ZN(n1194) );
NOR2_X1 U851 ( .A1(n1195), .A2(n1182), .ZN(n1192) );
XOR2_X1 U852 ( .A(n1196), .B(n1128), .Z(n1195) );
NAND2_X1 U853 ( .A1(KEYINPUT10), .A2(n1197), .ZN(n1196) );
NOR2_X1 U854 ( .A1(n1198), .A2(n1159), .ZN(n1188) );
NOR2_X1 U855 ( .A1(n1155), .A2(n1199), .ZN(G51) );
XOR2_X1 U856 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U857 ( .A(n1202), .B(n1203), .Z(n1200) );
NOR2_X1 U858 ( .A1(n1204), .A2(n1159), .ZN(n1203) );
OR2_X1 U859 ( .A1(n1205), .A2(n1053), .ZN(n1159) );
NOR3_X1 U860 ( .A1(n1148), .A2(n1121), .A3(n1120), .ZN(n1053) );
NAND4_X1 U861 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1120) );
AND4_X1 U862 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND3_X1 U863 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1208) );
XNOR2_X1 U864 ( .A(KEYINPUT14), .B(n1098), .ZN(n1214) );
INV_X1 U865 ( .A(n1217), .ZN(n1098) );
INV_X1 U866 ( .A(n1218), .ZN(n1121) );
NAND4_X1 U867 ( .A1(n1219), .A2(n1173), .A3(n1220), .A4(n1221), .ZN(n1148) );
AND4_X1 U868 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
OR2_X1 U869 ( .A1(n1226), .A2(n1227), .ZN(n1220) );
NAND3_X1 U870 ( .A1(n1050), .A2(n1052), .A3(n1109), .ZN(n1173) );
NAND2_X1 U871 ( .A1(n1050), .A2(n1108), .ZN(n1219) );
NAND2_X1 U872 ( .A1(n1228), .A2(n1229), .ZN(n1108) );
NAND2_X1 U873 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U874 ( .A1(n1049), .A2(n1052), .ZN(n1228) );
NAND2_X1 U875 ( .A1(KEYINPUT29), .A2(n1232), .ZN(n1202) );
XNOR2_X1 U876 ( .A(KEYINPUT18), .B(n1186), .ZN(n1232) );
NOR2_X1 U877 ( .A1(n1056), .A2(G952), .ZN(n1155) );
XNOR2_X1 U878 ( .A(G146), .B(n1206), .ZN(G48) );
NAND2_X1 U879 ( .A1(n1233), .A2(n1109), .ZN(n1206) );
XOR2_X1 U880 ( .A(n1234), .B(n1235), .Z(G45) );
XNOR2_X1 U881 ( .A(G143), .B(KEYINPUT40), .ZN(n1235) );
NAND3_X1 U882 ( .A1(n1216), .A2(n1236), .A3(KEYINPUT19), .ZN(n1234) );
AND4_X1 U883 ( .A1(n1237), .A2(n1110), .A3(n1103), .A4(n1238), .ZN(n1216) );
XNOR2_X1 U884 ( .A(G140), .B(n1207), .ZN(G42) );
NAND2_X1 U885 ( .A1(n1239), .A2(n1240), .ZN(n1207) );
XNOR2_X1 U886 ( .A(G137), .B(n1213), .ZN(G39) );
NAND3_X1 U887 ( .A1(n1239), .A2(n1241), .A3(n1230), .ZN(n1213) );
XNOR2_X1 U888 ( .A(G134), .B(n1212), .ZN(G36) );
NAND3_X1 U889 ( .A1(n1239), .A2(n1049), .A3(n1110), .ZN(n1212) );
XNOR2_X1 U890 ( .A(G131), .B(n1218), .ZN(G33) );
NAND3_X1 U891 ( .A1(n1239), .A2(n1109), .A3(n1110), .ZN(n1218) );
AND3_X1 U892 ( .A1(n1236), .A2(n1099), .A3(n1094), .ZN(n1239) );
XOR2_X1 U893 ( .A(n1211), .B(n1242), .Z(G30) );
NAND2_X1 U894 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1242) );
NAND2_X1 U895 ( .A1(n1233), .A2(n1049), .ZN(n1211) );
AND4_X1 U896 ( .A1(n1243), .A2(n1236), .A3(n1103), .A4(n1241), .ZN(n1233) );
AND2_X1 U897 ( .A1(n1217), .A2(n1215), .ZN(n1236) );
XNOR2_X1 U898 ( .A(G101), .B(n1225), .ZN(G3) );
NAND3_X1 U899 ( .A1(n1110), .A2(n1050), .A3(n1089), .ZN(n1225) );
AND3_X1 U900 ( .A1(n1217), .A2(n1244), .A3(n1103), .ZN(n1050) );
XOR2_X1 U901 ( .A(n1210), .B(n1245), .Z(G27) );
XNOR2_X1 U902 ( .A(G125), .B(KEYINPUT20), .ZN(n1245) );
NAND4_X1 U903 ( .A1(n1102), .A2(n1240), .A3(n1103), .A4(n1215), .ZN(n1210) );
NAND2_X1 U904 ( .A1(n1246), .A2(n1112), .ZN(n1215) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1124), .A4(n1247), .ZN(n1246) );
XOR2_X1 U906 ( .A(KEYINPUT57), .B(G900), .Z(n1124) );
AND3_X1 U907 ( .A1(n1231), .A2(n1243), .A3(n1109), .ZN(n1240) );
XNOR2_X1 U908 ( .A(G122), .B(n1224), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1237), .A2(n1248), .A3(n1052), .A4(n1238), .ZN(n1224) );
NOR2_X1 U910 ( .A1(n1241), .A2(n1243), .ZN(n1052) );
XNOR2_X1 U911 ( .A(G119), .B(n1223), .ZN(G21) );
NAND3_X1 U912 ( .A1(n1230), .A2(n1241), .A3(n1248), .ZN(n1223) );
INV_X1 U913 ( .A(n1249), .ZN(n1230) );
XNOR2_X1 U914 ( .A(G116), .B(n1222), .ZN(G18) );
NAND3_X1 U915 ( .A1(n1110), .A2(n1049), .A3(n1248), .ZN(n1222) );
AND3_X1 U916 ( .A1(n1103), .A2(n1244), .A3(n1102), .ZN(n1248) );
NOR2_X1 U917 ( .A1(n1237), .A2(n1250), .ZN(n1049) );
XNOR2_X1 U918 ( .A(n1251), .B(n1252), .ZN(G15) );
NOR2_X1 U919 ( .A1(n1253), .A2(n1227), .ZN(n1252) );
XOR2_X1 U920 ( .A(n1226), .B(KEYINPUT7), .Z(n1253) );
NAND4_X1 U921 ( .A1(n1110), .A2(n1102), .A3(n1109), .A4(n1244), .ZN(n1226) );
AND2_X1 U922 ( .A1(n1250), .A2(n1237), .ZN(n1109) );
INV_X1 U923 ( .A(n1238), .ZN(n1250) );
INV_X1 U924 ( .A(n1096), .ZN(n1102) );
NAND2_X1 U925 ( .A1(n1101), .A2(n1254), .ZN(n1096) );
NOR2_X1 U926 ( .A1(n1231), .A2(n1243), .ZN(n1110) );
INV_X1 U927 ( .A(n1241), .ZN(n1231) );
XNOR2_X1 U928 ( .A(G110), .B(n1255), .ZN(G12) );
NAND4_X1 U929 ( .A1(n1256), .A2(n1244), .A3(n1217), .A4(n1257), .ZN(n1255) );
NOR2_X1 U930 ( .A1(n1249), .A2(n1241), .ZN(n1257) );
XNOR2_X1 U931 ( .A(n1074), .B(n1071), .ZN(n1241) );
INV_X1 U932 ( .A(G472), .ZN(n1071) );
INV_X1 U933 ( .A(n1069), .ZN(n1074) );
NAND2_X1 U934 ( .A1(n1258), .A2(n1205), .ZN(n1069) );
XOR2_X1 U935 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U936 ( .A(n1186), .B(n1261), .Z(n1260) );
XNOR2_X1 U937 ( .A(KEYINPUT56), .B(KEYINPUT4), .ZN(n1261) );
XNOR2_X1 U938 ( .A(n1262), .B(n1183), .ZN(n1259) );
XOR2_X1 U939 ( .A(n1263), .B(n1264), .Z(n1183) );
XNOR2_X1 U940 ( .A(n1265), .B(G116), .ZN(n1264) );
NAND2_X1 U941 ( .A1(KEYINPUT37), .A2(n1251), .ZN(n1263) );
INV_X1 U942 ( .A(G113), .ZN(n1251) );
XNOR2_X1 U943 ( .A(n1182), .B(n1177), .ZN(n1262) );
XNOR2_X1 U944 ( .A(n1266), .B(G101), .ZN(n1177) );
NAND2_X1 U945 ( .A1(G210), .A2(n1267), .ZN(n1266) );
NAND2_X1 U946 ( .A1(n1089), .A2(n1243), .ZN(n1249) );
XOR2_X1 U947 ( .A(n1078), .B(n1268), .Z(n1243) );
NOR2_X1 U948 ( .A1(KEYINPUT38), .A2(n1269), .ZN(n1268) );
XOR2_X1 U949 ( .A(n1075), .B(KEYINPUT31), .Z(n1269) );
NAND2_X1 U950 ( .A1(n1270), .A2(n1158), .ZN(n1075) );
XNOR2_X1 U951 ( .A(n1271), .B(n1272), .ZN(n1158) );
XOR2_X1 U952 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR3_X1 U953 ( .A1(n1275), .A2(KEYINPUT1), .A3(n1276), .ZN(n1274) );
NOR4_X1 U954 ( .A1(G953), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1276) );
NOR2_X1 U955 ( .A1(n1280), .A2(n1281), .ZN(n1275) );
XNOR2_X1 U956 ( .A(G137), .B(KEYINPUT5), .ZN(n1281) );
NOR3_X1 U957 ( .A1(n1278), .A2(G953), .A3(n1277), .ZN(n1280) );
INV_X1 U958 ( .A(G221), .ZN(n1278) );
NAND2_X1 U959 ( .A1(n1282), .A2(n1283), .ZN(n1273) );
NAND2_X1 U960 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U961 ( .A(n1265), .B(n1286), .ZN(n1285) );
XNOR2_X1 U962 ( .A(KEYINPUT6), .B(G110), .ZN(n1284) );
XOR2_X1 U963 ( .A(n1287), .B(KEYINPUT33), .Z(n1282) );
NAND2_X1 U964 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U965 ( .A(KEYINPUT6), .B(G110), .Z(n1289) );
XNOR2_X1 U966 ( .A(G119), .B(n1286), .ZN(n1288) );
NOR2_X1 U967 ( .A1(G128), .A2(KEYINPUT9), .ZN(n1286) );
XNOR2_X1 U968 ( .A(G902), .B(KEYINPUT63), .ZN(n1270) );
NAND2_X1 U969 ( .A1(G217), .A2(n1290), .ZN(n1078) );
NOR2_X1 U970 ( .A1(n1238), .A2(n1237), .ZN(n1089) );
XNOR2_X1 U971 ( .A(n1291), .B(n1065), .ZN(n1237) );
INV_X1 U972 ( .A(G475), .ZN(n1065) );
NAND2_X1 U973 ( .A1(KEYINPUT32), .A2(n1292), .ZN(n1291) );
INV_X1 U974 ( .A(n1063), .ZN(n1292) );
NOR2_X1 U975 ( .A1(n1171), .A2(G902), .ZN(n1063) );
XNOR2_X1 U976 ( .A(n1293), .B(n1294), .ZN(n1171) );
NOR2_X1 U977 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U978 ( .A(n1297), .B(KEYINPUT24), .Z(n1296) );
NAND2_X1 U979 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR2_X1 U980 ( .A1(n1298), .A2(n1299), .ZN(n1295) );
XNOR2_X1 U981 ( .A(G113), .B(G122), .ZN(n1298) );
NAND2_X1 U982 ( .A1(KEYINPUT11), .A2(n1300), .ZN(n1293) );
XOR2_X1 U983 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U984 ( .A(n1303), .B(n1272), .Z(n1302) );
NAND2_X1 U985 ( .A1(n1304), .A2(n1305), .ZN(n1272) );
NAND2_X1 U986 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U987 ( .A1(n1308), .A2(n1309), .ZN(n1306) );
NAND2_X1 U988 ( .A1(G125), .A2(n1310), .ZN(n1309) );
INV_X1 U989 ( .A(n1131), .ZN(n1308) );
NOR2_X1 U990 ( .A1(n1310), .A2(G125), .ZN(n1131) );
NAND2_X1 U991 ( .A1(G146), .A2(n1311), .ZN(n1304) );
XNOR2_X1 U992 ( .A(G125), .B(G140), .ZN(n1311) );
NAND2_X1 U993 ( .A1(KEYINPUT46), .A2(n1312), .ZN(n1303) );
INV_X1 U994 ( .A(G131), .ZN(n1312) );
XOR2_X1 U995 ( .A(n1313), .B(G143), .Z(n1301) );
NAND2_X1 U996 ( .A1(G214), .A2(n1267), .ZN(n1313) );
NOR2_X1 U997 ( .A1(G953), .A2(G237), .ZN(n1267) );
XOR2_X1 U998 ( .A(G478), .B(n1314), .Z(n1238) );
NOR2_X1 U999 ( .A1(KEYINPUT62), .A2(n1082), .ZN(n1314) );
INV_X1 U1000 ( .A(n1161), .ZN(n1082) );
NOR2_X1 U1001 ( .A1(n1166), .A2(G902), .ZN(n1161) );
INV_X1 U1002 ( .A(n1164), .ZN(n1166) );
XNOR2_X1 U1003 ( .A(n1315), .B(n1316), .ZN(n1164) );
NOR2_X1 U1004 ( .A1(KEYINPUT23), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1005 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1006 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U1007 ( .A1(KEYINPUT61), .A2(G134), .ZN(n1320) );
XOR2_X1 U1008 ( .A(n1322), .B(KEYINPUT26), .Z(n1318) );
NAND2_X1 U1009 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND3_X1 U1010 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1324) );
XNOR2_X1 U1011 ( .A(n1328), .B(n1329), .ZN(n1327) );
INV_X1 U1012 ( .A(G107), .ZN(n1329) );
NAND2_X1 U1013 ( .A1(KEYINPUT43), .A2(G122), .ZN(n1328) );
NAND2_X1 U1014 ( .A1(n1330), .A2(n1331), .ZN(n1323) );
NAND2_X1 U1015 ( .A1(n1325), .A2(n1326), .ZN(n1331) );
INV_X1 U1016 ( .A(KEYINPUT58), .ZN(n1326) );
INV_X1 U1017 ( .A(G116), .ZN(n1325) );
XNOR2_X1 U1018 ( .A(G107), .B(n1332), .ZN(n1330) );
AND2_X1 U1019 ( .A1(n1333), .A2(KEYINPUT43), .ZN(n1332) );
NAND3_X1 U1020 ( .A1(n1334), .A2(n1056), .A3(G217), .ZN(n1315) );
INV_X1 U1021 ( .A(n1277), .ZN(n1334) );
XOR2_X1 U1022 ( .A(G234), .B(KEYINPUT15), .Z(n1277) );
NOR2_X1 U1023 ( .A1(n1101), .A2(n1100), .ZN(n1217) );
INV_X1 U1024 ( .A(n1254), .ZN(n1100) );
NAND2_X1 U1025 ( .A1(G221), .A2(n1290), .ZN(n1254) );
NAND2_X1 U1026 ( .A1(G234), .A2(n1205), .ZN(n1290) );
XNOR2_X1 U1027 ( .A(n1335), .B(n1198), .ZN(n1101) );
INV_X1 U1028 ( .A(G469), .ZN(n1198) );
NAND2_X1 U1029 ( .A1(n1336), .A2(n1205), .ZN(n1335) );
XOR2_X1 U1030 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1031 ( .A(n1197), .B(n1128), .ZN(n1338) );
XNOR2_X1 U1032 ( .A(n1339), .B(n1321), .ZN(n1128) );
XOR2_X1 U1033 ( .A(G128), .B(G143), .Z(n1321) );
XNOR2_X1 U1034 ( .A(G146), .B(KEYINPUT54), .ZN(n1339) );
XNOR2_X1 U1035 ( .A(n1340), .B(G101), .ZN(n1197) );
XNOR2_X1 U1036 ( .A(n1182), .B(n1190), .ZN(n1337) );
AND2_X1 U1037 ( .A1(n1341), .A2(n1342), .ZN(n1190) );
NAND3_X1 U1038 ( .A1(G227), .A2(n1056), .A3(n1343), .ZN(n1342) );
XNOR2_X1 U1039 ( .A(G110), .B(G140), .ZN(n1343) );
NAND2_X1 U1040 ( .A1(n1344), .A2(n1345), .ZN(n1341) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1056), .ZN(n1345) );
XNOR2_X1 U1042 ( .A(n1310), .B(G110), .ZN(n1344) );
INV_X1 U1043 ( .A(G140), .ZN(n1310) );
XNOR2_X1 U1044 ( .A(n1127), .B(KEYINPUT41), .ZN(n1182) );
XNOR2_X1 U1045 ( .A(G131), .B(n1346), .ZN(n1127) );
XNOR2_X1 U1046 ( .A(n1279), .B(G134), .ZN(n1346) );
INV_X1 U1047 ( .A(G137), .ZN(n1279) );
NAND2_X1 U1048 ( .A1(n1112), .A2(n1347), .ZN(n1244) );
NAND4_X1 U1049 ( .A1(G953), .A2(G902), .A3(n1247), .A4(n1143), .ZN(n1347) );
INV_X1 U1050 ( .A(G898), .ZN(n1143) );
NAND3_X1 U1051 ( .A1(n1247), .A2(n1056), .A3(G952), .ZN(n1112) );
INV_X1 U1052 ( .A(G953), .ZN(n1056) );
NAND2_X1 U1053 ( .A1(G237), .A2(G234), .ZN(n1247) );
XNOR2_X1 U1054 ( .A(KEYINPUT45), .B(n1227), .ZN(n1256) );
INV_X1 U1055 ( .A(n1103), .ZN(n1227) );
NOR2_X1 U1056 ( .A1(n1094), .A2(n1095), .ZN(n1103) );
INV_X1 U1057 ( .A(n1099), .ZN(n1095) );
NAND2_X1 U1058 ( .A1(G214), .A2(n1348), .ZN(n1099) );
INV_X1 U1059 ( .A(n1111), .ZN(n1094) );
XOR2_X1 U1060 ( .A(n1349), .B(n1204), .Z(n1111) );
NAND2_X1 U1061 ( .A1(G210), .A2(n1348), .ZN(n1204) );
NAND2_X1 U1062 ( .A1(n1205), .A2(n1350), .ZN(n1348) );
INV_X1 U1063 ( .A(G237), .ZN(n1350) );
NAND2_X1 U1064 ( .A1(n1351), .A2(n1205), .ZN(n1349) );
INV_X1 U1065 ( .A(G902), .ZN(n1205) );
XNOR2_X1 U1066 ( .A(n1201), .B(n1352), .ZN(n1351) );
XOR2_X1 U1067 ( .A(n1186), .B(KEYINPUT59), .Z(n1352) );
NAND3_X1 U1068 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1186) );
OR2_X1 U1069 ( .A1(n1356), .A2(KEYINPUT0), .ZN(n1355) );
NAND3_X1 U1070 ( .A1(KEYINPUT0), .A2(n1357), .A3(G128), .ZN(n1354) );
OR2_X1 U1071 ( .A1(n1357), .A2(G128), .ZN(n1353) );
AND2_X1 U1072 ( .A1(KEYINPUT30), .A2(n1356), .ZN(n1357) );
XNOR2_X1 U1073 ( .A(n1358), .B(G143), .ZN(n1356) );
NAND2_X1 U1074 ( .A1(KEYINPUT12), .A2(n1307), .ZN(n1358) );
INV_X1 U1075 ( .A(G146), .ZN(n1307) );
XNOR2_X1 U1076 ( .A(n1359), .B(n1360), .ZN(n1201) );
NOR2_X1 U1077 ( .A1(G953), .A2(n1142), .ZN(n1360) );
INV_X1 U1078 ( .A(G224), .ZN(n1142) );
XNOR2_X1 U1079 ( .A(n1361), .B(n1133), .ZN(n1359) );
INV_X1 U1080 ( .A(G125), .ZN(n1133) );
NAND2_X1 U1081 ( .A1(n1150), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1082 ( .A1(n1363), .A2(n1153), .ZN(n1362) );
XOR2_X1 U1083 ( .A(n1154), .B(KEYINPUT53), .Z(n1363) );
OR2_X1 U1084 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
XOR2_X1 U1085 ( .A(n1364), .B(n1365), .Z(n1154) );
XNOR2_X1 U1086 ( .A(n1333), .B(G110), .ZN(n1365) );
INV_X1 U1087 ( .A(G122), .ZN(n1333) );
XOR2_X1 U1088 ( .A(n1340), .B(n1366), .Z(n1364) );
NOR2_X1 U1089 ( .A1(G101), .A2(KEYINPUT49), .ZN(n1366) );
XNOR2_X1 U1090 ( .A(G107), .B(n1299), .ZN(n1340) );
XOR2_X1 U1091 ( .A(G104), .B(KEYINPUT55), .Z(n1299) );
XNOR2_X1 U1092 ( .A(n1367), .B(n1368), .ZN(n1153) );
NOR2_X1 U1093 ( .A1(KEYINPUT51), .A2(n1265), .ZN(n1368) );
INV_X1 U1094 ( .A(G119), .ZN(n1265) );
XNOR2_X1 U1095 ( .A(G113), .B(G116), .ZN(n1367) );
endmodule


