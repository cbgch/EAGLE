//Key = 1010110011100100011000110000000111011101100110011110010001010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366;

XOR2_X1 U751 ( .A(G107), .B(n1046), .Z(G9) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U753 ( .A1(G953), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1048) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR4_X1 U756 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
NOR2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
NOR2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR3_X1 U759 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1062) );
NOR2_X1 U761 ( .A1(n1069), .A2(n1070), .ZN(n1056) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1071), .ZN(n1069) );
NOR4_X1 U763 ( .A1(n1064), .A2(n1072), .A3(n1071), .A4(n1060), .ZN(n1054) );
NOR2_X1 U764 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U765 ( .A1(n1075), .A2(n1058), .ZN(n1074) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U768 ( .A1(n1080), .A2(n1059), .ZN(n1073) );
NOR2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
INV_X1 U771 ( .A(n1085), .ZN(n1052) );
NOR3_X1 U772 ( .A1(n1049), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U773 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1049) );
NOR4_X1 U774 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
XNOR2_X1 U775 ( .A(n1094), .B(n1095), .ZN(n1091) );
NAND2_X1 U776 ( .A1(KEYINPUT5), .A2(n1096), .ZN(n1094) );
INV_X1 U777 ( .A(G472), .ZN(n1096) );
XOR2_X1 U778 ( .A(n1070), .B(KEYINPUT13), .Z(n1090) );
XOR2_X1 U779 ( .A(n1097), .B(G475), .Z(n1088) );
XOR2_X1 U780 ( .A(n1068), .B(KEYINPUT45), .Z(n1086) );
XOR2_X1 U781 ( .A(n1098), .B(n1099), .Z(G72) );
XOR2_X1 U782 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U783 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U785 ( .A(KEYINPUT40), .B(KEYINPUT11), .Z(n1105) );
XNOR2_X1 U786 ( .A(n1106), .B(n1107), .ZN(n1104) );
NAND2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U789 ( .A(KEYINPUT53), .B(n1112), .Z(n1108) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1112) );
XOR2_X1 U791 ( .A(G137), .B(n1113), .Z(n1111) );
NOR2_X1 U792 ( .A1(G900), .A2(n1114), .ZN(n1102) );
NOR2_X1 U793 ( .A1(KEYINPUT20), .A2(n1115), .ZN(n1100) );
NOR2_X1 U794 ( .A1(n1116), .A2(G953), .ZN(n1115) );
NOR2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U796 ( .A(KEYINPUT59), .B(n1119), .ZN(n1118) );
NAND3_X1 U797 ( .A1(G953), .A2(n1120), .A3(KEYINPUT10), .ZN(n1098) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1121), .B(n1122), .Z(G69) );
NOR2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U801 ( .A(KEYINPUT42), .B(n1125), .Z(n1124) );
NOR3_X1 U802 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
AND3_X1 U803 ( .A1(n1126), .A2(n1114), .A3(n1128), .ZN(n1123) );
XNOR2_X1 U804 ( .A(n1129), .B(n1130), .ZN(n1126) );
NAND2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
INV_X1 U806 ( .A(n1133), .ZN(n1132) );
NAND2_X1 U807 ( .A1(G953), .A2(n1134), .ZN(n1121) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1134) );
NOR2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR3_X1 U811 ( .A1(n1139), .A2(KEYINPUT21), .A3(n1140), .ZN(n1138) );
XOR2_X1 U812 ( .A(KEYINPUT31), .B(G217), .Z(n1139) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1141), .ZN(G63) );
XOR2_X1 U814 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U815 ( .A1(n1144), .A2(G478), .ZN(n1142) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1145), .ZN(G60) );
NOR3_X1 U817 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1145) );
NOR2_X1 U818 ( .A1(KEYINPUT49), .A2(n1149), .ZN(n1148) );
NOR2_X1 U819 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NOR3_X1 U823 ( .A1(n1140), .A2(n1158), .A3(n1157), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1155), .A2(n1151), .ZN(n1158) );
INV_X1 U825 ( .A(KEYINPUT49), .ZN(n1151) );
XOR2_X1 U826 ( .A(G104), .B(n1159), .Z(G6) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U828 ( .A1(KEYINPUT52), .A2(n1162), .ZN(n1161) );
NOR2_X1 U829 ( .A1(KEYINPUT8), .A2(n1163), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1135), .A2(n1164), .ZN(G57) );
NOR2_X1 U831 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U832 ( .A(n1167), .B(KEYINPUT50), .Z(n1166) );
NAND2_X1 U833 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U834 ( .A1(n1169), .A2(n1168), .ZN(n1165) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1168) );
XNOR2_X1 U836 ( .A(n1172), .B(n1173), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1174), .B(KEYINPUT25), .Z(n1170) );
NAND2_X1 U838 ( .A1(n1144), .A2(G472), .ZN(n1174) );
NOR2_X1 U839 ( .A1(n1135), .A2(n1175), .ZN(G54) );
XOR2_X1 U840 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U841 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U842 ( .A(n1180), .B(n1181), .ZN(n1179) );
XNOR2_X1 U843 ( .A(n1182), .B(n1183), .ZN(n1178) );
NOR2_X1 U844 ( .A1(KEYINPUT61), .A2(n1184), .ZN(n1183) );
INV_X1 U845 ( .A(n1110), .ZN(n1184) );
XOR2_X1 U846 ( .A(n1185), .B(n1186), .Z(n1110) );
NOR2_X1 U847 ( .A1(G140), .A2(KEYINPUT28), .ZN(n1182) );
XOR2_X1 U848 ( .A(n1187), .B(n1188), .Z(n1176) );
XOR2_X1 U849 ( .A(KEYINPUT39), .B(G137), .Z(n1188) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1187) );
NOR2_X1 U851 ( .A1(n1191), .A2(KEYINPUT63), .ZN(n1190) );
AND2_X1 U852 ( .A1(G469), .A2(n1144), .ZN(n1191) );
NOR2_X1 U853 ( .A1(n1135), .A2(n1192), .ZN(G51) );
XOR2_X1 U854 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U855 ( .A1(KEYINPUT14), .A2(n1195), .ZN(n1194) );
XOR2_X1 U856 ( .A(n1196), .B(KEYINPUT18), .Z(n1195) );
NAND2_X1 U857 ( .A1(n1144), .A2(G210), .ZN(n1193) );
INV_X1 U858 ( .A(n1140), .ZN(n1144) );
NAND2_X1 U859 ( .A1(G902), .A2(n1051), .ZN(n1140) );
INV_X1 U860 ( .A(n1156), .ZN(n1051) );
NOR3_X1 U861 ( .A1(n1119), .A2(n1128), .A3(n1117), .ZN(n1156) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1117) );
NAND2_X1 U863 ( .A1(n1201), .A2(n1202), .ZN(n1128) );
NOR4_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR4_X1 U865 ( .A1(n1046), .A2(n1207), .A3(n1162), .A4(n1208), .ZN(n1201) );
NOR3_X1 U866 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
INV_X1 U867 ( .A(n1163), .ZN(n1162) );
NAND3_X1 U868 ( .A1(n1212), .A2(n1213), .A3(n1066), .ZN(n1163) );
INV_X1 U869 ( .A(n1214), .ZN(n1207) );
AND3_X1 U870 ( .A1(n1065), .A2(n1213), .A3(n1212), .ZN(n1046) );
INV_X1 U871 ( .A(n1058), .ZN(n1213) );
NAND4_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1119) );
NAND3_X1 U873 ( .A1(n1066), .A2(n1087), .A3(n1219), .ZN(n1215) );
AND2_X1 U874 ( .A1(n1220), .A2(n1221), .ZN(n1135) );
XOR2_X1 U875 ( .A(KEYINPUT12), .B(G953), .Z(n1221) );
XNOR2_X1 U876 ( .A(G952), .B(KEYINPUT27), .ZN(n1220) );
NAND2_X1 U877 ( .A1(n1222), .A2(n1223), .ZN(G48) );
NAND2_X1 U878 ( .A1(G146), .A2(n1197), .ZN(n1223) );
XOR2_X1 U879 ( .A(n1224), .B(KEYINPUT38), .Z(n1222) );
OR2_X1 U880 ( .A1(n1197), .A2(G146), .ZN(n1224) );
NAND2_X1 U881 ( .A1(n1225), .A2(n1066), .ZN(n1197) );
XNOR2_X1 U882 ( .A(G143), .B(n1198), .ZN(G45) );
NAND4_X1 U883 ( .A1(n1226), .A2(n1219), .A3(n1077), .A4(n1093), .ZN(n1198) );
XOR2_X1 U884 ( .A(G140), .B(n1227), .Z(G42) );
NOR2_X1 U885 ( .A1(KEYINPUT6), .A2(n1199), .ZN(n1227) );
NAND4_X1 U886 ( .A1(n1066), .A2(n1228), .A3(n1229), .A4(n1087), .ZN(n1199) );
INV_X1 U887 ( .A(n1230), .ZN(n1066) );
NAND3_X1 U888 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(G39) );
NAND2_X1 U889 ( .A1(G137), .A2(n1200), .ZN(n1233) );
NAND2_X1 U890 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
INV_X1 U891 ( .A(KEYINPUT47), .ZN(n1235) );
NAND2_X1 U892 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
INV_X1 U893 ( .A(n1200), .ZN(n1237) );
XOR2_X1 U894 ( .A(KEYINPUT3), .B(n1238), .Z(n1236) );
NAND2_X1 U895 ( .A1(KEYINPUT47), .A2(n1239), .ZN(n1231) );
NAND2_X1 U896 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
OR3_X1 U897 ( .A1(n1200), .A2(G137), .A3(KEYINPUT3), .ZN(n1241) );
NAND4_X1 U898 ( .A1(n1067), .A2(n1228), .A3(n1087), .A4(n1083), .ZN(n1200) );
NAND2_X1 U899 ( .A1(KEYINPUT3), .A2(G137), .ZN(n1240) );
XNOR2_X1 U900 ( .A(G134), .B(n1216), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1087), .A2(n1065), .A3(n1219), .ZN(n1216) );
INV_X1 U902 ( .A(n1242), .ZN(n1219) );
INV_X1 U903 ( .A(n1059), .ZN(n1087) );
XOR2_X1 U904 ( .A(G131), .B(n1243), .Z(G33) );
NOR4_X1 U905 ( .A1(KEYINPUT46), .A2(n1059), .A3(n1230), .A4(n1242), .ZN(n1243) );
NAND2_X1 U906 ( .A1(n1082), .A2(n1244), .ZN(n1242) );
NAND2_X1 U907 ( .A1(n1245), .A2(n1079), .ZN(n1059) );
INV_X1 U908 ( .A(n1078), .ZN(n1245) );
NAND2_X1 U909 ( .A1(n1246), .A2(n1247), .ZN(G30) );
NAND2_X1 U910 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U911 ( .A(KEYINPUT32), .B(n1250), .Z(n1246) );
NOR2_X1 U912 ( .A1(n1248), .A2(n1249), .ZN(n1250) );
INV_X1 U913 ( .A(n1217), .ZN(n1248) );
NAND2_X1 U914 ( .A1(n1225), .A2(n1065), .ZN(n1217) );
INV_X1 U915 ( .A(n1210), .ZN(n1065) );
AND3_X1 U916 ( .A1(n1077), .A2(n1083), .A3(n1228), .ZN(n1225) );
AND2_X1 U917 ( .A1(n1244), .A2(n1251), .ZN(n1228) );
NOR3_X1 U918 ( .A1(n1070), .A2(n1064), .A3(n1252), .ZN(n1244) );
XOR2_X1 U919 ( .A(n1253), .B(n1254), .Z(G3) );
XNOR2_X1 U920 ( .A(G101), .B(KEYINPUT54), .ZN(n1254) );
NAND2_X1 U921 ( .A1(KEYINPUT33), .A2(n1206), .ZN(n1253) );
AND3_X1 U922 ( .A1(n1067), .A2(n1212), .A3(n1082), .ZN(n1206) );
XNOR2_X1 U923 ( .A(G125), .B(n1218), .ZN(G27) );
NAND3_X1 U924 ( .A1(n1251), .A2(n1255), .A3(n1256), .ZN(n1218) );
NOR3_X1 U925 ( .A1(n1252), .A2(n1257), .A3(n1083), .ZN(n1256) );
NAND2_X1 U926 ( .A1(n1258), .A2(n1085), .ZN(n1252) );
NAND2_X1 U927 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
OR3_X1 U928 ( .A1(n1114), .A2(G900), .A3(n1261), .ZN(n1260) );
NAND3_X1 U929 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(G24) );
NAND2_X1 U930 ( .A1(n1205), .A2(n1265), .ZN(n1264) );
NAND2_X1 U931 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U932 ( .A(KEYINPUT58), .ZN(n1267) );
XOR2_X1 U933 ( .A(n1268), .B(KEYINPUT37), .Z(n1266) );
OR3_X1 U934 ( .A1(n1268), .A2(n1205), .A3(KEYINPUT58), .ZN(n1263) );
NOR4_X1 U935 ( .A1(n1269), .A2(n1209), .A3(n1058), .A4(n1270), .ZN(n1205) );
NAND2_X1 U936 ( .A1(n1229), .A2(n1084), .ZN(n1058) );
NAND2_X1 U937 ( .A1(KEYINPUT58), .A2(n1268), .ZN(n1262) );
XOR2_X1 U938 ( .A(G119), .B(n1204), .Z(G21) );
NOR4_X1 U939 ( .A1(n1209), .A2(n1071), .A3(n1084), .A4(n1229), .ZN(n1204) );
XOR2_X1 U940 ( .A(n1271), .B(n1272), .Z(G18) );
NOR2_X1 U941 ( .A1(KEYINPUT41), .A2(n1273), .ZN(n1272) );
NOR3_X1 U942 ( .A1(n1209), .A2(n1274), .A3(n1211), .ZN(n1271) );
XOR2_X1 U943 ( .A(n1210), .B(KEYINPUT15), .Z(n1274) );
NAND2_X1 U944 ( .A1(n1269), .A2(n1093), .ZN(n1210) );
NAND4_X1 U945 ( .A1(n1070), .A2(n1275), .A3(n1077), .A4(n1068), .ZN(n1209) );
INV_X1 U946 ( .A(n1257), .ZN(n1077) );
XOR2_X1 U947 ( .A(n1276), .B(n1214), .Z(G15) );
NAND4_X1 U948 ( .A1(n1255), .A2(n1082), .A3(n1277), .A4(n1275), .ZN(n1214) );
INV_X1 U949 ( .A(n1211), .ZN(n1082) );
NAND2_X1 U950 ( .A1(n1084), .A2(n1083), .ZN(n1211) );
INV_X1 U951 ( .A(n1229), .ZN(n1083) );
INV_X1 U952 ( .A(n1251), .ZN(n1084) );
NOR3_X1 U953 ( .A1(n1060), .A2(n1064), .A3(n1230), .ZN(n1255) );
NAND2_X1 U954 ( .A1(n1226), .A2(n1278), .ZN(n1230) );
XOR2_X1 U955 ( .A(KEYINPUT43), .B(n1093), .Z(n1278) );
INV_X1 U956 ( .A(n1270), .ZN(n1093) );
INV_X1 U957 ( .A(n1068), .ZN(n1064) );
XOR2_X1 U958 ( .A(G110), .B(n1203), .Z(G12) );
AND4_X1 U959 ( .A1(n1251), .A2(n1067), .A3(n1229), .A4(n1212), .ZN(n1203) );
AND4_X1 U960 ( .A1(n1277), .A2(n1275), .A3(n1060), .A4(n1068), .ZN(n1212) );
NAND2_X1 U961 ( .A1(G221), .A2(n1279), .ZN(n1068) );
INV_X1 U962 ( .A(n1070), .ZN(n1060) );
XOR2_X1 U963 ( .A(n1280), .B(n1281), .Z(n1070) );
XOR2_X1 U964 ( .A(KEYINPUT29), .B(G469), .Z(n1281) );
NAND2_X1 U965 ( .A1(n1282), .A2(n1261), .ZN(n1280) );
XOR2_X1 U966 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U967 ( .A(n1285), .B(n1286), .Z(n1284) );
INV_X1 U968 ( .A(n1185), .ZN(n1286) );
XNOR2_X1 U969 ( .A(KEYINPUT0), .B(n1287), .ZN(n1185) );
NOR2_X1 U970 ( .A1(KEYINPUT24), .A2(n1288), .ZN(n1287) );
XNOR2_X1 U971 ( .A(n1289), .B(n1181), .ZN(n1285) );
XOR2_X1 U972 ( .A(n1290), .B(n1291), .Z(n1181) );
XOR2_X1 U973 ( .A(n1292), .B(n1293), .Z(n1290) );
AND2_X1 U974 ( .A1(n1114), .A2(G227), .ZN(n1293) );
NAND2_X1 U975 ( .A1(KEYINPUT48), .A2(G101), .ZN(n1292) );
XOR2_X1 U976 ( .A(n1294), .B(n1295), .Z(n1283) );
NOR2_X1 U977 ( .A1(G140), .A2(KEYINPUT19), .ZN(n1295) );
XOR2_X1 U978 ( .A(n1189), .B(G143), .Z(n1294) );
AND2_X1 U979 ( .A1(n1296), .A2(n1085), .ZN(n1275) );
NAND2_X1 U980 ( .A1(G237), .A2(G234), .ZN(n1085) );
NAND2_X1 U981 ( .A1(n1259), .A2(n1297), .ZN(n1296) );
NAND2_X1 U982 ( .A1(G902), .A2(n1127), .ZN(n1297) );
NOR2_X1 U983 ( .A1(n1114), .A2(G898), .ZN(n1127) );
NAND2_X1 U984 ( .A1(n1298), .A2(n1114), .ZN(n1259) );
XOR2_X1 U985 ( .A(KEYINPUT34), .B(G952), .Z(n1298) );
XOR2_X1 U986 ( .A(n1257), .B(KEYINPUT22), .Z(n1277) );
NAND2_X1 U987 ( .A1(n1079), .A2(n1078), .ZN(n1257) );
NAND3_X1 U988 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1078) );
OR2_X1 U989 ( .A1(n1302), .A2(n1196), .ZN(n1301) );
NAND3_X1 U990 ( .A1(n1196), .A2(n1302), .A3(n1261), .ZN(n1300) );
NAND2_X1 U991 ( .A1(G210), .A2(G237), .ZN(n1302) );
XOR2_X1 U992 ( .A(n1303), .B(n1304), .Z(n1196) );
XNOR2_X1 U993 ( .A(n1130), .B(n1305), .ZN(n1304) );
XOR2_X1 U994 ( .A(n1306), .B(n1307), .Z(n1305) );
NOR2_X1 U995 ( .A1(n1133), .A2(n1308), .ZN(n1307) );
XOR2_X1 U996 ( .A(n1131), .B(KEYINPUT4), .Z(n1308) );
NAND2_X1 U997 ( .A1(n1309), .A2(n1310), .ZN(n1131) );
NOR2_X1 U998 ( .A1(n1310), .A2(n1309), .ZN(n1133) );
XNOR2_X1 U999 ( .A(n1311), .B(n1312), .ZN(n1309) );
XOR2_X1 U1000 ( .A(G113), .B(n1313), .Z(n1312) );
NOR2_X1 U1001 ( .A1(KEYINPUT51), .A2(n1314), .ZN(n1313) );
INV_X1 U1002 ( .A(G119), .ZN(n1314) );
XOR2_X1 U1003 ( .A(G101), .B(n1291), .Z(n1310) );
XOR2_X1 U1004 ( .A(G104), .B(G107), .Z(n1291) );
NAND2_X1 U1005 ( .A1(G224), .A2(n1114), .ZN(n1306) );
XOR2_X1 U1006 ( .A(n1189), .B(n1268), .Z(n1130) );
INV_X1 U1007 ( .A(G122), .ZN(n1268) );
INV_X1 U1008 ( .A(G110), .ZN(n1189) );
XOR2_X1 U1009 ( .A(n1315), .B(n1316), .Z(n1303) );
XOR2_X1 U1010 ( .A(G128), .B(G125), .Z(n1316) );
NAND2_X1 U1011 ( .A1(G210), .A2(G902), .ZN(n1299) );
NAND2_X1 U1012 ( .A1(n1317), .A2(G214), .ZN(n1079) );
XOR2_X1 U1013 ( .A(n1318), .B(KEYINPUT26), .Z(n1317) );
OR2_X1 U1014 ( .A1(G902), .A2(G237), .ZN(n1318) );
XOR2_X1 U1015 ( .A(n1095), .B(G472), .Z(n1229) );
NAND2_X1 U1016 ( .A1(n1319), .A2(n1261), .ZN(n1095) );
XOR2_X1 U1017 ( .A(n1320), .B(n1169), .Z(n1319) );
XOR2_X1 U1018 ( .A(n1321), .B(G101), .Z(n1169) );
NAND2_X1 U1019 ( .A1(n1322), .A2(G210), .ZN(n1321) );
NAND2_X1 U1020 ( .A1(n1323), .A2(n1324), .ZN(n1320) );
NAND2_X1 U1021 ( .A1(n1173), .A2(n1172), .ZN(n1324) );
XOR2_X1 U1022 ( .A(n1325), .B(KEYINPUT16), .Z(n1323) );
OR2_X1 U1023 ( .A1(n1172), .A2(n1173), .ZN(n1325) );
XNOR2_X1 U1024 ( .A(n1289), .B(n1315), .ZN(n1173) );
NAND2_X1 U1025 ( .A1(n1326), .A2(KEYINPUT17), .ZN(n1315) );
XOR2_X1 U1026 ( .A(G143), .B(n1288), .Z(n1326) );
XNOR2_X1 U1027 ( .A(n1327), .B(n1180), .ZN(n1289) );
XOR2_X1 U1028 ( .A(n1113), .B(KEYINPUT1), .Z(n1180) );
XOR2_X1 U1029 ( .A(G131), .B(G134), .Z(n1113) );
XNOR2_X1 U1030 ( .A(n1276), .B(n1328), .ZN(n1172) );
NOR2_X1 U1031 ( .A1(KEYINPUT56), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1032 ( .A(G119), .B(n1311), .Z(n1329) );
XNOR2_X1 U1033 ( .A(n1273), .B(KEYINPUT57), .ZN(n1311) );
INV_X1 U1034 ( .A(G113), .ZN(n1276) );
INV_X1 U1035 ( .A(n1071), .ZN(n1067) );
NAND2_X1 U1036 ( .A1(n1330), .A2(n1269), .ZN(n1071) );
INV_X1 U1037 ( .A(n1226), .ZN(n1269) );
XOR2_X1 U1038 ( .A(n1331), .B(n1153), .Z(n1226) );
INV_X1 U1039 ( .A(n1097), .ZN(n1153) );
NAND2_X1 U1040 ( .A1(n1149), .A2(n1261), .ZN(n1097) );
INV_X1 U1041 ( .A(n1155), .ZN(n1149) );
XOR2_X1 U1042 ( .A(n1332), .B(n1333), .Z(n1155) );
XOR2_X1 U1043 ( .A(G122), .B(G113), .Z(n1333) );
XOR2_X1 U1044 ( .A(n1334), .B(G104), .Z(n1332) );
NAND2_X1 U1045 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1046 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1047 ( .A(KEYINPUT35), .B(n1339), .Z(n1335) );
NOR2_X1 U1048 ( .A1(n1337), .A2(n1338), .ZN(n1339) );
NAND2_X1 U1049 ( .A1(n1340), .A2(n1341), .ZN(n1338) );
NAND2_X1 U1050 ( .A1(n1107), .A2(n1288), .ZN(n1341) );
XOR2_X1 U1051 ( .A(KEYINPUT9), .B(n1342), .Z(n1340) );
NOR2_X1 U1052 ( .A1(n1107), .A2(n1288), .ZN(n1342) );
INV_X1 U1053 ( .A(G146), .ZN(n1288) );
XOR2_X1 U1054 ( .A(n1343), .B(n1344), .Z(n1337) );
XOR2_X1 U1055 ( .A(G143), .B(G131), .Z(n1344) );
NAND3_X1 U1056 ( .A1(n1322), .A2(G214), .A3(KEYINPUT2), .ZN(n1343) );
NOR2_X1 U1057 ( .A1(G953), .A2(G237), .ZN(n1322) );
NAND2_X1 U1058 ( .A1(KEYINPUT36), .A2(n1157), .ZN(n1331) );
INV_X1 U1059 ( .A(G475), .ZN(n1157) );
XOR2_X1 U1060 ( .A(n1270), .B(KEYINPUT30), .Z(n1330) );
XOR2_X1 U1061 ( .A(n1345), .B(G478), .Z(n1270) );
NAND2_X1 U1062 ( .A1(n1143), .A2(n1261), .ZN(n1345) );
XNOR2_X1 U1063 ( .A(n1346), .B(n1347), .ZN(n1143) );
AND2_X1 U1064 ( .A1(n1348), .A2(G217), .ZN(n1347) );
NAND3_X1 U1065 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1346) );
OR2_X1 U1066 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND3_X1 U1067 ( .A1(n1354), .A2(n1352), .A3(n1355), .ZN(n1350) );
INV_X1 U1068 ( .A(KEYINPUT7), .ZN(n1352) );
OR2_X1 U1069 ( .A1(n1355), .A2(n1354), .ZN(n1349) );
AND2_X1 U1070 ( .A1(KEYINPUT44), .A2(n1353), .ZN(n1354) );
XOR2_X1 U1071 ( .A(n1186), .B(n1356), .Z(n1353) );
NOR2_X1 U1072 ( .A1(G134), .A2(KEYINPUT60), .ZN(n1356) );
XOR2_X1 U1073 ( .A(G128), .B(G143), .Z(n1186) );
XNOR2_X1 U1074 ( .A(n1357), .B(n1358), .ZN(n1355) );
NOR2_X1 U1075 ( .A1(G122), .A2(KEYINPUT55), .ZN(n1358) );
XOR2_X1 U1076 ( .A(G107), .B(n1273), .Z(n1357) );
INV_X1 U1077 ( .A(G116), .ZN(n1273) );
XNOR2_X1 U1078 ( .A(n1092), .B(KEYINPUT23), .ZN(n1251) );
XNOR2_X1 U1079 ( .A(n1359), .B(n1360), .ZN(n1092) );
AND2_X1 U1080 ( .A1(n1279), .A2(G217), .ZN(n1360) );
NAND2_X1 U1081 ( .A1(G234), .A2(n1261), .ZN(n1279) );
INV_X1 U1082 ( .A(G902), .ZN(n1261) );
NAND2_X1 U1083 ( .A1(n1361), .A2(n1137), .ZN(n1359) );
XNOR2_X1 U1084 ( .A(n1362), .B(n1363), .ZN(n1137) );
XOR2_X1 U1085 ( .A(G110), .B(n1364), .Z(n1363) );
XOR2_X1 U1086 ( .A(G146), .B(G119), .Z(n1364) );
XOR2_X1 U1087 ( .A(n1365), .B(n1327), .Z(n1362) );
XOR2_X1 U1088 ( .A(n1249), .B(n1238), .Z(n1327) );
INV_X1 U1089 ( .A(G137), .ZN(n1238) );
INV_X1 U1090 ( .A(G128), .ZN(n1249) );
XNOR2_X1 U1091 ( .A(n1366), .B(n1107), .ZN(n1365) );
XNOR2_X1 U1092 ( .A(G125), .B(G140), .ZN(n1107) );
NAND2_X1 U1093 ( .A1(n1348), .A2(G221), .ZN(n1366) );
AND2_X1 U1094 ( .A1(G234), .A2(n1114), .ZN(n1348) );
INV_X1 U1095 ( .A(G953), .ZN(n1114) );
XOR2_X1 U1096 ( .A(KEYINPUT62), .B(G902), .Z(n1361) );
endmodule


