//Key = 1110000001101111011101101000100000111101110110100100110100100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309;

XNOR2_X1 U726 ( .A(n1009), .B(n1010), .ZN(G9) );
NAND3_X1 U727 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(G75) );
NAND2_X1 U728 ( .A1(G952), .A2(n1014), .ZN(n1013) );
NAND3_X1 U729 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND2_X1 U730 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NAND2_X1 U731 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND4_X1 U732 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
NAND2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1020) );
NAND2_X1 U734 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U735 ( .A1(n1025), .A2(n1030), .A3(n1022), .ZN(n1029) );
NAND2_X1 U736 ( .A1(n1024), .A2(n1031), .ZN(n1028) );
NAND2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U738 ( .A1(n1022), .A2(n1034), .ZN(n1033) );
NAND2_X1 U739 ( .A1(n1025), .A2(n1035), .ZN(n1032) );
INV_X1 U740 ( .A(n1036), .ZN(n1018) );
XOR2_X1 U741 ( .A(KEYINPUT5), .B(n1037), .Z(n1015) );
NOR2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR4_X1 U743 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1036), .ZN(n1039) );
NOR2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
NOR2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR3_X1 U746 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1043) );
NOR4_X1 U747 ( .A1(n1050), .A2(n1049), .A3(n1046), .A4(n1036), .ZN(n1038) );
XNOR2_X1 U748 ( .A(n1051), .B(KEYINPUT20), .ZN(n1036) );
NOR2_X1 U749 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
AND3_X1 U750 ( .A1(n1054), .A2(n1025), .A3(n1055), .ZN(n1052) );
NAND4_X1 U751 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1011) );
NOR4_X1 U752 ( .A1(n1060), .A2(n1054), .A3(n1061), .A4(n1062), .ZN(n1059) );
NOR2_X1 U753 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U754 ( .A1(G902), .A2(n1065), .ZN(n1063) );
NOR2_X1 U755 ( .A1(n1066), .A2(n1049), .ZN(n1058) );
INV_X1 U756 ( .A(n1026), .ZN(n1049) );
XOR2_X1 U757 ( .A(n1067), .B(n1068), .Z(n1066) );
XNOR2_X1 U758 ( .A(KEYINPUT28), .B(n1069), .ZN(n1068) );
XOR2_X1 U759 ( .A(n1070), .B(n1071), .Z(n1057) );
NAND2_X1 U760 ( .A1(KEYINPUT35), .A2(n1072), .ZN(n1070) );
XNOR2_X1 U761 ( .A(n1073), .B(n1074), .ZN(n1056) );
XNOR2_X1 U762 ( .A(KEYINPUT63), .B(KEYINPUT17), .ZN(n1073) );
XOR2_X1 U763 ( .A(n1075), .B(n1076), .Z(G72) );
XOR2_X1 U764 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U766 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U767 ( .A(n1083), .B(n1084), .Z(n1082) );
XNOR2_X1 U768 ( .A(n1085), .B(G131), .ZN(n1084) );
XOR2_X1 U769 ( .A(KEYINPUT25), .B(KEYINPUT16), .Z(n1083) );
XNOR2_X1 U770 ( .A(n1086), .B(n1087), .ZN(n1081) );
XOR2_X1 U771 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U772 ( .A1(KEYINPUT41), .A2(n1090), .ZN(n1089) );
NAND2_X1 U773 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U774 ( .A1(G137), .A2(n1093), .ZN(n1092) );
XOR2_X1 U775 ( .A(n1094), .B(KEYINPUT47), .Z(n1091) );
OR2_X1 U776 ( .A1(n1093), .A2(G137), .ZN(n1094) );
NOR2_X1 U777 ( .A1(G900), .A2(n1012), .ZN(n1079) );
NAND3_X1 U778 ( .A1(n1095), .A2(n1096), .A3(KEYINPUT58), .ZN(n1077) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1096) );
NAND2_X1 U780 ( .A1(n1012), .A2(n1097), .ZN(n1075) );
XOR2_X1 U781 ( .A(n1098), .B(n1099), .Z(G69) );
NOR2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U783 ( .A(n1095), .ZN(n1101) );
XOR2_X1 U784 ( .A(G953), .B(KEYINPUT57), .Z(n1095) );
NOR2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND3_X1 U786 ( .A1(n1104), .A2(n1105), .A3(KEYINPUT13), .ZN(n1098) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1012), .ZN(n1105) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND3_X1 U789 ( .A1(n1107), .A2(G898), .A3(G953), .ZN(n1104) );
NOR2_X1 U790 ( .A1(KEYINPUT42), .A2(n1109), .ZN(n1107) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
XOR2_X1 U795 ( .A(n1115), .B(KEYINPUT49), .Z(n1116) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U797 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U798 ( .A1(KEYINPUT0), .A2(n1122), .ZN(n1120) );
NAND2_X1 U799 ( .A1(n1123), .A2(n1071), .ZN(n1122) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U801 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U802 ( .A1(G478), .A2(n1123), .ZN(n1125) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1127), .ZN(G60) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
AND2_X1 U805 ( .A1(G475), .A2(n1123), .ZN(n1128) );
XOR2_X1 U806 ( .A(G104), .B(n1130), .Z(G6) );
NOR2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U808 ( .A1(n1118), .A2(n1133), .ZN(G57) );
XNOR2_X1 U809 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U810 ( .A(n1136), .B(n1137), .Z(n1134) );
NAND2_X1 U811 ( .A1(n1123), .A2(G472), .ZN(n1136) );
NOR2_X1 U812 ( .A1(n1118), .A2(n1138), .ZN(G54) );
XOR2_X1 U813 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U814 ( .A(n1141), .B(n1142), .Z(n1139) );
NOR2_X1 U815 ( .A1(KEYINPUT26), .A2(n1143), .ZN(n1142) );
NAND2_X1 U816 ( .A1(n1123), .A2(G469), .ZN(n1141) );
NOR3_X1 U817 ( .A1(n1118), .A2(n1144), .A3(n1145), .ZN(G51) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U819 ( .A(n1148), .B(n1149), .Z(n1146) );
NOR2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
INV_X1 U821 ( .A(KEYINPUT40), .ZN(n1151) );
NOR2_X1 U822 ( .A1(n1152), .A2(n1153), .ZN(n1144) );
XOR2_X1 U823 ( .A(n1148), .B(n1154), .Z(n1153) );
AND2_X1 U824 ( .A1(n1150), .A2(KEYINPUT40), .ZN(n1154) );
AND2_X1 U825 ( .A1(n1123), .A2(n1155), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1017), .ZN(n1123) );
NOR2_X1 U827 ( .A1(n1108), .A2(n1097), .ZN(n1017) );
NAND4_X1 U828 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1097) );
AND4_X1 U829 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND3_X1 U830 ( .A1(n1165), .A2(n1023), .A3(n1053), .ZN(n1159) );
NAND2_X1 U831 ( .A1(n1022), .A2(n1166), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XNOR2_X1 U833 ( .A(n1169), .B(KEYINPUT50), .ZN(n1167) );
NAND4_X1 U834 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1108) );
NOR4_X1 U835 ( .A1(n1174), .A2(n1175), .A3(n1010), .A4(n1176), .ZN(n1173) );
INV_X1 U836 ( .A(n1177), .ZN(n1176) );
NOR2_X1 U837 ( .A1(n1045), .A2(n1131), .ZN(n1010) );
NAND2_X1 U838 ( .A1(n1178), .A2(n1025), .ZN(n1131) );
INV_X1 U839 ( .A(n1179), .ZN(n1045) );
NOR4_X1 U840 ( .A1(n1180), .A2(n1181), .A3(n1041), .A4(n1132), .ZN(n1175) );
INV_X1 U841 ( .A(n1025), .ZN(n1041) );
NOR2_X1 U842 ( .A1(KEYINPUT43), .A2(n1182), .ZN(n1181) );
NOR3_X1 U843 ( .A1(n1183), .A2(n1035), .A3(n1184), .ZN(n1182) );
NOR2_X1 U844 ( .A1(n1178), .A2(n1185), .ZN(n1180) );
INV_X1 U845 ( .A(KEYINPUT43), .ZN(n1185) );
NOR2_X1 U846 ( .A1(n1186), .A2(n1187), .ZN(n1172) );
INV_X1 U847 ( .A(n1147), .ZN(n1152) );
NAND2_X1 U848 ( .A1(KEYINPUT24), .A2(n1188), .ZN(n1147) );
XOR2_X1 U849 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U850 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U851 ( .A1(KEYINPUT54), .A2(n1090), .ZN(n1192) );
NOR2_X1 U852 ( .A1(n1012), .A2(G952), .ZN(n1118) );
XNOR2_X1 U853 ( .A(G146), .B(n1158), .ZN(G48) );
NAND2_X1 U854 ( .A1(n1193), .A2(n1023), .ZN(n1158) );
XOR2_X1 U855 ( .A(n1164), .B(n1194), .Z(G45) );
XNOR2_X1 U856 ( .A(G143), .B(KEYINPUT38), .ZN(n1194) );
NAND4_X1 U857 ( .A1(n1195), .A2(n1035), .A3(n1196), .A4(n1197), .ZN(n1164) );
XNOR2_X1 U858 ( .A(G140), .B(n1198), .ZN(G42) );
NAND3_X1 U859 ( .A1(n1053), .A2(n1165), .A3(n1199), .ZN(n1198) );
XNOR2_X1 U860 ( .A(n1023), .B(KEYINPUT18), .ZN(n1199) );
AND3_X1 U861 ( .A1(n1200), .A2(n1201), .A3(n1022), .ZN(n1053) );
XNOR2_X1 U862 ( .A(G137), .B(n1202), .ZN(G39) );
NAND2_X1 U863 ( .A1(n1169), .A2(n1022), .ZN(n1202) );
AND2_X1 U864 ( .A1(n1165), .A2(n1203), .ZN(n1169) );
XNOR2_X1 U865 ( .A(n1093), .B(n1204), .ZN(G36) );
NOR3_X1 U866 ( .A1(n1042), .A2(KEYINPUT32), .A3(n1205), .ZN(n1204) );
XOR2_X1 U867 ( .A(n1168), .B(KEYINPUT27), .Z(n1205) );
NAND2_X1 U868 ( .A1(n1195), .A2(n1179), .ZN(n1168) );
XNOR2_X1 U869 ( .A(n1206), .B(n1163), .ZN(G33) );
NAND3_X1 U870 ( .A1(n1195), .A2(n1023), .A3(n1022), .ZN(n1163) );
INV_X1 U871 ( .A(n1042), .ZN(n1022) );
NAND2_X1 U872 ( .A1(n1055), .A2(n1207), .ZN(n1042) );
AND2_X1 U873 ( .A1(n1165), .A2(n1034), .ZN(n1195) );
NAND2_X1 U874 ( .A1(KEYINPUT53), .A2(n1208), .ZN(n1206) );
XOR2_X1 U875 ( .A(G128), .B(n1209), .Z(G30) );
NOR2_X1 U876 ( .A1(KEYINPUT45), .A2(n1162), .ZN(n1209) );
NAND2_X1 U877 ( .A1(n1193), .A2(n1179), .ZN(n1162) );
AND4_X1 U878 ( .A1(n1074), .A2(n1165), .A3(n1035), .A4(n1201), .ZN(n1193) );
AND2_X1 U879 ( .A1(n1030), .A2(n1210), .ZN(n1165) );
INV_X1 U880 ( .A(n1183), .ZN(n1030) );
XOR2_X1 U881 ( .A(G101), .B(n1174), .Z(G3) );
AND3_X1 U882 ( .A1(n1026), .A2(n1178), .A3(n1034), .ZN(n1174) );
XOR2_X1 U883 ( .A(n1161), .B(n1211), .Z(G27) );
XOR2_X1 U884 ( .A(KEYINPUT9), .B(G125), .Z(n1211) );
NAND4_X1 U885 ( .A1(n1201), .A2(n1210), .A3(n1200), .A4(n1212), .ZN(n1161) );
NOR3_X1 U886 ( .A1(n1132), .A2(n1213), .A3(n1046), .ZN(n1212) );
NAND2_X1 U887 ( .A1(n1214), .A2(n1215), .ZN(n1210) );
NAND2_X1 U888 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
INV_X1 U889 ( .A(G900), .ZN(n1217) );
XNOR2_X1 U890 ( .A(G122), .B(n1170), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1218), .A2(n1025), .A3(n1196), .A4(n1197), .ZN(n1170) );
NOR2_X1 U892 ( .A1(n1201), .A2(n1074), .ZN(n1025) );
XNOR2_X1 U893 ( .A(G119), .B(n1171), .ZN(G21) );
NAND2_X1 U894 ( .A1(n1203), .A2(n1218), .ZN(n1171) );
AND3_X1 U895 ( .A1(n1074), .A2(n1201), .A3(n1026), .ZN(n1203) );
XNOR2_X1 U896 ( .A(n1219), .B(n1220), .ZN(G18) );
NOR2_X1 U897 ( .A1(KEYINPUT56), .A2(n1177), .ZN(n1220) );
NAND3_X1 U898 ( .A1(n1034), .A2(n1179), .A3(n1218), .ZN(n1177) );
NOR2_X1 U899 ( .A1(n1197), .A2(n1221), .ZN(n1179) );
XNOR2_X1 U900 ( .A(G113), .B(n1222), .ZN(G15) );
NAND2_X1 U901 ( .A1(KEYINPUT1), .A2(n1187), .ZN(n1222) );
AND3_X1 U902 ( .A1(n1218), .A2(n1034), .A3(n1023), .ZN(n1187) );
INV_X1 U903 ( .A(n1132), .ZN(n1023) );
NAND2_X1 U904 ( .A1(n1221), .A2(n1197), .ZN(n1132) );
INV_X1 U905 ( .A(n1196), .ZN(n1221) );
AND2_X1 U906 ( .A1(n1074), .A2(n1223), .ZN(n1034) );
XOR2_X1 U907 ( .A(KEYINPUT55), .B(n1201), .Z(n1223) );
INV_X1 U908 ( .A(n1200), .ZN(n1074) );
NOR3_X1 U909 ( .A1(n1213), .A2(n1184), .A3(n1046), .ZN(n1218) );
INV_X1 U910 ( .A(n1024), .ZN(n1046) );
NOR2_X1 U911 ( .A1(n1048), .A2(n1061), .ZN(n1024) );
INV_X1 U912 ( .A(n1047), .ZN(n1061) );
NAND2_X1 U913 ( .A1(n1224), .A2(n1225), .ZN(G12) );
NAND2_X1 U914 ( .A1(n1186), .A2(n1226), .ZN(n1225) );
XOR2_X1 U915 ( .A(KEYINPUT10), .B(n1227), .Z(n1224) );
NOR2_X1 U916 ( .A1(n1186), .A2(n1226), .ZN(n1227) );
INV_X1 U917 ( .A(G110), .ZN(n1226) );
AND4_X1 U918 ( .A1(n1026), .A2(n1178), .A3(n1200), .A4(n1201), .ZN(n1186) );
XOR2_X1 U919 ( .A(n1072), .B(n1071), .Z(n1201) );
AND2_X1 U920 ( .A1(G217), .A2(n1228), .ZN(n1071) );
NOR2_X1 U921 ( .A1(n1121), .A2(G902), .ZN(n1072) );
XOR2_X1 U922 ( .A(n1229), .B(n1230), .Z(n1121) );
XOR2_X1 U923 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U924 ( .A(G128), .B(G119), .Z(n1232) );
XOR2_X1 U925 ( .A(KEYINPUT51), .B(G137), .Z(n1231) );
XOR2_X1 U926 ( .A(n1233), .B(n1234), .Z(n1229) );
AND3_X1 U927 ( .A1(G221), .A2(n1012), .A3(G234), .ZN(n1234) );
XNOR2_X1 U928 ( .A(G110), .B(n1235), .ZN(n1233) );
NOR2_X1 U929 ( .A1(KEYINPUT59), .A2(n1236), .ZN(n1235) );
XOR2_X1 U930 ( .A(n1237), .B(n1238), .Z(n1236) );
NAND2_X1 U931 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
NAND2_X1 U932 ( .A1(n1241), .A2(n1085), .ZN(n1240) );
XOR2_X1 U933 ( .A(KEYINPUT14), .B(n1242), .Z(n1239) );
NOR2_X1 U934 ( .A1(n1241), .A2(n1085), .ZN(n1242) );
XNOR2_X1 U935 ( .A(n1243), .B(n1244), .ZN(n1200) );
XOR2_X1 U936 ( .A(KEYINPUT19), .B(G472), .Z(n1244) );
NAND2_X1 U937 ( .A1(n1245), .A2(n1156), .ZN(n1243) );
XOR2_X1 U938 ( .A(n1246), .B(n1137), .Z(n1245) );
XNOR2_X1 U939 ( .A(n1247), .B(G101), .ZN(n1137) );
NAND2_X1 U940 ( .A1(G210), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U941 ( .A(KEYINPUT36), .B(n1249), .ZN(n1246) );
NOR2_X1 U942 ( .A1(KEYINPUT6), .A2(n1135), .ZN(n1249) );
XOR2_X1 U943 ( .A(n1250), .B(n1251), .Z(n1135) );
XNOR2_X1 U944 ( .A(G113), .B(n1252), .ZN(n1251) );
XNOR2_X1 U945 ( .A(KEYINPUT30), .B(KEYINPUT21), .ZN(n1252) );
XOR2_X1 U946 ( .A(n1253), .B(n1254), .Z(n1250) );
XNOR2_X1 U947 ( .A(n1255), .B(n1189), .ZN(n1253) );
NOR3_X1 U948 ( .A1(n1183), .A2(n1184), .A3(n1213), .ZN(n1178) );
INV_X1 U949 ( .A(n1035), .ZN(n1213) );
NOR2_X1 U950 ( .A1(n1054), .A2(n1055), .ZN(n1035) );
NOR2_X1 U951 ( .A1(n1256), .A2(n1060), .ZN(n1055) );
NOR3_X1 U952 ( .A1(n1155), .A2(G902), .A3(n1065), .ZN(n1060) );
INV_X1 U953 ( .A(n1064), .ZN(n1155) );
AND2_X1 U954 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
OR2_X1 U955 ( .A1(n1065), .A2(G902), .ZN(n1258) );
XNOR2_X1 U956 ( .A(n1259), .B(n1260), .ZN(n1065) );
XNOR2_X1 U957 ( .A(n1090), .B(n1150), .ZN(n1260) );
XOR2_X1 U958 ( .A(n1111), .B(n1261), .Z(n1150) );
NOR2_X1 U959 ( .A1(KEYINPUT8), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U960 ( .A(n1115), .B(n1117), .ZN(n1262) );
INV_X1 U961 ( .A(n1114), .ZN(n1117) );
XNOR2_X1 U962 ( .A(n1263), .B(n1264), .ZN(n1114) );
XNOR2_X1 U963 ( .A(KEYINPUT12), .B(n1265), .ZN(n1263) );
NOR2_X1 U964 ( .A1(KEYINPUT23), .A2(n1009), .ZN(n1265) );
INV_X1 U965 ( .A(G107), .ZN(n1009) );
NAND2_X1 U966 ( .A1(n1266), .A2(n1267), .ZN(n1115) );
NAND2_X1 U967 ( .A1(n1268), .A2(n1255), .ZN(n1267) );
XOR2_X1 U968 ( .A(n1269), .B(KEYINPUT3), .Z(n1266) );
OR2_X1 U969 ( .A1(n1255), .A2(n1268), .ZN(n1269) );
XOR2_X1 U970 ( .A(G113), .B(KEYINPUT4), .Z(n1268) );
XOR2_X1 U971 ( .A(G116), .B(n1270), .Z(n1255) );
XOR2_X1 U972 ( .A(KEYINPUT33), .B(G119), .Z(n1270) );
XNOR2_X1 U973 ( .A(G110), .B(G122), .ZN(n1111) );
XOR2_X1 U974 ( .A(n1271), .B(n1189), .Z(n1259) );
XNOR2_X1 U975 ( .A(n1272), .B(KEYINPUT22), .ZN(n1189) );
INV_X1 U976 ( .A(n1086), .ZN(n1272) );
XOR2_X1 U977 ( .A(n1273), .B(KEYINPUT52), .Z(n1271) );
NAND2_X1 U978 ( .A1(KEYINPUT62), .A2(n1191), .ZN(n1273) );
NOR2_X1 U979 ( .A1(n1102), .A2(G953), .ZN(n1191) );
INV_X1 U980 ( .A(G224), .ZN(n1102) );
XNOR2_X1 U981 ( .A(KEYINPUT60), .B(n1064), .ZN(n1257) );
NAND2_X1 U982 ( .A1(G210), .A2(n1274), .ZN(n1064) );
INV_X1 U983 ( .A(n1207), .ZN(n1054) );
NAND2_X1 U984 ( .A1(G214), .A2(n1274), .ZN(n1207) );
NAND2_X1 U985 ( .A1(n1275), .A2(n1156), .ZN(n1274) );
INV_X1 U986 ( .A(G237), .ZN(n1275) );
AND2_X1 U987 ( .A1(n1214), .A2(n1276), .ZN(n1184) );
NAND2_X1 U988 ( .A1(n1216), .A2(n1103), .ZN(n1276) );
INV_X1 U989 ( .A(G898), .ZN(n1103) );
AND3_X1 U990 ( .A1(G902), .A2(n1051), .A3(G953), .ZN(n1216) );
NAND3_X1 U991 ( .A1(n1051), .A2(n1012), .A3(G952), .ZN(n1214) );
NAND2_X1 U992 ( .A1(G237), .A2(n1277), .ZN(n1051) );
NAND2_X1 U993 ( .A1(n1048), .A2(n1047), .ZN(n1183) );
NAND2_X1 U994 ( .A1(G221), .A2(n1228), .ZN(n1047) );
NAND2_X1 U995 ( .A1(n1277), .A2(n1156), .ZN(n1228) );
XNOR2_X1 U996 ( .A(G234), .B(KEYINPUT61), .ZN(n1277) );
XNOR2_X1 U997 ( .A(n1278), .B(n1067), .ZN(n1048) );
NAND2_X1 U998 ( .A1(n1279), .A2(n1156), .ZN(n1067) );
INV_X1 U999 ( .A(G902), .ZN(n1156) );
XOR2_X1 U1000 ( .A(n1143), .B(n1280), .Z(n1279) );
XNOR2_X1 U1001 ( .A(n1140), .B(KEYINPUT11), .ZN(n1280) );
XNOR2_X1 U1002 ( .A(n1281), .B(n1282), .ZN(n1140) );
XNOR2_X1 U1003 ( .A(n1085), .B(G110), .ZN(n1282) );
XOR2_X1 U1004 ( .A(n1283), .B(n1254), .Z(n1281) );
XNOR2_X1 U1005 ( .A(n1284), .B(n1285), .ZN(n1254) );
XOR2_X1 U1006 ( .A(KEYINPUT15), .B(G137), .Z(n1285) );
XNOR2_X1 U1007 ( .A(G131), .B(G134), .ZN(n1284) );
NAND2_X1 U1008 ( .A1(G227), .A2(n1012), .ZN(n1283) );
XOR2_X1 U1009 ( .A(n1286), .B(n1264), .Z(n1143) );
XOR2_X1 U1010 ( .A(G101), .B(G104), .Z(n1264) );
XNOR2_X1 U1011 ( .A(G107), .B(n1086), .ZN(n1286) );
XNOR2_X1 U1012 ( .A(n1287), .B(n1288), .ZN(n1086) );
XNOR2_X1 U1013 ( .A(G146), .B(KEYINPUT46), .ZN(n1287) );
NAND2_X1 U1014 ( .A1(KEYINPUT2), .A2(n1069), .ZN(n1278) );
INV_X1 U1015 ( .A(G469), .ZN(n1069) );
NOR2_X1 U1016 ( .A1(n1196), .A2(n1197), .ZN(n1026) );
XNOR2_X1 U1017 ( .A(n1289), .B(G475), .ZN(n1197) );
OR2_X1 U1018 ( .A1(n1129), .A2(G902), .ZN(n1289) );
XNOR2_X1 U1019 ( .A(n1290), .B(n1291), .ZN(n1129) );
XOR2_X1 U1020 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U1021 ( .A(G122), .B(G113), .Z(n1293) );
XNOR2_X1 U1022 ( .A(KEYINPUT34), .B(n1085), .ZN(n1292) );
INV_X1 U1023 ( .A(G140), .ZN(n1085) );
XOR2_X1 U1024 ( .A(n1294), .B(n1295), .Z(n1290) );
XOR2_X1 U1025 ( .A(G104), .B(n1296), .Z(n1295) );
NOR2_X1 U1026 ( .A1(KEYINPUT48), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1027 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U1028 ( .A(G143), .B(n1300), .ZN(n1299) );
NAND2_X1 U1029 ( .A1(n1248), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1030 ( .A(KEYINPUT29), .B(G214), .Z(n1301) );
NOR2_X1 U1031 ( .A1(G953), .A2(G237), .ZN(n1248) );
NOR2_X1 U1032 ( .A1(KEYINPUT31), .A2(n1208), .ZN(n1298) );
INV_X1 U1033 ( .A(G131), .ZN(n1208) );
XNOR2_X1 U1034 ( .A(n1238), .B(n1241), .ZN(n1294) );
INV_X1 U1035 ( .A(n1090), .ZN(n1241) );
XOR2_X1 U1036 ( .A(G125), .B(KEYINPUT37), .Z(n1090) );
XNOR2_X1 U1037 ( .A(G146), .B(KEYINPUT7), .ZN(n1238) );
XNOR2_X1 U1038 ( .A(n1302), .B(G478), .ZN(n1196) );
OR2_X1 U1039 ( .A1(n1126), .A2(G902), .ZN(n1302) );
XNOR2_X1 U1040 ( .A(n1303), .B(n1304), .ZN(n1126) );
XOR2_X1 U1041 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1042 ( .A(G107), .B(G122), .ZN(n1306) );
NAND3_X1 U1043 ( .A1(G217), .A2(n1012), .A3(G234), .ZN(n1305) );
INV_X1 U1044 ( .A(G953), .ZN(n1012) );
XNOR2_X1 U1045 ( .A(n1307), .B(n1308), .ZN(n1303) );
NAND2_X1 U1046 ( .A1(KEYINPUT39), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1047 ( .A(n1093), .B(n1288), .ZN(n1309) );
XOR2_X1 U1048 ( .A(G128), .B(G143), .Z(n1288) );
INV_X1 U1049 ( .A(G134), .ZN(n1093) );
NAND2_X1 U1050 ( .A1(KEYINPUT44), .A2(n1219), .ZN(n1307) );
INV_X1 U1051 ( .A(G116), .ZN(n1219) );
endmodule


