//Key = 1101011111010111101001100010011001011111110100010000011000011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321;

XNOR2_X1 U731 ( .A(G107), .B(n1008), .ZN(G9) );
NAND2_X1 U732 ( .A1(KEYINPUT22), .A2(n1009), .ZN(n1008) );
NOR2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U734 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NOR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND4_X1 U736 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1012) );
NAND3_X1 U737 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1019) );
XNOR2_X1 U738 ( .A(KEYINPUT28), .B(n1017), .ZN(n1023) );
NAND3_X1 U739 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1017) );
NAND2_X1 U740 ( .A1(n1028), .A2(n1029), .ZN(n1018) );
NAND3_X1 U741 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
XOR2_X1 U742 ( .A(KEYINPUT16), .B(n1033), .Z(n1032) );
NOR2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND4_X1 U744 ( .A1(n1025), .A2(n1036), .A3(n1026), .A4(n1037), .ZN(n1031) );
NAND2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
OR2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1027), .A2(n1050), .ZN(n1030) );
INV_X1 U752 ( .A(n1035), .ZN(n1027) );
NAND3_X1 U753 ( .A1(n1040), .A2(n1044), .A3(n1036), .ZN(n1035) );
INV_X1 U754 ( .A(n1051), .ZN(n1036) );
INV_X1 U755 ( .A(n1052), .ZN(n1028) );
NOR3_X1 U756 ( .A1(n1053), .A2(G953), .A3(G952), .ZN(n1010) );
INV_X1 U757 ( .A(n1020), .ZN(n1053) );
NAND4_X1 U758 ( .A1(n1054), .A2(n1048), .A3(n1025), .A4(n1055), .ZN(n1020) );
NOR3_X1 U759 ( .A1(n1056), .A2(n1052), .A3(n1057), .ZN(n1055) );
XNOR2_X1 U760 ( .A(n1026), .B(n1058), .ZN(n1056) );
XOR2_X1 U761 ( .A(KEYINPUT45), .B(KEYINPUT42), .Z(n1058) );
XNOR2_X1 U762 ( .A(G469), .B(n1059), .ZN(n1054) );
NAND2_X1 U763 ( .A1(KEYINPUT63), .A2(n1060), .ZN(n1059) );
XOR2_X1 U764 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XOR2_X1 U767 ( .A(KEYINPUT40), .B(n1067), .Z(n1066) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
NOR3_X1 U769 ( .A1(n1069), .A2(n1068), .A3(n1067), .ZN(n1063) );
AND2_X1 U770 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NAND2_X1 U771 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U772 ( .A(n1074), .B(n1075), .Z(n1070) );
XOR2_X1 U773 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U774 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U775 ( .A1(KEYINPUT8), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U776 ( .A(n1081), .B(n1082), .ZN(n1074) );
XOR2_X1 U777 ( .A(KEYINPUT17), .B(G134), .Z(n1082) );
XNOR2_X1 U778 ( .A(n1021), .B(KEYINPUT62), .ZN(n1069) );
NAND2_X1 U779 ( .A1(G953), .A2(n1083), .ZN(n1061) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1083) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(G69) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U783 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U786 ( .A1(n1073), .A2(n1091), .ZN(n1090) );
NOR2_X1 U787 ( .A1(n1092), .A2(G953), .ZN(n1084) );
NOR2_X1 U788 ( .A1(n1093), .A2(n1094), .ZN(G66) );
XNOR2_X1 U789 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1093), .A2(n1099), .ZN(G63) );
XOR2_X1 U792 ( .A(n1100), .B(n1101), .Z(n1099) );
AND2_X1 U793 ( .A1(G478), .A2(n1102), .ZN(n1100) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1103), .ZN(G60) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND3_X1 U796 ( .A1(n1102), .A2(G475), .A3(KEYINPUT37), .ZN(n1104) );
XOR2_X1 U797 ( .A(n1106), .B(n1107), .Z(G6) );
NAND2_X1 U798 ( .A1(KEYINPUT35), .A2(n1108), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1093), .A2(n1109), .ZN(G57) );
XOR2_X1 U800 ( .A(n1110), .B(n1111), .Z(n1109) );
XNOR2_X1 U801 ( .A(n1112), .B(n1113), .ZN(n1111) );
NOR2_X1 U802 ( .A1(KEYINPUT31), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U803 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND3_X1 U804 ( .A1(n1102), .A2(G472), .A3(KEYINPUT3), .ZN(n1112) );
XNOR2_X1 U805 ( .A(n1117), .B(n1118), .ZN(n1110) );
NOR2_X1 U806 ( .A1(n1093), .A2(n1119), .ZN(G54) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1122) );
NOR2_X1 U810 ( .A1(G110), .A2(KEYINPUT48), .ZN(n1125) );
NAND2_X1 U811 ( .A1(KEYINPUT18), .A2(n1076), .ZN(n1124) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(n1120) );
AND2_X1 U813 ( .A1(G469), .A2(n1102), .ZN(n1127) );
XNOR2_X1 U814 ( .A(G140), .B(n1128), .ZN(n1126) );
NOR3_X1 U815 ( .A1(n1129), .A2(KEYINPUT20), .A3(G953), .ZN(n1128) );
INV_X1 U816 ( .A(G227), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1093), .A2(n1130), .ZN(G51) );
XOR2_X1 U818 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U819 ( .A1(G210), .A2(n1102), .ZN(n1132) );
INV_X1 U820 ( .A(n1098), .ZN(n1102) );
NAND2_X1 U821 ( .A1(G902), .A2(n1133), .ZN(n1098) );
NAND2_X1 U822 ( .A1(n1092), .A2(n1068), .ZN(n1133) );
INV_X1 U823 ( .A(n1015), .ZN(n1068) );
NAND4_X1 U824 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1015) );
NOR4_X1 U825 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
NOR2_X1 U826 ( .A1(KEYINPUT4), .A2(n1142), .ZN(n1141) );
NOR2_X1 U827 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
INV_X1 U828 ( .A(n1145), .ZN(n1144) );
NOR2_X1 U829 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
NOR2_X1 U830 ( .A1(n1057), .A2(n1148), .ZN(n1147) );
INV_X1 U831 ( .A(n1044), .ZN(n1057) );
NOR3_X1 U832 ( .A1(n1149), .A2(n1043), .A3(n1150), .ZN(n1146) );
INV_X1 U833 ( .A(KEYINPUT4), .ZN(n1150) );
INV_X1 U834 ( .A(n1151), .ZN(n1043) );
NAND3_X1 U835 ( .A1(n1152), .A2(n1046), .A3(n1153), .ZN(n1149) );
NOR3_X1 U836 ( .A1(n1148), .A2(n1042), .A3(n1034), .ZN(n1139) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1155), .ZN(n1136) );
INV_X1 U838 ( .A(n1013), .ZN(n1092) );
NAND4_X1 U839 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1013) );
NOR4_X1 U840 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1107), .ZN(n1159) );
AND3_X1 U841 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1107) );
NOR2_X1 U842 ( .A1(n1009), .A2(n1166), .ZN(n1158) );
INV_X1 U843 ( .A(n1167), .ZN(n1166) );
AND3_X1 U844 ( .A1(n1163), .A2(n1164), .A3(n1151), .ZN(n1009) );
NOR2_X1 U845 ( .A1(n1168), .A2(n1169), .ZN(n1131) );
XOR2_X1 U846 ( .A(KEYINPUT56), .B(n1170), .Z(n1169) );
AND2_X1 U847 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U848 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
XNOR2_X1 U849 ( .A(n1173), .B(n1174), .ZN(n1172) );
XOR2_X1 U850 ( .A(KEYINPUT24), .B(n1175), .Z(n1174) );
NAND2_X1 U851 ( .A1(KEYINPUT38), .A2(n1176), .ZN(n1173) );
XNOR2_X1 U852 ( .A(n1177), .B(n1178), .ZN(n1176) );
NOR2_X1 U853 ( .A1(G125), .A2(KEYINPUT10), .ZN(n1178) );
NOR2_X1 U854 ( .A1(n1021), .A2(G952), .ZN(n1093) );
NAND2_X1 U855 ( .A1(n1179), .A2(n1180), .ZN(G48) );
NAND2_X1 U856 ( .A1(G146), .A2(n1181), .ZN(n1180) );
XOR2_X1 U857 ( .A(n1182), .B(KEYINPUT27), .Z(n1179) );
NAND2_X1 U858 ( .A1(n1138), .A2(n1183), .ZN(n1182) );
INV_X1 U859 ( .A(n1181), .ZN(n1138) );
NAND3_X1 U860 ( .A1(n1145), .A2(n1165), .A3(n1184), .ZN(n1181) );
XNOR2_X1 U861 ( .A(G143), .B(n1134), .ZN(G45) );
NAND4_X1 U862 ( .A1(n1184), .A2(n1050), .A3(n1185), .A4(n1186), .ZN(n1134) );
XNOR2_X1 U863 ( .A(G140), .B(n1187), .ZN(G42) );
NAND4_X1 U864 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1165), .ZN(n1187) );
XNOR2_X1 U865 ( .A(n1191), .B(KEYINPUT55), .ZN(n1188) );
XNOR2_X1 U866 ( .A(G137), .B(n1192), .ZN(G39) );
NAND4_X1 U867 ( .A1(n1189), .A2(n1145), .A3(n1044), .A4(n1193), .ZN(n1192) );
XNOR2_X1 U868 ( .A(KEYINPUT13), .B(n1152), .ZN(n1193) );
XOR2_X1 U869 ( .A(G134), .B(n1155), .Z(G36) );
AND3_X1 U870 ( .A1(n1050), .A2(n1151), .A3(n1194), .ZN(n1155) );
XNOR2_X1 U871 ( .A(n1081), .B(n1154), .ZN(G33) );
AND3_X1 U872 ( .A1(n1165), .A2(n1050), .A3(n1194), .ZN(n1154) );
INV_X1 U873 ( .A(n1148), .ZN(n1194) );
NAND2_X1 U874 ( .A1(n1189), .A2(n1152), .ZN(n1148) );
NOR2_X1 U875 ( .A1(n1052), .A2(n1046), .ZN(n1189) );
NAND2_X1 U876 ( .A1(n1022), .A2(n1195), .ZN(n1052) );
XOR2_X1 U877 ( .A(n1142), .B(n1196), .Z(G30) );
XNOR2_X1 U878 ( .A(KEYINPUT14), .B(n1197), .ZN(n1196) );
NAND3_X1 U879 ( .A1(n1145), .A2(n1151), .A3(n1184), .ZN(n1142) );
NOR3_X1 U880 ( .A1(n1016), .A2(n1191), .A3(n1046), .ZN(n1184) );
XOR2_X1 U881 ( .A(G101), .B(n1162), .Z(G3) );
AND3_X1 U882 ( .A1(n1044), .A2(n1163), .A3(n1198), .ZN(n1162) );
XOR2_X1 U883 ( .A(n1199), .B(G125), .Z(G27) );
NAND2_X1 U884 ( .A1(KEYINPUT59), .A2(n1135), .ZN(n1199) );
NAND3_X1 U885 ( .A1(n1190), .A2(n1040), .A3(n1200), .ZN(n1135) );
NOR3_X1 U886 ( .A1(n1042), .A2(n1191), .A3(n1016), .ZN(n1200) );
INV_X1 U887 ( .A(n1153), .ZN(n1016) );
INV_X1 U888 ( .A(n1152), .ZN(n1191) );
NAND2_X1 U889 ( .A1(n1051), .A2(n1201), .ZN(n1152) );
NAND4_X1 U890 ( .A1(G902), .A2(n1072), .A3(n1073), .A4(n1202), .ZN(n1201) );
XOR2_X1 U891 ( .A(KEYINPUT6), .B(G900), .Z(n1072) );
XNOR2_X1 U892 ( .A(G122), .B(n1156), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1040), .A2(n1164), .A3(n1185), .A4(n1186), .ZN(n1156) );
AND3_X1 U894 ( .A1(n1025), .A2(n1026), .A3(n1203), .ZN(n1164) );
XNOR2_X1 U895 ( .A(G119), .B(n1157), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1145), .A2(n1040), .A3(n1044), .A4(n1203), .ZN(n1157) );
NOR2_X1 U897 ( .A1(n1026), .A2(n1025), .ZN(n1145) );
INV_X1 U898 ( .A(n1204), .ZN(n1026) );
XOR2_X1 U899 ( .A(G116), .B(n1161), .Z(G18) );
AND3_X1 U900 ( .A1(n1198), .A2(n1151), .A3(n1040), .ZN(n1161) );
NOR2_X1 U901 ( .A1(n1186), .A2(n1205), .ZN(n1151) );
XNOR2_X1 U902 ( .A(G113), .B(n1206), .ZN(G15) );
NAND2_X1 U903 ( .A1(KEYINPUT53), .A2(n1160), .ZN(n1206) );
AND3_X1 U904 ( .A1(n1165), .A2(n1198), .A3(n1040), .ZN(n1160) );
NOR2_X1 U905 ( .A1(n1049), .A2(n1207), .ZN(n1040) );
INV_X1 U906 ( .A(n1048), .ZN(n1207) );
AND2_X1 U907 ( .A1(n1050), .A2(n1203), .ZN(n1198) );
NOR2_X1 U908 ( .A1(n1204), .A2(n1025), .ZN(n1050) );
INV_X1 U909 ( .A(n1042), .ZN(n1165) );
NAND2_X1 U910 ( .A1(n1205), .A2(n1186), .ZN(n1042) );
INV_X1 U911 ( .A(n1185), .ZN(n1205) );
XOR2_X1 U912 ( .A(G110), .B(n1208), .Z(G12) );
NOR2_X1 U913 ( .A1(KEYINPUT50), .A2(n1167), .ZN(n1208) );
NAND4_X1 U914 ( .A1(n1190), .A2(n1044), .A3(n1163), .A4(n1203), .ZN(n1167) );
AND2_X1 U915 ( .A1(n1153), .A2(n1209), .ZN(n1203) );
NAND2_X1 U916 ( .A1(n1051), .A2(n1210), .ZN(n1209) );
NAND4_X1 U917 ( .A1(G902), .A2(n1073), .A3(n1202), .A4(n1091), .ZN(n1210) );
INV_X1 U918 ( .A(G898), .ZN(n1091) );
XNOR2_X1 U919 ( .A(n1021), .B(KEYINPUT12), .ZN(n1073) );
NAND3_X1 U920 ( .A1(n1202), .A2(n1021), .A3(G952), .ZN(n1051) );
NAND2_X1 U921 ( .A1(G237), .A2(G234), .ZN(n1202) );
NOR2_X1 U922 ( .A1(n1022), .A2(n1024), .ZN(n1153) );
INV_X1 U923 ( .A(n1195), .ZN(n1024) );
NAND2_X1 U924 ( .A1(G214), .A2(n1211), .ZN(n1195) );
XOR2_X1 U925 ( .A(n1212), .B(n1213), .Z(n1022) );
AND2_X1 U926 ( .A1(n1211), .A2(G210), .ZN(n1213) );
NAND2_X1 U927 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
XNOR2_X1 U928 ( .A(G237), .B(KEYINPUT23), .ZN(n1214) );
NAND3_X1 U929 ( .A1(n1216), .A2(n1215), .A3(n1217), .ZN(n1212) );
XOR2_X1 U930 ( .A(KEYINPUT21), .B(n1218), .Z(n1217) );
NOR2_X1 U931 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U932 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
XNOR2_X1 U933 ( .A(n1116), .B(n1221), .ZN(n1220) );
XOR2_X1 U934 ( .A(G125), .B(n1175), .Z(n1221) );
AND2_X1 U935 ( .A1(G224), .A2(n1021), .ZN(n1175) );
INV_X1 U936 ( .A(n1171), .ZN(n1219) );
XNOR2_X1 U937 ( .A(n1089), .B(KEYINPUT57), .ZN(n1171) );
XOR2_X1 U938 ( .A(n1222), .B(n1223), .Z(n1089) );
XOR2_X1 U939 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U940 ( .A(G110), .B(G116), .ZN(n1225) );
NAND2_X1 U941 ( .A1(KEYINPUT0), .A2(n1226), .ZN(n1224) );
INV_X1 U942 ( .A(G119), .ZN(n1226) );
XNOR2_X1 U943 ( .A(n1227), .B(n1228), .ZN(n1222) );
XOR2_X1 U944 ( .A(n1229), .B(n1230), .Z(n1227) );
NAND2_X1 U945 ( .A1(KEYINPUT39), .A2(n1231), .ZN(n1229) );
INV_X1 U946 ( .A(n1046), .ZN(n1163) );
NAND2_X1 U947 ( .A1(n1049), .A2(n1048), .ZN(n1046) );
NAND2_X1 U948 ( .A1(G221), .A2(n1232), .ZN(n1048) );
NAND2_X1 U949 ( .A1(n1233), .A2(n1234), .ZN(n1049) );
NAND2_X1 U950 ( .A1(G469), .A2(n1060), .ZN(n1234) );
XOR2_X1 U951 ( .A(KEYINPUT15), .B(n1235), .Z(n1233) );
NOR2_X1 U952 ( .A1(G469), .A2(n1060), .ZN(n1235) );
NAND2_X1 U953 ( .A1(n1236), .A2(n1215), .ZN(n1060) );
XOR2_X1 U954 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U955 ( .A(n1239), .B(n1240), .ZN(n1238) );
NAND2_X1 U956 ( .A1(KEYINPUT30), .A2(n1241), .ZN(n1240) );
XOR2_X1 U957 ( .A(n1123), .B(n1076), .Z(n1241) );
XNOR2_X1 U958 ( .A(n1242), .B(G128), .ZN(n1076) );
NAND2_X1 U959 ( .A1(KEYINPUT36), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U960 ( .A(n1244), .B(n1245), .ZN(n1243) );
XNOR2_X1 U961 ( .A(KEYINPUT32), .B(n1183), .ZN(n1245) );
XOR2_X1 U962 ( .A(n1230), .B(n1246), .Z(n1123) );
XNOR2_X1 U963 ( .A(G104), .B(n1115), .ZN(n1246) );
XOR2_X1 U964 ( .A(G101), .B(n1247), .Z(n1230) );
XOR2_X1 U965 ( .A(KEYINPUT44), .B(G107), .Z(n1247) );
NAND2_X1 U966 ( .A1(n1248), .A2(KEYINPUT1), .ZN(n1239) );
XNOR2_X1 U967 ( .A(G110), .B(n1249), .ZN(n1248) );
XOR2_X1 U968 ( .A(KEYINPUT11), .B(G140), .Z(n1249) );
NAND2_X1 U969 ( .A1(G227), .A2(n1021), .ZN(n1237) );
NOR2_X1 U970 ( .A1(n1185), .A2(n1186), .ZN(n1044) );
XNOR2_X1 U971 ( .A(n1250), .B(G475), .ZN(n1186) );
NAND2_X1 U972 ( .A1(n1105), .A2(n1215), .ZN(n1250) );
XNOR2_X1 U973 ( .A(n1228), .B(n1251), .ZN(n1105) );
XNOR2_X1 U974 ( .A(n1231), .B(n1252), .ZN(n1251) );
NOR2_X1 U975 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U976 ( .A(n1255), .B(KEYINPUT47), .Z(n1254) );
NAND2_X1 U977 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NOR2_X1 U978 ( .A1(n1256), .A2(n1257), .ZN(n1253) );
NAND2_X1 U979 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
OR2_X1 U980 ( .A1(n1260), .A2(G146), .ZN(n1259) );
XOR2_X1 U981 ( .A(n1261), .B(KEYINPUT61), .Z(n1258) );
NAND2_X1 U982 ( .A1(G146), .A2(n1260), .ZN(n1261) );
AND2_X1 U983 ( .A1(n1262), .A2(n1263), .ZN(n1256) );
NAND2_X1 U984 ( .A1(n1264), .A2(n1081), .ZN(n1263) );
XOR2_X1 U985 ( .A(KEYINPUT60), .B(n1265), .Z(n1262) );
NOR2_X1 U986 ( .A1(n1264), .A2(n1081), .ZN(n1265) );
INV_X1 U987 ( .A(G131), .ZN(n1081) );
AND2_X1 U988 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND2_X1 U989 ( .A1(n1268), .A2(n1244), .ZN(n1267) );
NAND2_X1 U990 ( .A1(G214), .A2(n1269), .ZN(n1268) );
NAND3_X1 U991 ( .A1(G214), .A2(n1269), .A3(G143), .ZN(n1266) );
XOR2_X1 U992 ( .A(n1108), .B(G113), .Z(n1228) );
INV_X1 U993 ( .A(G104), .ZN(n1108) );
XOR2_X1 U994 ( .A(G478), .B(n1270), .Z(n1185) );
NOR2_X1 U995 ( .A1(G902), .A2(n1101), .ZN(n1270) );
XNOR2_X1 U996 ( .A(n1271), .B(n1272), .ZN(n1101) );
XOR2_X1 U997 ( .A(G107), .B(n1273), .Z(n1272) );
XNOR2_X1 U998 ( .A(n1231), .B(G116), .ZN(n1273) );
INV_X1 U999 ( .A(G122), .ZN(n1231) );
XOR2_X1 U1000 ( .A(n1274), .B(n1275), .Z(n1271) );
NOR2_X1 U1001 ( .A1(KEYINPUT34), .A2(n1276), .ZN(n1275) );
XOR2_X1 U1002 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U1003 ( .A(G134), .B(n1197), .ZN(n1278) );
XNOR2_X1 U1004 ( .A(KEYINPUT51), .B(n1244), .ZN(n1277) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1279), .ZN(n1274) );
INV_X1 U1006 ( .A(n1034), .ZN(n1190) );
NAND2_X1 U1007 ( .A1(n1025), .A2(n1204), .ZN(n1034) );
XOR2_X1 U1008 ( .A(n1280), .B(n1097), .Z(n1204) );
NAND2_X1 U1009 ( .A1(G217), .A2(n1232), .ZN(n1097) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1215), .ZN(n1232) );
NAND2_X1 U1011 ( .A1(n1215), .A2(n1095), .ZN(n1280) );
NAND2_X1 U1012 ( .A1(n1281), .A2(n1282), .ZN(n1095) );
NAND2_X1 U1013 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U1014 ( .A(KEYINPUT26), .B(n1285), .Z(n1281) );
NOR2_X1 U1015 ( .A1(n1283), .A2(n1284), .ZN(n1285) );
XNOR2_X1 U1016 ( .A(n1286), .B(n1287), .ZN(n1284) );
XNOR2_X1 U1017 ( .A(KEYINPUT25), .B(n1080), .ZN(n1287) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1279), .ZN(n1286) );
AND2_X1 U1019 ( .A1(G234), .A2(n1021), .ZN(n1279) );
INV_X1 U1020 ( .A(G953), .ZN(n1021) );
XOR2_X1 U1021 ( .A(n1288), .B(n1289), .Z(n1283) );
XNOR2_X1 U1022 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U1023 ( .A1(KEYINPUT52), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U1024 ( .A(G146), .B(n1260), .ZN(n1292) );
XNOR2_X1 U1025 ( .A(n1079), .B(KEYINPUT49), .ZN(n1260) );
XNOR2_X1 U1026 ( .A(G125), .B(G140), .ZN(n1079) );
NAND2_X1 U1027 ( .A1(n1293), .A2(KEYINPUT41), .ZN(n1290) );
XNOR2_X1 U1028 ( .A(G119), .B(n1294), .ZN(n1293) );
XNOR2_X1 U1029 ( .A(KEYINPUT7), .B(n1197), .ZN(n1294) );
XNOR2_X1 U1030 ( .A(G110), .B(KEYINPUT19), .ZN(n1288) );
XOR2_X1 U1031 ( .A(n1295), .B(G472), .Z(n1025) );
NAND3_X1 U1032 ( .A1(n1296), .A2(n1297), .A3(n1215), .ZN(n1295) );
INV_X1 U1033 ( .A(G902), .ZN(n1215) );
NAND2_X1 U1034 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1035 ( .A(KEYINPUT54), .B(n1300), .ZN(n1298) );
NAND2_X1 U1036 ( .A1(KEYINPUT29), .A2(n1117), .ZN(n1300) );
NAND3_X1 U1037 ( .A1(n1117), .A2(n1301), .A3(n1302), .ZN(n1296) );
INV_X1 U1038 ( .A(n1299), .ZN(n1302) );
NAND2_X1 U1039 ( .A1(n1303), .A2(n1304), .ZN(n1299) );
NAND2_X1 U1040 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U1041 ( .A(KEYINPUT5), .B(n1118), .Z(n1306) );
XNOR2_X1 U1042 ( .A(n1177), .B(n1307), .ZN(n1305) );
NAND2_X1 U1043 ( .A1(n1308), .A2(n1309), .ZN(n1303) );
XNOR2_X1 U1044 ( .A(n1116), .B(n1307), .ZN(n1309) );
NAND2_X1 U1045 ( .A1(KEYINPUT9), .A2(n1115), .ZN(n1307) );
NAND2_X1 U1046 ( .A1(n1310), .A2(n1311), .ZN(n1115) );
NAND2_X1 U1047 ( .A1(G131), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1048 ( .A(n1313), .B(KEYINPUT46), .Z(n1310) );
OR2_X1 U1049 ( .A1(n1312), .A2(G131), .ZN(n1313) );
XNOR2_X1 U1050 ( .A(G134), .B(n1080), .ZN(n1312) );
INV_X1 U1051 ( .A(G137), .ZN(n1080) );
INV_X1 U1052 ( .A(n1177), .ZN(n1116) );
NAND2_X1 U1053 ( .A1(n1314), .A2(n1315), .ZN(n1177) );
NAND2_X1 U1054 ( .A1(n1316), .A2(n1197), .ZN(n1315) );
XOR2_X1 U1055 ( .A(n1317), .B(KEYINPUT58), .Z(n1314) );
OR2_X1 U1056 ( .A1(n1316), .A2(n1197), .ZN(n1317) );
INV_X1 U1057 ( .A(G128), .ZN(n1197) );
XOR2_X1 U1058 ( .A(n1318), .B(n1244), .Z(n1316) );
INV_X1 U1059 ( .A(G143), .ZN(n1244) );
NAND2_X1 U1060 ( .A1(KEYINPUT43), .A2(n1183), .ZN(n1318) );
INV_X1 U1061 ( .A(G146), .ZN(n1183) );
XNOR2_X1 U1062 ( .A(n1118), .B(KEYINPUT33), .ZN(n1308) );
XNOR2_X1 U1063 ( .A(n1319), .B(n1320), .ZN(n1118) );
NOR2_X1 U1064 ( .A1(KEYINPUT2), .A2(G113), .ZN(n1320) );
XNOR2_X1 U1065 ( .A(G116), .B(G119), .ZN(n1319) );
XNOR2_X1 U1066 ( .A(KEYINPUT29), .B(KEYINPUT54), .ZN(n1301) );
XNOR2_X1 U1067 ( .A(n1321), .B(G101), .ZN(n1117) );
NAND2_X1 U1068 ( .A1(G210), .A2(n1269), .ZN(n1321) );
NOR2_X1 U1069 ( .A1(G953), .A2(G237), .ZN(n1269) );
endmodule


