//Key = 0011110101111101100011011000100010101001110010000001000111110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359;

XOR2_X1 U755 ( .A(n1041), .B(n1042), .Z(G9) );
XNOR2_X1 U756 ( .A(KEYINPUT41), .B(n1043), .ZN(n1042) );
NAND4_X1 U757 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1041) );
XOR2_X1 U758 ( .A(n1048), .B(KEYINPUT61), .Z(n1044) );
NOR2_X1 U759 ( .A1(n1049), .A2(n1050), .ZN(G75) );
NOR4_X1 U760 ( .A1(G953), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1050) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR3_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1061) );
NOR2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR3_X1 U769 ( .A1(n1064), .A2(n1072), .A3(n1065), .ZN(n1056) );
NOR2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR3_X1 U771 ( .A1(n1058), .A2(n1075), .A3(n1076), .ZN(n1074) );
AND2_X1 U772 ( .A1(n1077), .A2(n1070), .ZN(n1076) );
NOR3_X1 U773 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1070) );
NOR2_X1 U774 ( .A1(n1045), .A2(n1077), .ZN(n1075) );
NOR3_X1 U775 ( .A1(n1060), .A2(n1066), .A3(n1081), .ZN(n1073) );
NOR2_X1 U776 ( .A1(n1046), .A2(n1082), .ZN(n1081) );
XNOR2_X1 U777 ( .A(n1083), .B(KEYINPUT24), .ZN(n1082) );
NOR3_X1 U778 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1049) );
AND4_X1 U779 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1051) );
NOR4_X1 U780 ( .A1(n1066), .A2(n1088), .A3(n1078), .A4(n1089), .ZN(n1087) );
NOR3_X1 U781 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR3_X1 U783 ( .A1(G469), .A2(KEYINPUT46), .A3(n1095), .ZN(n1091) );
INV_X1 U784 ( .A(n1093), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1096), .A2(KEYINPUT49), .ZN(n1093) );
AND2_X1 U786 ( .A1(n1096), .A2(KEYINPUT46), .ZN(n1090) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1088) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U789 ( .A(KEYINPUT30), .B(n1101), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1086) );
XNOR2_X1 U791 ( .A(KEYINPUT31), .B(n1104), .ZN(n1103) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1102) );
XNOR2_X1 U793 ( .A(KEYINPUT43), .B(n1107), .ZN(n1106) );
NOR3_X1 U794 ( .A1(n1108), .A2(KEYINPUT22), .A3(G902), .ZN(n1105) );
XNOR2_X1 U795 ( .A(KEYINPUT55), .B(n1109), .ZN(n1085) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1116), .B(KEYINPUT0), .Z(n1114) );
NAND3_X1 U800 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
XOR2_X1 U801 ( .A(KEYINPUT62), .B(n1120), .Z(n1118) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1112) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U804 ( .A(n1125), .B(n1126), .Z(n1121) );
XOR2_X1 U805 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U806 ( .A(G131), .B(n1129), .ZN(n1127) );
XNOR2_X1 U807 ( .A(G134), .B(n1130), .ZN(n1125) );
XNOR2_X1 U808 ( .A(G140), .B(n1131), .ZN(n1130) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1115), .ZN(n1110) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1124), .ZN(n1132) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(G69) );
NAND2_X1 U812 ( .A1(G953), .A2(n1136), .ZN(n1135) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1136) );
NAND2_X1 U814 ( .A1(KEYINPUT23), .A2(n1137), .ZN(n1134) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
XNOR2_X1 U818 ( .A(G953), .B(KEYINPUT16), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR3_X1 U822 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
XNOR2_X1 U823 ( .A(KEYINPUT44), .B(n1153), .ZN(n1150) );
NAND2_X1 U824 ( .A1(KEYINPUT40), .A2(n1154), .ZN(n1148) );
NOR2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(G63) );
XOR2_X1 U826 ( .A(KEYINPUT42), .B(n1146), .Z(n1156) );
XNOR2_X1 U827 ( .A(n1157), .B(n1158), .ZN(n1155) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1152), .ZN(n1158) );
NOR2_X1 U829 ( .A1(n1146), .A2(n1160), .ZN(G60) );
XOR2_X1 U830 ( .A(n1161), .B(n1108), .Z(n1160) );
NOR2_X1 U831 ( .A1(n1107), .A2(n1152), .ZN(n1161) );
INV_X1 U832 ( .A(G475), .ZN(n1107) );
XNOR2_X1 U833 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1164), .ZN(G57) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U836 ( .A(n1167), .B(n1168), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1165) );
XOR2_X1 U839 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U840 ( .A1(n1175), .A2(n1152), .ZN(n1174) );
NAND2_X1 U841 ( .A1(n1176), .A2(KEYINPUT39), .ZN(n1171) );
XNOR2_X1 U842 ( .A(G101), .B(KEYINPUT3), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(n1163) );
XOR2_X1 U844 ( .A(KEYINPUT8), .B(G952), .Z(n1178) );
XNOR2_X1 U845 ( .A(G953), .B(KEYINPUT37), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1146), .A2(n1179), .ZN(G54) );
XOR2_X1 U847 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U848 ( .A(n1182), .B(n1183), .Z(n1180) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1182) );
NOR2_X1 U850 ( .A1(n1094), .A2(n1152), .ZN(n1185) );
NAND2_X1 U851 ( .A1(KEYINPUT2), .A2(n1186), .ZN(n1184) );
NOR2_X1 U852 ( .A1(n1146), .A2(n1187), .ZN(G51) );
NOR2_X1 U853 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U854 ( .A(n1190), .B(KEYINPUT32), .Z(n1189) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
OR2_X1 U856 ( .A1(n1152), .A2(n1101), .ZN(n1192) );
XOR2_X1 U857 ( .A(KEYINPUT38), .B(n1193), .Z(n1191) );
NOR3_X1 U858 ( .A1(n1193), .A2(n1101), .A3(n1152), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1194), .A2(n1053), .ZN(n1152) );
NAND4_X1 U860 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1119), .ZN(n1053) );
AND3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1119) );
NOR2_X1 U862 ( .A1(n1120), .A2(n1201), .ZN(n1197) );
XOR2_X1 U863 ( .A(n1144), .B(KEYINPUT26), .Z(n1201) );
NAND4_X1 U864 ( .A1(n1202), .A2(n1162), .A3(n1203), .A4(n1204), .ZN(n1144) );
NAND3_X1 U865 ( .A1(n1083), .A2(n1045), .A3(n1205), .ZN(n1162) );
NAND3_X1 U866 ( .A1(n1045), .A2(n1046), .A3(n1205), .ZN(n1202) );
INV_X1 U867 ( .A(n1145), .ZN(n1196) );
NAND4_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1145) );
NAND3_X1 U869 ( .A1(n1210), .A2(n1083), .A3(n1080), .ZN(n1206) );
XNOR2_X1 U870 ( .A(n1117), .B(KEYINPUT15), .ZN(n1195) );
AND4_X1 U871 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1117) );
NAND3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1211) );
XNOR2_X1 U873 ( .A(KEYINPUT45), .B(n1218), .ZN(n1194) );
XOR2_X1 U874 ( .A(n1219), .B(n1220), .Z(n1193) );
XNOR2_X1 U875 ( .A(n1141), .B(KEYINPUT52), .ZN(n1219) );
AND2_X1 U876 ( .A1(n1221), .A2(G953), .ZN(n1146) );
XNOR2_X1 U877 ( .A(KEYINPUT8), .B(G952), .ZN(n1221) );
XNOR2_X1 U878 ( .A(G146), .B(n1212), .ZN(G48) );
NAND4_X1 U879 ( .A1(n1215), .A2(n1083), .A3(n1047), .A4(n1222), .ZN(n1212) );
XNOR2_X1 U880 ( .A(n1223), .B(n1224), .ZN(G45) );
NAND2_X1 U881 ( .A1(KEYINPUT56), .A2(n1213), .ZN(n1223) );
NAND4_X1 U882 ( .A1(n1225), .A2(n1222), .A3(n1047), .A4(n1226), .ZN(n1213) );
NOR2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
INV_X1 U884 ( .A(n1080), .ZN(n1227) );
XNOR2_X1 U885 ( .A(G140), .B(n1214), .ZN(G42) );
NAND3_X1 U886 ( .A1(n1079), .A2(n1083), .A3(n1217), .ZN(n1214) );
XNOR2_X1 U887 ( .A(G137), .B(n1229), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1215), .A2(n1230), .A3(n1217), .ZN(n1229) );
XNOR2_X1 U889 ( .A(KEYINPUT33), .B(n1058), .ZN(n1230) );
XNOR2_X1 U890 ( .A(G134), .B(n1200), .ZN(G36) );
NAND3_X1 U891 ( .A1(n1080), .A2(n1046), .A3(n1217), .ZN(n1200) );
XNOR2_X1 U892 ( .A(G131), .B(n1198), .ZN(G33) );
NAND3_X1 U893 ( .A1(n1080), .A2(n1083), .A3(n1217), .ZN(n1198) );
NOR3_X1 U894 ( .A1(n1063), .A2(n1231), .A3(n1064), .ZN(n1217) );
OR2_X1 U895 ( .A1(n1071), .A2(n1078), .ZN(n1064) );
INV_X1 U896 ( .A(n1232), .ZN(n1071) );
XNOR2_X1 U897 ( .A(G128), .B(n1199), .ZN(G30) );
NAND4_X1 U898 ( .A1(n1215), .A2(n1046), .A3(n1047), .A4(n1222), .ZN(n1199) );
XOR2_X1 U899 ( .A(n1203), .B(n1233), .Z(G3) );
XNOR2_X1 U900 ( .A(G101), .B(KEYINPUT50), .ZN(n1233) );
NAND3_X1 U901 ( .A1(n1216), .A2(n1080), .A3(n1205), .ZN(n1203) );
XOR2_X1 U902 ( .A(G125), .B(n1120), .Z(G27) );
AND4_X1 U903 ( .A1(n1234), .A2(n1083), .A3(n1079), .A4(n1235), .ZN(n1120) );
NOR3_X1 U904 ( .A1(n1236), .A2(n1066), .A3(n1231), .ZN(n1235) );
INV_X1 U905 ( .A(n1222), .ZN(n1231) );
NAND2_X1 U906 ( .A1(n1237), .A2(n1055), .ZN(n1222) );
NAND4_X1 U907 ( .A1(n1123), .A2(G902), .A3(n1238), .A4(n1124), .ZN(n1237) );
INV_X1 U908 ( .A(G900), .ZN(n1124) );
INV_X1 U909 ( .A(n1239), .ZN(n1123) );
XNOR2_X1 U910 ( .A(G122), .B(n1207), .ZN(G24) );
OR4_X1 U911 ( .A1(n1228), .A2(n1240), .A3(n1060), .A4(n1084), .ZN(n1207) );
INV_X1 U912 ( .A(n1045), .ZN(n1060) );
NOR2_X1 U913 ( .A1(n1241), .A2(n1242), .ZN(n1045) );
XNOR2_X1 U914 ( .A(G119), .B(n1208), .ZN(G21) );
NAND3_X1 U915 ( .A1(n1216), .A2(n1210), .A3(n1215), .ZN(n1208) );
NOR2_X1 U916 ( .A1(n1104), .A2(n1109), .ZN(n1215) );
XNOR2_X1 U917 ( .A(G116), .B(n1209), .ZN(G18) );
NAND3_X1 U918 ( .A1(n1210), .A2(n1046), .A3(n1080), .ZN(n1209) );
AND2_X1 U919 ( .A1(n1243), .A2(n1225), .ZN(n1046) );
INV_X1 U920 ( .A(n1240), .ZN(n1210) );
XOR2_X1 U921 ( .A(n1244), .B(n1245), .Z(G15) );
NOR2_X1 U922 ( .A1(KEYINPUT54), .A2(n1246), .ZN(n1245) );
INV_X1 U923 ( .A(G113), .ZN(n1246) );
NOR3_X1 U924 ( .A1(n1240), .A2(n1247), .A3(n1248), .ZN(n1244) );
INV_X1 U925 ( .A(n1083), .ZN(n1248) );
NOR2_X1 U926 ( .A1(n1228), .A2(n1225), .ZN(n1083) );
XNOR2_X1 U927 ( .A(n1243), .B(KEYINPUT57), .ZN(n1228) );
XNOR2_X1 U928 ( .A(n1080), .B(KEYINPUT1), .ZN(n1247) );
NOR2_X1 U929 ( .A1(n1242), .A2(n1109), .ZN(n1080) );
INV_X1 U930 ( .A(n1241), .ZN(n1109) );
NAND4_X1 U931 ( .A1(n1234), .A2(n1069), .A3(n1048), .A4(n1077), .ZN(n1240) );
INV_X1 U932 ( .A(n1065), .ZN(n1234) );
XNOR2_X1 U933 ( .A(G110), .B(n1204), .ZN(G12) );
NAND3_X1 U934 ( .A1(n1216), .A2(n1079), .A3(n1205), .ZN(n1204) );
AND2_X1 U935 ( .A1(n1047), .A2(n1048), .ZN(n1205) );
NAND2_X1 U936 ( .A1(n1055), .A2(n1249), .ZN(n1048) );
NAND3_X1 U937 ( .A1(n1140), .A2(n1238), .A3(G902), .ZN(n1249) );
NOR2_X1 U938 ( .A1(n1239), .A2(G898), .ZN(n1140) );
XOR2_X1 U939 ( .A(G953), .B(KEYINPUT34), .Z(n1239) );
NAND3_X1 U940 ( .A1(n1238), .A2(n1115), .A3(G952), .ZN(n1055) );
INV_X1 U941 ( .A(G953), .ZN(n1115) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1238) );
NOR2_X1 U943 ( .A1(n1236), .A2(n1063), .ZN(n1047) );
NAND2_X1 U944 ( .A1(n1065), .A2(n1077), .ZN(n1063) );
INV_X1 U945 ( .A(n1066), .ZN(n1077) );
NOR2_X1 U946 ( .A1(n1250), .A2(n1151), .ZN(n1066) );
XOR2_X1 U947 ( .A(n1096), .B(n1251), .Z(n1065) );
NOR2_X1 U948 ( .A1(KEYINPUT17), .A2(n1094), .ZN(n1251) );
INV_X1 U949 ( .A(G469), .ZN(n1094) );
AND2_X1 U950 ( .A1(n1252), .A2(n1218), .ZN(n1096) );
XOR2_X1 U951 ( .A(n1253), .B(n1181), .Z(n1252) );
XNOR2_X1 U952 ( .A(n1254), .B(n1167), .ZN(n1181) );
XNOR2_X1 U953 ( .A(G110), .B(G140), .ZN(n1254) );
XNOR2_X1 U954 ( .A(n1255), .B(n1186), .ZN(n1253) );
NOR2_X1 U955 ( .A1(n1133), .A2(n1256), .ZN(n1186) );
INV_X1 U956 ( .A(G227), .ZN(n1133) );
NAND2_X1 U957 ( .A1(KEYINPUT13), .A2(n1183), .ZN(n1255) );
XNOR2_X1 U958 ( .A(n1257), .B(n1258), .ZN(n1183) );
XOR2_X1 U959 ( .A(G104), .B(n1259), .Z(n1258) );
XNOR2_X1 U960 ( .A(KEYINPUT25), .B(n1043), .ZN(n1259) );
XOR2_X1 U961 ( .A(n1260), .B(n1129), .Z(n1257) );
XNOR2_X1 U962 ( .A(n1261), .B(KEYINPUT6), .ZN(n1129) );
NAND2_X1 U963 ( .A1(KEYINPUT5), .A2(n1224), .ZN(n1261) );
XNOR2_X1 U964 ( .A(G101), .B(n1262), .ZN(n1260) );
INV_X1 U965 ( .A(n1069), .ZN(n1236) );
NOR2_X1 U966 ( .A1(n1232), .A2(n1078), .ZN(n1069) );
AND2_X1 U967 ( .A1(G214), .A2(n1263), .ZN(n1078) );
NAND2_X1 U968 ( .A1(n1264), .A2(n1265), .ZN(n1232) );
NAND2_X1 U969 ( .A1(KEYINPUT4), .A2(n1266), .ZN(n1265) );
NAND2_X1 U970 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U971 ( .A1(n1101), .A2(n1269), .ZN(n1268) );
INV_X1 U972 ( .A(n1097), .ZN(n1267) );
NOR2_X1 U973 ( .A1(n1101), .A2(n1269), .ZN(n1097) );
NAND2_X1 U974 ( .A1(n1270), .A2(n1271), .ZN(n1264) );
INV_X1 U975 ( .A(KEYINPUT4), .ZN(n1271) );
XNOR2_X1 U976 ( .A(n1099), .B(n1101), .ZN(n1270) );
NAND2_X1 U977 ( .A1(G210), .A2(n1263), .ZN(n1101) );
NAND2_X1 U978 ( .A1(n1272), .A2(n1218), .ZN(n1263) );
INV_X1 U979 ( .A(n1269), .ZN(n1099) );
NAND2_X1 U980 ( .A1(n1273), .A2(n1218), .ZN(n1269) );
XNOR2_X1 U981 ( .A(n1274), .B(n1275), .ZN(n1273) );
INV_X1 U982 ( .A(n1141), .ZN(n1275) );
XNOR2_X1 U983 ( .A(n1276), .B(n1277), .ZN(n1141) );
XOR2_X1 U984 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U985 ( .A(n1280), .B(n1043), .ZN(n1279) );
NAND2_X1 U986 ( .A1(KEYINPUT51), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U987 ( .A(G110), .B(KEYINPUT48), .ZN(n1278) );
XNOR2_X1 U988 ( .A(n1170), .B(n1282), .ZN(n1276) );
XNOR2_X1 U989 ( .A(n1283), .B(n1284), .ZN(n1282) );
NOR2_X1 U990 ( .A1(G101), .A2(KEYINPUT63), .ZN(n1284) );
NAND2_X1 U991 ( .A1(KEYINPUT59), .A2(G104), .ZN(n1283) );
NAND2_X1 U992 ( .A1(KEYINPUT36), .A2(n1220), .ZN(n1274) );
XOR2_X1 U993 ( .A(n1285), .B(n1128), .Z(n1220) );
XOR2_X1 U994 ( .A(G125), .B(n1262), .Z(n1128) );
XNOR2_X1 U995 ( .A(G143), .B(n1286), .ZN(n1285) );
AND2_X1 U996 ( .A1(n1287), .A2(G224), .ZN(n1286) );
NOR2_X1 U997 ( .A1(n1241), .A2(n1104), .ZN(n1079) );
INV_X1 U998 ( .A(n1242), .ZN(n1104) );
XNOR2_X1 U999 ( .A(n1288), .B(n1289), .ZN(n1242) );
NOR2_X1 U1000 ( .A1(n1151), .A2(n1153), .ZN(n1289) );
NOR2_X1 U1001 ( .A1(n1290), .A2(G902), .ZN(n1151) );
NAND2_X1 U1002 ( .A1(n1154), .A2(n1218), .ZN(n1288) );
XNOR2_X1 U1003 ( .A(n1291), .B(n1292), .ZN(n1154) );
NOR2_X1 U1004 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NOR2_X1 U1005 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U1006 ( .A(KEYINPUT18), .B(n1131), .ZN(n1296) );
AND2_X1 U1007 ( .A1(G137), .A2(n1295), .ZN(n1293) );
NOR3_X1 U1008 ( .A1(n1256), .A2(n1250), .A3(n1290), .ZN(n1295) );
INV_X1 U1009 ( .A(G221), .ZN(n1250) );
NAND3_X1 U1010 ( .A1(n1297), .A2(n1298), .A3(KEYINPUT20), .ZN(n1291) );
NAND3_X1 U1011 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1298) );
INV_X1 U1012 ( .A(KEYINPUT11), .ZN(n1301) );
NAND2_X1 U1013 ( .A1(n1302), .A2(KEYINPUT11), .ZN(n1297) );
XOR2_X1 U1014 ( .A(n1300), .B(n1299), .Z(n1302) );
XNOR2_X1 U1015 ( .A(n1303), .B(n1304), .ZN(n1299) );
XOR2_X1 U1016 ( .A(G119), .B(G110), .Z(n1304) );
NAND2_X1 U1017 ( .A1(KEYINPUT28), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1018 ( .A(n1306), .B(n1307), .Z(n1300) );
NAND2_X1 U1019 ( .A1(KEYINPUT7), .A2(G146), .ZN(n1306) );
XOR2_X1 U1020 ( .A(n1308), .B(n1175), .Z(n1241) );
INV_X1 U1021 ( .A(G472), .ZN(n1175) );
NAND2_X1 U1022 ( .A1(n1309), .A2(n1218), .ZN(n1308) );
XNOR2_X1 U1023 ( .A(n1173), .B(n1310), .ZN(n1309) );
XOR2_X1 U1024 ( .A(G101), .B(n1311), .Z(n1310) );
NOR2_X1 U1025 ( .A1(KEYINPUT47), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1026 ( .A(n1313), .B(n1170), .ZN(n1312) );
XOR2_X1 U1027 ( .A(G113), .B(n1314), .Z(n1170) );
XOR2_X1 U1028 ( .A(G119), .B(G116), .Z(n1314) );
NAND2_X1 U1029 ( .A1(n1315), .A2(KEYINPUT9), .ZN(n1313) );
XOR2_X1 U1030 ( .A(n1169), .B(n1316), .Z(n1315) );
NOR2_X1 U1031 ( .A1(KEYINPUT35), .A2(n1167), .ZN(n1316) );
AND2_X1 U1032 ( .A1(n1317), .A2(n1318), .ZN(n1167) );
NAND2_X1 U1033 ( .A1(G137), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1034 ( .A1(n1320), .A2(n1131), .ZN(n1317) );
INV_X1 U1035 ( .A(G137), .ZN(n1131) );
XNOR2_X1 U1036 ( .A(KEYINPUT14), .B(n1319), .ZN(n1320) );
XOR2_X1 U1037 ( .A(n1321), .B(n1322), .Z(n1319) );
XOR2_X1 U1038 ( .A(KEYINPUT27), .B(G134), .Z(n1322) );
XNOR2_X1 U1039 ( .A(G143), .B(n1262), .ZN(n1169) );
XNOR2_X1 U1040 ( .A(n1305), .B(G146), .ZN(n1262) );
NAND3_X1 U1041 ( .A1(n1287), .A2(n1272), .A3(G210), .ZN(n1173) );
INV_X1 U1042 ( .A(G237), .ZN(n1272) );
INV_X1 U1043 ( .A(n1256), .ZN(n1287) );
INV_X1 U1044 ( .A(n1058), .ZN(n1216) );
NAND2_X1 U1045 ( .A1(n1084), .A2(n1243), .ZN(n1058) );
XNOR2_X1 U1046 ( .A(G475), .B(n1323), .ZN(n1243) );
NOR2_X1 U1047 ( .A1(G902), .A2(n1108), .ZN(n1323) );
XNOR2_X1 U1048 ( .A(n1324), .B(n1325), .ZN(n1108) );
XOR2_X1 U1049 ( .A(G104), .B(n1326), .Z(n1325) );
NOR3_X1 U1050 ( .A1(KEYINPUT53), .A2(n1327), .A3(n1328), .ZN(n1326) );
NOR2_X1 U1051 ( .A1(n1321), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1052 ( .A(n1330), .B(n1331), .ZN(n1329) );
NAND2_X1 U1053 ( .A1(KEYINPUT58), .A2(n1332), .ZN(n1330) );
INV_X1 U1054 ( .A(G131), .ZN(n1321) );
NOR2_X1 U1055 ( .A1(G131), .A2(n1333), .ZN(n1327) );
XOR2_X1 U1056 ( .A(n1331), .B(n1334), .Z(n1333) );
NOR2_X1 U1057 ( .A1(n1332), .A2(n1335), .ZN(n1334) );
INV_X1 U1058 ( .A(KEYINPUT58), .ZN(n1335) );
NOR2_X1 U1059 ( .A1(KEYINPUT19), .A2(n1336), .ZN(n1332) );
XNOR2_X1 U1060 ( .A(n1224), .B(n1337), .ZN(n1336) );
NOR3_X1 U1061 ( .A1(n1338), .A2(G237), .A3(n1256), .ZN(n1337) );
XOR2_X1 U1062 ( .A(KEYINPUT21), .B(G214), .Z(n1338) );
NAND2_X1 U1063 ( .A1(n1339), .A2(n1340), .ZN(n1331) );
NAND2_X1 U1064 ( .A1(n1307), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1065 ( .A(KEYINPUT12), .B(n1342), .Z(n1339) );
NOR2_X1 U1066 ( .A1(n1307), .A2(n1341), .ZN(n1342) );
INV_X1 U1067 ( .A(G146), .ZN(n1341) );
XNOR2_X1 U1068 ( .A(G125), .B(G140), .ZN(n1307) );
XNOR2_X1 U1069 ( .A(G113), .B(G122), .ZN(n1324) );
INV_X1 U1070 ( .A(n1225), .ZN(n1084) );
XOR2_X1 U1071 ( .A(n1343), .B(n1159), .Z(n1225) );
INV_X1 U1072 ( .A(G478), .ZN(n1159) );
NAND2_X1 U1073 ( .A1(n1157), .A2(n1218), .ZN(n1343) );
INV_X1 U1074 ( .A(G902), .ZN(n1218) );
XNOR2_X1 U1075 ( .A(n1344), .B(n1345), .ZN(n1157) );
XNOR2_X1 U1076 ( .A(n1305), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1077 ( .A(n1224), .B(G134), .ZN(n1346) );
INV_X1 U1078 ( .A(G143), .ZN(n1224) );
INV_X1 U1079 ( .A(G128), .ZN(n1305) );
XOR2_X1 U1080 ( .A(n1347), .B(n1348), .Z(n1344) );
NOR3_X1 U1081 ( .A1(n1153), .A2(n1290), .A3(n1256), .ZN(n1348) );
XOR2_X1 U1082 ( .A(G953), .B(KEYINPUT60), .Z(n1256) );
INV_X1 U1083 ( .A(G234), .ZN(n1290) );
INV_X1 U1084 ( .A(G217), .ZN(n1153) );
NAND3_X1 U1085 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1347) );
NAND2_X1 U1086 ( .A1(G107), .A2(n1352), .ZN(n1351) );
NAND2_X1 U1087 ( .A1(KEYINPUT29), .A2(n1353), .ZN(n1350) );
NAND2_X1 U1088 ( .A1(n1354), .A2(n1043), .ZN(n1353) );
INV_X1 U1089 ( .A(G107), .ZN(n1043) );
XNOR2_X1 U1090 ( .A(n1355), .B(n1352), .ZN(n1354) );
NAND2_X1 U1091 ( .A1(n1356), .A2(n1357), .ZN(n1349) );
INV_X1 U1092 ( .A(KEYINPUT29), .ZN(n1357) );
NAND2_X1 U1093 ( .A1(n1358), .A2(n1359), .ZN(n1356) );
NAND2_X1 U1094 ( .A1(n1352), .A2(n1355), .ZN(n1359) );
OR3_X1 U1095 ( .A1(n1352), .A2(G107), .A3(n1355), .ZN(n1358) );
INV_X1 U1096 ( .A(KEYINPUT10), .ZN(n1355) );
XNOR2_X1 U1097 ( .A(G116), .B(n1281), .ZN(n1352) );
INV_X1 U1098 ( .A(G122), .ZN(n1281) );
endmodule


