//Key = 0001100011011011010010010000101000000110111111110010001001010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275;

XOR2_X1 U705 ( .A(G107), .B(n977), .Z(G9) );
NAND3_X1 U706 ( .A1(n978), .A2(n979), .A3(n980), .ZN(G75) );
NAND2_X1 U707 ( .A1(G952), .A2(n981), .ZN(n980) );
NAND4_X1 U708 ( .A1(n982), .A2(n983), .A3(n984), .A4(n985), .ZN(n981) );
NAND2_X1 U709 ( .A1(n986), .A2(n987), .ZN(n985) );
NAND2_X1 U710 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND4_X1 U711 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n989) );
NAND2_X1 U712 ( .A1(n994), .A2(n995), .ZN(n988) );
NAND2_X1 U713 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND3_X1 U714 ( .A1(n998), .A2(n999), .A3(n992), .ZN(n997) );
NAND2_X1 U715 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U716 ( .A1(n990), .A2(n1002), .ZN(n1000) );
NAND2_X1 U717 ( .A1(n1003), .A2(n1004), .ZN(n998) );
NAND2_X1 U718 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
XOR2_X1 U719 ( .A(n1007), .B(KEYINPUT45), .Z(n1005) );
NAND2_X1 U720 ( .A1(n991), .A2(n1008), .ZN(n996) );
NAND2_X1 U721 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U722 ( .A1(n992), .A2(n1011), .ZN(n1010) );
NAND2_X1 U723 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U724 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
INV_X1 U725 ( .A(n1016), .ZN(n1012) );
NAND2_X1 U726 ( .A1(n990), .A2(n1017), .ZN(n1009) );
NAND2_X1 U727 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
INV_X1 U728 ( .A(n1020), .ZN(n1019) );
XOR2_X1 U729 ( .A(KEYINPUT41), .B(n1021), .Z(n1018) );
INV_X1 U730 ( .A(n1022), .ZN(n986) );
NAND2_X1 U731 ( .A1(KEYINPUT19), .A2(n1023), .ZN(n984) );
XOR2_X1 U732 ( .A(n1024), .B(KEYINPUT0), .Z(n982) );
NAND4_X1 U733 ( .A1(n991), .A2(n992), .A3(n1025), .A4(n1026), .ZN(n1024) );
NOR2_X1 U734 ( .A1(n1007), .A2(n1022), .ZN(n1026) );
NAND2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n978) );
NAND2_X1 U736 ( .A1(KEYINPUT19), .A2(G952), .ZN(n1028) );
INV_X1 U737 ( .A(n1023), .ZN(n1027) );
NAND4_X1 U738 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1023) );
NOR4_X1 U739 ( .A1(n1014), .A2(n1003), .A3(n1033), .A4(n1034), .ZN(n1032) );
XOR2_X1 U740 ( .A(KEYINPUT17), .B(n1035), .Z(n1034) );
NOR2_X1 U741 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR3_X1 U742 ( .A1(n1038), .A2(KEYINPUT60), .A3(n1039), .ZN(n1037) );
INV_X1 U743 ( .A(G478), .ZN(n1038) );
NOR2_X1 U744 ( .A1(G478), .A2(n1040), .ZN(n1036) );
NOR2_X1 U745 ( .A1(KEYINPUT60), .A2(n1039), .ZN(n1040) );
XNOR2_X1 U746 ( .A(n1041), .B(n1042), .ZN(n1033) );
NOR2_X1 U747 ( .A1(G475), .A2(KEYINPUT13), .ZN(n1042) );
INV_X1 U748 ( .A(n1001), .ZN(n1003) );
NOR2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1031) );
XOR2_X1 U750 ( .A(n1045), .B(n1046), .Z(n1044) );
NAND2_X1 U751 ( .A1(KEYINPUT50), .A2(n1047), .ZN(n1046) );
XOR2_X1 U752 ( .A(n1048), .B(G469), .Z(n1030) );
XOR2_X1 U753 ( .A(n1049), .B(n1050), .Z(n1029) );
XOR2_X1 U754 ( .A(n1051), .B(n1052), .Z(G72) );
NOR2_X1 U755 ( .A1(n1053), .A2(n979), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1051) );
NAND2_X1 U758 ( .A1(n1058), .A2(n979), .ZN(n1057) );
XOR2_X1 U759 ( .A(n1059), .B(n1060), .Z(n1058) );
NAND3_X1 U760 ( .A1(G900), .A2(n1060), .A3(G953), .ZN(n1056) );
XNOR2_X1 U761 ( .A(n1061), .B(n1062), .ZN(n1060) );
XOR2_X1 U762 ( .A(G125), .B(n1063), .Z(n1062) );
XOR2_X1 U763 ( .A(G140), .B(G131), .Z(n1063) );
XOR2_X1 U764 ( .A(n1064), .B(n1065), .Z(n1061) );
NAND2_X1 U765 ( .A1(KEYINPUT54), .A2(n1066), .ZN(n1064) );
XOR2_X1 U766 ( .A(n1067), .B(n1068), .Z(G69) );
XOR2_X1 U767 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U768 ( .A1(G953), .A2(n1071), .ZN(n1070) );
NAND2_X1 U769 ( .A1(G898), .A2(G224), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
NAND2_X1 U771 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1075), .B(n1076), .Z(n1072) );
XOR2_X1 U773 ( .A(n1077), .B(G122), .Z(n1075) );
NAND2_X1 U774 ( .A1(KEYINPUT62), .A2(n1078), .ZN(n1077) );
XOR2_X1 U775 ( .A(G113), .B(n1079), .Z(n1078) );
AND2_X1 U776 ( .A1(n1080), .A2(n979), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1081), .A2(n1082), .ZN(G66) );
XOR2_X1 U778 ( .A(n1083), .B(n1084), .Z(n1082) );
AND2_X1 U779 ( .A1(G217), .A2(n1085), .ZN(n1083) );
NOR2_X1 U780 ( .A1(G952), .A2(n1086), .ZN(n1081) );
XOR2_X1 U781 ( .A(n979), .B(KEYINPUT5), .Z(n1086) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(G63) );
XOR2_X1 U783 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U784 ( .A1(KEYINPUT32), .A2(n1091), .ZN(n1090) );
NAND2_X1 U785 ( .A1(n1085), .A2(G478), .ZN(n1089) );
NOR2_X1 U786 ( .A1(n1087), .A2(n1092), .ZN(G60) );
NOR3_X1 U787 ( .A1(n1041), .A2(n1093), .A3(n1094), .ZN(n1092) );
AND3_X1 U788 ( .A1(n1095), .A2(G475), .A3(n1085), .ZN(n1094) );
INV_X1 U789 ( .A(n1096), .ZN(n1085) );
NOR2_X1 U790 ( .A1(n1097), .A2(n1095), .ZN(n1093) );
AND2_X1 U791 ( .A1(n1098), .A2(G475), .ZN(n1097) );
XOR2_X1 U792 ( .A(G104), .B(n1099), .Z(G6) );
NOR2_X1 U793 ( .A1(n1087), .A2(n1100), .ZN(G57) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U795 ( .A(KEYINPUT29), .B(n1103), .Z(n1102) );
AND2_X1 U796 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
XNOR2_X1 U798 ( .A(n1106), .B(n1107), .ZN(n1105) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND4_X1 U800 ( .A1(KEYINPUT44), .A2(G472), .A3(n1110), .A4(n1098), .ZN(n1109) );
XOR2_X1 U801 ( .A(KEYINPUT53), .B(G902), .Z(n1110) );
NAND2_X1 U802 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
OR2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U804 ( .A(n1115), .B(KEYINPUT22), .Z(n1111) );
NAND2_X1 U805 ( .A1(n1114), .A2(n1113), .ZN(n1115) );
NOR3_X1 U806 ( .A1(n1116), .A2(n1087), .A3(n1117), .ZN(G54) );
NOR3_X1 U807 ( .A1(n1118), .A2(n1119), .A3(n1096), .ZN(n1117) );
NOR2_X1 U808 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
XNOR2_X1 U809 ( .A(KEYINPUT2), .B(n1118), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1122), .B(n1123), .Z(n1118) );
XNOR2_X1 U811 ( .A(n1066), .B(n1124), .ZN(n1123) );
XNOR2_X1 U812 ( .A(G140), .B(n1125), .ZN(n1124) );
XOR2_X1 U813 ( .A(n1126), .B(n1127), .Z(n1122) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U815 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1129) );
AND2_X1 U816 ( .A1(KEYINPUT16), .A2(G110), .ZN(n1128) );
NOR2_X1 U817 ( .A1(n1119), .A2(n1096), .ZN(n1120) );
NAND2_X1 U818 ( .A1(G902), .A2(n1098), .ZN(n1096) );
INV_X1 U819 ( .A(n983), .ZN(n1098) );
INV_X1 U820 ( .A(G469), .ZN(n1119) );
NOR2_X1 U821 ( .A1(n1130), .A2(n1131), .ZN(G51) );
XNOR2_X1 U822 ( .A(n1087), .B(KEYINPUT61), .ZN(n1131) );
NOR2_X1 U823 ( .A1(n979), .A2(G952), .ZN(n1087) );
XOR2_X1 U824 ( .A(n1132), .B(n1133), .Z(n1130) );
XOR2_X1 U825 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U826 ( .A(n1136), .B(KEYINPUT25), .Z(n1135) );
NAND3_X1 U827 ( .A1(n1050), .A2(n1137), .A3(G902), .ZN(n1134) );
XOR2_X1 U828 ( .A(KEYINPUT30), .B(n983), .Z(n1137) );
NOR2_X1 U829 ( .A1(n1080), .A2(n1059), .ZN(n983) );
NAND4_X1 U830 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1059) );
AND4_X1 U831 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
AND2_X1 U832 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
NAND2_X1 U833 ( .A1(n1148), .A2(n1016), .ZN(n1139) );
XOR2_X1 U834 ( .A(n1149), .B(KEYINPUT15), .Z(n1148) );
NAND4_X1 U835 ( .A1(n1021), .A2(n991), .A3(n1150), .A4(n1151), .ZN(n1149) );
XOR2_X1 U836 ( .A(KEYINPUT63), .B(n993), .Z(n1150) );
OR2_X1 U837 ( .A1(n1152), .A2(n1007), .ZN(n1138) );
NAND2_X1 U838 ( .A1(n1153), .A2(n1154), .ZN(n1080) );
NOR4_X1 U839 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
NOR4_X1 U840 ( .A1(n977), .A2(n1159), .A3(n1099), .A4(n1160), .ZN(n1153) );
AND3_X1 U841 ( .A1(n1025), .A2(n1161), .A3(n992), .ZN(n1160) );
AND3_X1 U842 ( .A1(n1161), .A2(n994), .A3(n1021), .ZN(n1099) );
AND3_X1 U843 ( .A1(n1020), .A2(n994), .A3(n1161), .ZN(n977) );
INV_X1 U844 ( .A(n1162), .ZN(n1050) );
XOR2_X1 U845 ( .A(n1163), .B(n1164), .Z(n1132) );
NAND2_X1 U846 ( .A1(KEYINPUT12), .A2(n1165), .ZN(n1163) );
XOR2_X1 U847 ( .A(G146), .B(n1166), .Z(G48) );
NOR2_X1 U848 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
AND2_X1 U849 ( .A1(KEYINPUT23), .A2(n1147), .ZN(n1168) );
NOR2_X1 U850 ( .A1(KEYINPUT43), .A2(n1147), .ZN(n1167) );
NAND3_X1 U851 ( .A1(n1021), .A2(n1016), .A3(n1169), .ZN(n1147) );
XOR2_X1 U852 ( .A(n1170), .B(n1146), .Z(G45) );
NAND4_X1 U853 ( .A1(n1171), .A2(n1016), .A3(n1172), .A4(n1173), .ZN(n1146) );
XNOR2_X1 U854 ( .A(G140), .B(n1145), .ZN(G42) );
NAND4_X1 U855 ( .A1(n990), .A2(n1174), .A3(n1021), .A4(n993), .ZN(n1145) );
XOR2_X1 U856 ( .A(n1175), .B(G137), .Z(G39) );
NAND2_X1 U857 ( .A1(KEYINPUT38), .A2(n1144), .ZN(n1175) );
NAND3_X1 U858 ( .A1(n1169), .A2(n992), .A3(n990), .ZN(n1144) );
XNOR2_X1 U859 ( .A(G134), .B(n1143), .ZN(G36) );
NAND3_X1 U860 ( .A1(n1171), .A2(n1020), .A3(n990), .ZN(n1143) );
INV_X1 U861 ( .A(n1007), .ZN(n990) );
XOR2_X1 U862 ( .A(G131), .B(n1176), .Z(G33) );
NOR2_X1 U863 ( .A1(n1177), .A2(n1007), .ZN(n1176) );
NAND2_X1 U864 ( .A1(n1015), .A2(n1178), .ZN(n1007) );
XOR2_X1 U865 ( .A(n1152), .B(KEYINPUT18), .Z(n1177) );
NAND2_X1 U866 ( .A1(n1171), .A2(n1021), .ZN(n1152) );
AND2_X1 U867 ( .A1(n1174), .A2(n1025), .ZN(n1171) );
XNOR2_X1 U868 ( .A(G128), .B(n1142), .ZN(G30) );
NAND3_X1 U869 ( .A1(n1020), .A2(n1016), .A3(n1169), .ZN(n1142) );
AND3_X1 U870 ( .A1(n1043), .A2(n1179), .A3(n1174), .ZN(n1169) );
AND3_X1 U871 ( .A1(n1151), .A2(n1001), .A3(n1002), .ZN(n1174) );
XNOR2_X1 U872 ( .A(G101), .B(n1180), .ZN(G3) );
NAND4_X1 U873 ( .A1(KEYINPUT57), .A2(n1025), .A3(n1161), .A4(n1181), .ZN(n1180) );
XOR2_X1 U874 ( .A(KEYINPUT34), .B(n992), .Z(n1181) );
XOR2_X1 U875 ( .A(n1182), .B(n1183), .Z(G27) );
NAND3_X1 U876 ( .A1(n1021), .A2(n991), .A3(n1184), .ZN(n1183) );
AND3_X1 U877 ( .A1(n993), .A2(n1151), .A3(n1016), .ZN(n1184) );
NAND2_X1 U878 ( .A1(n1022), .A2(n1185), .ZN(n1151) );
NAND4_X1 U879 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1055), .ZN(n1185) );
INV_X1 U880 ( .A(G900), .ZN(n1055) );
XNOR2_X1 U881 ( .A(n1159), .B(n1187), .ZN(G24) );
XOR2_X1 U882 ( .A(KEYINPUT4), .B(G122), .Z(n1187) );
AND4_X1 U883 ( .A1(n1188), .A2(n994), .A3(n1172), .A4(n1173), .ZN(n1159) );
NOR2_X1 U884 ( .A1(n1179), .A2(n1043), .ZN(n994) );
XNOR2_X1 U885 ( .A(n1158), .B(n1189), .ZN(G21) );
XOR2_X1 U886 ( .A(KEYINPUT9), .B(G119), .Z(n1189) );
AND4_X1 U887 ( .A1(n1188), .A2(n992), .A3(n1043), .A4(n1179), .ZN(n1158) );
INV_X1 U888 ( .A(n1190), .ZN(n1043) );
XOR2_X1 U889 ( .A(G116), .B(n1157), .Z(G18) );
AND3_X1 U890 ( .A1(n1188), .A2(n1020), .A3(n1025), .ZN(n1157) );
NOR2_X1 U891 ( .A1(n1173), .A2(n1191), .ZN(n1020) );
XOR2_X1 U892 ( .A(n1156), .B(n1192), .Z(G15) );
NOR2_X1 U893 ( .A1(KEYINPUT56), .A2(n1193), .ZN(n1192) );
AND3_X1 U894 ( .A1(n1021), .A2(n1188), .A3(n1025), .ZN(n1156) );
NOR2_X1 U895 ( .A1(n1179), .A2(n1190), .ZN(n1025) );
AND3_X1 U896 ( .A1(n1016), .A2(n1194), .A3(n991), .ZN(n1188) );
AND2_X1 U897 ( .A1(n1006), .A2(n1001), .ZN(n991) );
XNOR2_X1 U898 ( .A(n1002), .B(KEYINPUT58), .ZN(n1006) );
AND2_X1 U899 ( .A1(n1191), .A2(n1173), .ZN(n1021) );
INV_X1 U900 ( .A(n1172), .ZN(n1191) );
XOR2_X1 U901 ( .A(n1155), .B(n1195), .Z(G12) );
NOR2_X1 U902 ( .A1(KEYINPUT48), .A2(n1196), .ZN(n1195) );
AND3_X1 U903 ( .A1(n993), .A2(n1161), .A3(n992), .ZN(n1155) );
NOR2_X1 U904 ( .A1(n1172), .A2(n1173), .ZN(n992) );
XOR2_X1 U905 ( .A(n1041), .B(G475), .Z(n1173) );
NOR2_X1 U906 ( .A1(n1095), .A2(G902), .ZN(n1041) );
XOR2_X1 U907 ( .A(n1197), .B(n1198), .Z(n1095) );
XOR2_X1 U908 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U909 ( .A(n1201), .B(n1202), .ZN(n1200) );
NOR2_X1 U910 ( .A1(KEYINPUT24), .A2(n1203), .ZN(n1202) );
XOR2_X1 U911 ( .A(n1204), .B(n1205), .Z(n1199) );
NOR3_X1 U912 ( .A1(n1206), .A2(G237), .A3(n1207), .ZN(n1205) );
INV_X1 U913 ( .A(G214), .ZN(n1207) );
XOR2_X1 U914 ( .A(KEYINPUT7), .B(G953), .Z(n1206) );
NAND2_X1 U915 ( .A1(KEYINPUT8), .A2(n1170), .ZN(n1204) );
XOR2_X1 U916 ( .A(n1208), .B(n1209), .Z(n1197) );
XOR2_X1 U917 ( .A(KEYINPUT3), .B(G140), .Z(n1209) );
XNOR2_X1 U918 ( .A(G104), .B(G131), .ZN(n1208) );
XOR2_X1 U919 ( .A(n1039), .B(G478), .Z(n1172) );
NOR2_X1 U920 ( .A1(n1091), .A2(G902), .ZN(n1039) );
XOR2_X1 U921 ( .A(n1210), .B(n1211), .Z(n1091) );
XNOR2_X1 U922 ( .A(n1212), .B(n1213), .ZN(n1211) );
NAND2_X1 U923 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
XOR2_X1 U924 ( .A(KEYINPUT59), .B(KEYINPUT26), .Z(n1215) );
XNOR2_X1 U925 ( .A(G134), .B(n1216), .ZN(n1214) );
XOR2_X1 U926 ( .A(n1217), .B(n1218), .Z(n1210) );
XOR2_X1 U927 ( .A(G122), .B(G107), .Z(n1218) );
NAND2_X1 U928 ( .A1(G217), .A2(n1219), .ZN(n1217) );
AND4_X1 U929 ( .A1(n1002), .A2(n1016), .A3(n1001), .A4(n1194), .ZN(n1161) );
NAND2_X1 U930 ( .A1(n1220), .A2(n1022), .ZN(n1194) );
NAND3_X1 U931 ( .A1(n1186), .A2(n979), .A3(G952), .ZN(n1022) );
XOR2_X1 U932 ( .A(n1221), .B(KEYINPUT51), .Z(n1220) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1074), .ZN(n1221) );
INV_X1 U934 ( .A(G898), .ZN(n1074) );
NAND2_X1 U935 ( .A1(G237), .A2(G234), .ZN(n1186) );
NAND2_X1 U936 ( .A1(G221), .A2(n1222), .ZN(n1001) );
NOR2_X1 U937 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
INV_X1 U938 ( .A(n1178), .ZN(n1014) );
NAND2_X1 U939 ( .A1(G214), .A2(n1223), .ZN(n1178) );
XOR2_X1 U940 ( .A(n1049), .B(n1224), .Z(n1015) );
NOR2_X1 U941 ( .A1(KEYINPUT39), .A2(n1162), .ZN(n1224) );
NAND2_X1 U942 ( .A1(G210), .A2(n1223), .ZN(n1162) );
NAND2_X1 U943 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NAND2_X1 U944 ( .A1(n1227), .A2(n1225), .ZN(n1049) );
XOR2_X1 U945 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U946 ( .A(n1164), .B(n1165), .Z(n1229) );
XNOR2_X1 U947 ( .A(G125), .B(n1114), .ZN(n1165) );
XNOR2_X1 U948 ( .A(n1230), .B(n1076), .ZN(n1164) );
XOR2_X1 U949 ( .A(n1231), .B(n1232), .Z(n1076) );
XOR2_X1 U950 ( .A(G110), .B(n1233), .Z(n1232) );
NOR2_X1 U951 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1233) );
XOR2_X1 U952 ( .A(n1079), .B(n1203), .Z(n1230) );
XOR2_X1 U953 ( .A(n1193), .B(G122), .Z(n1203) );
XOR2_X1 U954 ( .A(n1136), .B(KEYINPUT28), .Z(n1228) );
NAND2_X1 U955 ( .A1(n1234), .A2(n979), .ZN(n1136) );
XOR2_X1 U956 ( .A(KEYINPUT21), .B(G224), .Z(n1234) );
XOR2_X1 U957 ( .A(n1048), .B(n1235), .Z(n1002) );
NOR2_X1 U958 ( .A1(G469), .A2(n1236), .ZN(n1235) );
XNOR2_X1 U959 ( .A(KEYINPUT47), .B(KEYINPUT36), .ZN(n1236) );
NAND2_X1 U960 ( .A1(n1237), .A2(n1225), .ZN(n1048) );
XOR2_X1 U961 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U962 ( .A(n1240), .B(n1125), .Z(n1239) );
XOR2_X1 U963 ( .A(n1113), .B(n1241), .Z(n1125) );
NOR2_X1 U964 ( .A1(G953), .A2(n1054), .ZN(n1241) );
INV_X1 U965 ( .A(G227), .ZN(n1054) );
NAND2_X1 U966 ( .A1(n1242), .A2(KEYINPUT42), .ZN(n1240) );
XOR2_X1 U967 ( .A(n1066), .B(n1243), .Z(n1242) );
XNOR2_X1 U968 ( .A(n1244), .B(KEYINPUT52), .ZN(n1243) );
NAND2_X1 U969 ( .A1(KEYINPUT14), .A2(n1126), .ZN(n1244) );
XNOR2_X1 U970 ( .A(G101), .B(n1231), .ZN(n1126) );
XOR2_X1 U971 ( .A(G104), .B(G107), .Z(n1231) );
XOR2_X1 U972 ( .A(n1245), .B(n1216), .Z(n1066) );
XOR2_X1 U973 ( .A(G128), .B(G143), .Z(n1216) );
XOR2_X1 U974 ( .A(n1246), .B(KEYINPUT33), .Z(n1245) );
XOR2_X1 U975 ( .A(G110), .B(n1247), .Z(n1238) );
XOR2_X1 U976 ( .A(KEYINPUT1), .B(G140), .Z(n1247) );
AND2_X1 U977 ( .A1(n1190), .A2(n1179), .ZN(n993) );
XNOR2_X1 U978 ( .A(n1047), .B(n1045), .ZN(n1179) );
NAND2_X1 U979 ( .A1(n1248), .A2(n1222), .ZN(n1045) );
NAND2_X1 U980 ( .A1(G234), .A2(n1225), .ZN(n1222) );
XOR2_X1 U981 ( .A(KEYINPUT35), .B(G217), .Z(n1248) );
NOR2_X1 U982 ( .A1(n1084), .A2(G902), .ZN(n1047) );
XNOR2_X1 U983 ( .A(n1249), .B(n1250), .ZN(n1084) );
XOR2_X1 U984 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U985 ( .A(G137), .B(n1196), .Z(n1252) );
INV_X1 U986 ( .A(G110), .ZN(n1196) );
NAND2_X1 U987 ( .A1(KEYINPUT11), .A2(n1253), .ZN(n1251) );
XOR2_X1 U988 ( .A(G128), .B(G119), .Z(n1253) );
XOR2_X1 U989 ( .A(n1254), .B(n1201), .Z(n1249) );
XOR2_X1 U990 ( .A(n1182), .B(n1246), .Z(n1201) );
INV_X1 U991 ( .A(G125), .ZN(n1182) );
XOR2_X1 U992 ( .A(n1255), .B(n1256), .Z(n1254) );
NOR2_X1 U993 ( .A1(G140), .A2(KEYINPUT10), .ZN(n1256) );
NAND2_X1 U994 ( .A1(n1219), .A2(G221), .ZN(n1255) );
AND2_X1 U995 ( .A1(G234), .A2(n979), .ZN(n1219) );
XOR2_X1 U996 ( .A(n1257), .B(G472), .Z(n1190) );
NAND2_X1 U997 ( .A1(n1258), .A2(n1225), .ZN(n1257) );
INV_X1 U998 ( .A(G902), .ZN(n1225) );
XOR2_X1 U999 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U1000 ( .A(n1261), .B(n1104), .Z(n1260) );
XNOR2_X1 U1001 ( .A(n1262), .B(G101), .ZN(n1104) );
NAND3_X1 U1002 ( .A1(n1226), .A2(n979), .A3(G210), .ZN(n1262) );
INV_X1 U1003 ( .A(G953), .ZN(n979) );
INV_X1 U1004 ( .A(G237), .ZN(n1226) );
INV_X1 U1005 ( .A(n1106), .ZN(n1261) );
XNOR2_X1 U1006 ( .A(n1079), .B(n1263), .ZN(n1106) );
XNOR2_X1 U1007 ( .A(n1264), .B(KEYINPUT46), .ZN(n1263) );
NAND2_X1 U1008 ( .A1(KEYINPUT20), .A2(n1193), .ZN(n1264) );
INV_X1 U1009 ( .A(G113), .ZN(n1193) );
XOR2_X1 U1010 ( .A(G119), .B(n1213), .Z(n1079) );
XOR2_X1 U1011 ( .A(G116), .B(KEYINPUT37), .Z(n1213) );
XNOR2_X1 U1012 ( .A(n1265), .B(n1114), .ZN(n1259) );
XNOR2_X1 U1013 ( .A(n1266), .B(n1267), .ZN(n1114) );
NOR2_X1 U1014 ( .A1(G128), .A2(KEYINPUT55), .ZN(n1267) );
NAND2_X1 U1015 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
NAND2_X1 U1016 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
INV_X1 U1017 ( .A(KEYINPUT31), .ZN(n1271) );
XOR2_X1 U1018 ( .A(n1170), .B(G146), .Z(n1270) );
INV_X1 U1019 ( .A(G143), .ZN(n1170) );
NAND3_X1 U1020 ( .A1(G143), .A2(n1246), .A3(KEYINPUT31), .ZN(n1268) );
INV_X1 U1021 ( .A(G146), .ZN(n1246) );
NAND2_X1 U1022 ( .A1(KEYINPUT40), .A2(n1272), .ZN(n1265) );
INV_X1 U1023 ( .A(n1113), .ZN(n1272) );
NAND2_X1 U1024 ( .A1(n1273), .A2(n1274), .ZN(n1113) );
NAND2_X1 U1025 ( .A1(G131), .A2(n1065), .ZN(n1274) );
XOR2_X1 U1026 ( .A(n1275), .B(KEYINPUT27), .Z(n1273) );
OR2_X1 U1027 ( .A1(n1065), .A2(G131), .ZN(n1275) );
XOR2_X1 U1028 ( .A(G134), .B(G137), .Z(n1065) );
endmodule


