//Key = 1101011001101000111000111110001010111001101101111100010100110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326;

XNOR2_X1 U733 ( .A(G107), .B(n1004), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
NOR2_X1 U736 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U737 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
XOR2_X1 U738 ( .A(KEYINPUT56), .B(n1015), .Z(n1014) );
NOR2_X1 U739 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U740 ( .A(n1018), .ZN(n1016) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1017), .ZN(n1013) );
NAND3_X1 U742 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1017) );
NAND4_X1 U743 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1007) );
NAND3_X1 U744 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1024) );
INV_X1 U745 ( .A(KEYINPUT16), .ZN(n1028) );
NAND4_X1 U746 ( .A1(n1030), .A2(n1022), .A3(n1021), .A4(n1031), .ZN(n1027) );
NAND3_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1022), .ZN(n1023) );
INV_X1 U748 ( .A(n1033), .ZN(n1022) );
NAND2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND3_X1 U750 ( .A1(n1020), .A2(n1036), .A3(n1037), .ZN(n1035) );
OR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1021), .A2(n1040), .ZN(n1034) );
NAND3_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1037), .A2(n1044), .ZN(n1043) );
NAND2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U757 ( .A1(n1030), .A2(n1029), .A3(KEYINPUT16), .ZN(n1042) );
XNOR2_X1 U758 ( .A(n1020), .B(KEYINPUT58), .ZN(n1030) );
NAND3_X1 U759 ( .A1(n1049), .A2(n1020), .A3(n1050), .ZN(n1041) );
AND3_X1 U760 ( .A1(n1025), .A2(n1026), .A3(n1051), .ZN(n1005) );
NAND4_X1 U761 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1025) );
NOR4_X1 U762 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
XOR2_X1 U763 ( .A(KEYINPUT62), .B(n1060), .Z(n1059) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XNOR2_X1 U765 ( .A(G469), .B(n1063), .ZN(n1056) );
NOR2_X1 U766 ( .A1(n1064), .A2(KEYINPUT54), .ZN(n1063) );
NOR3_X1 U767 ( .A1(n1047), .A2(n1065), .A3(n1050), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1062), .A2(n1061), .ZN(n1053) );
XNOR2_X1 U769 ( .A(KEYINPUT4), .B(n1066), .ZN(n1062) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1052) );
XOR2_X1 U771 ( .A(n1069), .B(n1070), .Z(G72) );
XOR2_X1 U772 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U773 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U774 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U775 ( .A(n1026), .B(KEYINPUT53), .Z(n1075) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(n1073) );
XOR2_X1 U777 ( .A(KEYINPUT60), .B(n1079), .Z(n1078) );
XNOR2_X1 U778 ( .A(n1080), .B(n1081), .ZN(n1077) );
NAND2_X1 U779 ( .A1(G953), .A2(n1082), .ZN(n1071) );
XOR2_X1 U780 ( .A(KEYINPUT34), .B(n1083), .Z(n1082) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1083) );
NOR2_X1 U782 ( .A1(n1084), .A2(G953), .ZN(n1069) );
XOR2_X1 U783 ( .A(n1085), .B(n1086), .Z(G69) );
NAND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U785 ( .A1(G898), .A2(G224), .ZN(n1088) );
XOR2_X1 U786 ( .A(n1026), .B(KEYINPUT40), .Z(n1087) );
NAND2_X1 U787 ( .A1(KEYINPUT59), .A2(n1089), .ZN(n1085) );
XOR2_X1 U788 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U789 ( .A1(n1092), .A2(G953), .ZN(n1091) );
NOR2_X1 U790 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
XNOR2_X1 U791 ( .A(n1095), .B(n1096), .ZN(n1094) );
XOR2_X1 U792 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U793 ( .A1(G898), .A2(n1026), .ZN(n1093) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U796 ( .A1(KEYINPUT23), .A2(n1103), .ZN(n1102) );
NAND2_X1 U797 ( .A1(n1104), .A2(G217), .ZN(n1101) );
NOR2_X1 U798 ( .A1(n1099), .A2(n1105), .ZN(G63) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR3_X1 U800 ( .A1(n1108), .A2(KEYINPUT7), .A3(n1109), .ZN(n1106) );
INV_X1 U801 ( .A(G478), .ZN(n1109) );
NOR2_X1 U802 ( .A1(n1099), .A2(n1110), .ZN(G60) );
XOR2_X1 U803 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U804 ( .A1(n1104), .A2(G475), .ZN(n1112) );
NAND2_X1 U805 ( .A1(KEYINPUT1), .A2(n1113), .ZN(n1111) );
INV_X1 U806 ( .A(n1114), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1115), .B(n1116), .Z(G6) );
NOR2_X1 U808 ( .A1(KEYINPUT57), .A2(n1117), .ZN(n1116) );
XOR2_X1 U809 ( .A(n1118), .B(KEYINPUT50), .Z(n1117) );
NOR2_X1 U810 ( .A1(n1099), .A2(n1119), .ZN(G57) );
XOR2_X1 U811 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U812 ( .A(n1081), .B(n1122), .ZN(n1121) );
XOR2_X1 U813 ( .A(n1123), .B(n1124), .Z(n1120) );
NOR2_X1 U814 ( .A1(n1061), .A2(n1108), .ZN(n1124) );
INV_X1 U815 ( .A(G472), .ZN(n1061) );
NOR2_X1 U816 ( .A1(n1099), .A2(n1125), .ZN(G54) );
XOR2_X1 U817 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U818 ( .A(n1128), .B(n1129), .ZN(n1127) );
XOR2_X1 U819 ( .A(n1130), .B(n1131), .Z(n1126) );
AND2_X1 U820 ( .A1(G469), .A2(n1104), .ZN(n1131) );
INV_X1 U821 ( .A(n1108), .ZN(n1104) );
NOR2_X1 U822 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
XOR2_X1 U823 ( .A(KEYINPUT41), .B(n1134), .Z(n1133) );
AND2_X1 U824 ( .A1(n1080), .A2(n1135), .ZN(n1134) );
NOR2_X1 U825 ( .A1(n1080), .A2(n1135), .ZN(n1132) );
XNOR2_X1 U826 ( .A(n1136), .B(KEYINPUT33), .ZN(n1135) );
NOR2_X1 U827 ( .A1(n1099), .A2(n1137), .ZN(G51) );
XNOR2_X1 U828 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U829 ( .A1(n1140), .A2(n1108), .ZN(n1139) );
NAND2_X1 U830 ( .A1(G902), .A2(n1141), .ZN(n1108) );
NAND2_X1 U831 ( .A1(n1092), .A2(n1084), .ZN(n1141) );
INV_X1 U832 ( .A(n1010), .ZN(n1084) );
NAND2_X1 U833 ( .A1(n1142), .A2(n1143), .ZN(n1010) );
NOR4_X1 U834 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
AND4_X1 U835 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1142) );
INV_X1 U836 ( .A(n1008), .ZN(n1092) );
NAND2_X1 U837 ( .A1(n1152), .A2(n1153), .ZN(n1008) );
NOR4_X1 U838 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1115), .ZN(n1153) );
AND3_X1 U839 ( .A1(n1031), .A2(n1157), .A3(n1038), .ZN(n1115) );
INV_X1 U840 ( .A(n1158), .ZN(n1156) );
INV_X1 U841 ( .A(n1159), .ZN(n1154) );
AND4_X1 U842 ( .A1(n1004), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1152) );
OR3_X1 U843 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
XOR2_X1 U844 ( .A(KEYINPUT29), .B(n1166), .Z(n1163) );
NAND3_X1 U845 ( .A1(n1157), .A2(n1039), .A3(n1031), .ZN(n1004) );
AND2_X1 U846 ( .A1(n1167), .A2(n1051), .ZN(n1099) );
INV_X1 U847 ( .A(G952), .ZN(n1051) );
XOR2_X1 U848 ( .A(KEYINPUT31), .B(G953), .Z(n1167) );
XOR2_X1 U849 ( .A(G146), .B(n1168), .Z(G48) );
NOR2_X1 U850 ( .A1(KEYINPUT8), .A2(n1151), .ZN(n1168) );
NAND3_X1 U851 ( .A1(n1038), .A2(n1029), .A3(n1169), .ZN(n1151) );
XOR2_X1 U852 ( .A(n1170), .B(n1147), .Z(G45) );
AND3_X1 U853 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1147) );
NOR3_X1 U854 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NAND2_X1 U855 ( .A1(KEYINPUT12), .A2(n1177), .ZN(n1170) );
INV_X1 U856 ( .A(G143), .ZN(n1177) );
XOR2_X1 U857 ( .A(G140), .B(n1146), .Z(G42) );
AND4_X1 U858 ( .A1(n1037), .A2(n1171), .A3(n1038), .A4(n1018), .ZN(n1146) );
XOR2_X1 U859 ( .A(G137), .B(n1145), .Z(G39) );
AND3_X1 U860 ( .A1(n1037), .A2(n1021), .A3(n1169), .ZN(n1145) );
XOR2_X1 U861 ( .A(n1144), .B(n1178), .Z(G36) );
NOR2_X1 U862 ( .A1(KEYINPUT38), .A2(n1179), .ZN(n1178) );
NOR3_X1 U863 ( .A1(n1180), .A2(n1165), .A3(n1012), .ZN(n1144) );
INV_X1 U864 ( .A(n1037), .ZN(n1012) );
NAND2_X1 U865 ( .A1(n1181), .A2(n1182), .ZN(G33) );
NAND2_X1 U866 ( .A1(G131), .A2(n1150), .ZN(n1182) );
XOR2_X1 U867 ( .A(KEYINPUT46), .B(n1183), .Z(n1181) );
NOR2_X1 U868 ( .A1(G131), .A2(n1150), .ZN(n1183) );
NAND4_X1 U869 ( .A1(n1037), .A2(n1171), .A3(n1038), .A4(n1172), .ZN(n1150) );
NOR2_X1 U870 ( .A1(n1184), .A2(n1050), .ZN(n1037) );
XNOR2_X1 U871 ( .A(G128), .B(n1149), .ZN(G30) );
NAND3_X1 U872 ( .A1(n1039), .A2(n1029), .A3(n1169), .ZN(n1149) );
AND3_X1 U873 ( .A1(n1185), .A2(n1057), .A3(n1171), .ZN(n1169) );
INV_X1 U874 ( .A(n1180), .ZN(n1171) );
NAND2_X1 U875 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NAND2_X1 U876 ( .A1(n1188), .A2(n1189), .ZN(G3) );
OR2_X1 U877 ( .A1(n1158), .A2(G101), .ZN(n1189) );
XOR2_X1 U878 ( .A(n1190), .B(KEYINPUT20), .Z(n1188) );
NAND2_X1 U879 ( .A1(G101), .A2(n1158), .ZN(n1190) );
NAND3_X1 U880 ( .A1(n1021), .A2(n1157), .A3(n1172), .ZN(n1158) );
XOR2_X1 U881 ( .A(n1191), .B(n1148), .Z(G27) );
NAND4_X1 U882 ( .A1(n1038), .A2(n1192), .A3(n1018), .A4(n1187), .ZN(n1148) );
NAND2_X1 U883 ( .A1(n1033), .A2(n1193), .ZN(n1187) );
NAND4_X1 U884 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1076), .ZN(n1193) );
INV_X1 U885 ( .A(G900), .ZN(n1076) );
XOR2_X1 U886 ( .A(n1195), .B(G122), .Z(G24) );
NAND2_X1 U887 ( .A1(KEYINPUT61), .A2(n1161), .ZN(n1195) );
NAND4_X1 U888 ( .A1(n1196), .A2(n1031), .A3(n1197), .A4(n1198), .ZN(n1161) );
NOR2_X1 U889 ( .A1(n1057), .A2(n1185), .ZN(n1031) );
XNOR2_X1 U890 ( .A(G119), .B(n1160), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1185), .A2(n1196), .A3(n1021), .A4(n1057), .ZN(n1160) );
XOR2_X1 U892 ( .A(n1199), .B(n1200), .Z(G18) );
XOR2_X1 U893 ( .A(KEYINPUT13), .B(G116), .Z(n1200) );
NOR2_X1 U894 ( .A1(n1201), .A2(n1165), .ZN(n1199) );
NAND2_X1 U895 ( .A1(n1172), .A2(n1039), .ZN(n1165) );
NOR2_X1 U896 ( .A1(n1197), .A2(n1175), .ZN(n1039) );
INV_X1 U897 ( .A(n1176), .ZN(n1197) );
XOR2_X1 U898 ( .A(G113), .B(n1155), .Z(G15) );
AND3_X1 U899 ( .A1(n1172), .A2(n1196), .A3(n1038), .ZN(n1155) );
NOR2_X1 U900 ( .A1(n1198), .A2(n1176), .ZN(n1038) );
INV_X1 U901 ( .A(n1175), .ZN(n1198) );
INV_X1 U902 ( .A(n1201), .ZN(n1196) );
NAND2_X1 U903 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
INV_X1 U904 ( .A(n1164), .ZN(n1192) );
NAND2_X1 U905 ( .A1(n1020), .A2(n1029), .ZN(n1164) );
NOR2_X1 U906 ( .A1(n1203), .A2(n1047), .ZN(n1020) );
INV_X1 U907 ( .A(n1048), .ZN(n1203) );
INV_X1 U908 ( .A(n1019), .ZN(n1172) );
NAND2_X1 U909 ( .A1(n1185), .A2(n1204), .ZN(n1019) );
XOR2_X1 U910 ( .A(n1205), .B(n1159), .Z(G12) );
NAND3_X1 U911 ( .A1(n1021), .A2(n1157), .A3(n1018), .ZN(n1159) );
NOR2_X1 U912 ( .A1(n1185), .A2(n1204), .ZN(n1018) );
INV_X1 U913 ( .A(n1057), .ZN(n1204) );
NAND3_X1 U914 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1057) );
OR2_X1 U915 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND3_X1 U916 ( .A1(n1210), .A2(n1209), .A3(n1211), .ZN(n1207) );
NAND2_X1 U917 ( .A1(G217), .A2(n1212), .ZN(n1209) );
INV_X1 U918 ( .A(n1103), .ZN(n1210) );
XOR2_X1 U919 ( .A(n1213), .B(n1214), .Z(n1103) );
XOR2_X1 U920 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U921 ( .A(n1217), .B(n1218), .ZN(n1216) );
NAND2_X1 U922 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
NAND2_X1 U923 ( .A1(G140), .A2(n1191), .ZN(n1220) );
XOR2_X1 U924 ( .A(KEYINPUT32), .B(n1221), .Z(n1219) );
NOR2_X1 U925 ( .A1(G140), .A2(n1191), .ZN(n1221) );
INV_X1 U926 ( .A(G125), .ZN(n1191) );
XOR2_X1 U927 ( .A(n1222), .B(n1223), .Z(n1213) );
XOR2_X1 U928 ( .A(KEYINPUT27), .B(G110), .Z(n1223) );
NAND2_X1 U929 ( .A1(KEYINPUT6), .A2(n1224), .ZN(n1222) );
XOR2_X1 U930 ( .A(G137), .B(n1225), .Z(n1224) );
NOR4_X1 U931 ( .A1(KEYINPUT44), .A2(G953), .A3(n1226), .A4(n1212), .ZN(n1225) );
INV_X1 U932 ( .A(G234), .ZN(n1212) );
INV_X1 U933 ( .A(G221), .ZN(n1226) );
NAND2_X1 U934 ( .A1(G902), .A2(G217), .ZN(n1206) );
XOR2_X1 U935 ( .A(n1066), .B(n1227), .Z(n1185) );
XOR2_X1 U936 ( .A(KEYINPUT39), .B(G472), .Z(n1227) );
NAND2_X1 U937 ( .A1(n1228), .A2(n1211), .ZN(n1066) );
XNOR2_X1 U938 ( .A(n1229), .B(n1122), .ZN(n1228) );
XOR2_X1 U939 ( .A(n1230), .B(n1231), .Z(n1122) );
XOR2_X1 U940 ( .A(n1232), .B(n1218), .Z(n1231) );
XOR2_X1 U941 ( .A(n1233), .B(n1234), .Z(n1230) );
XOR2_X1 U942 ( .A(G113), .B(G101), .Z(n1234) );
NAND2_X1 U943 ( .A1(G210), .A2(n1235), .ZN(n1233) );
NAND2_X1 U944 ( .A1(n1236), .A2(KEYINPUT43), .ZN(n1229) );
XNOR2_X1 U945 ( .A(n1081), .B(n1237), .ZN(n1236) );
NOR2_X1 U946 ( .A1(KEYINPUT2), .A2(n1123), .ZN(n1237) );
NOR3_X1 U947 ( .A1(n1174), .A2(n1166), .A3(n1045), .ZN(n1157) );
INV_X1 U948 ( .A(n1186), .ZN(n1045) );
NOR2_X1 U949 ( .A1(n1048), .A2(n1047), .ZN(n1186) );
AND2_X1 U950 ( .A1(G221), .A2(n1238), .ZN(n1047) );
NAND2_X1 U951 ( .A1(G234), .A2(n1211), .ZN(n1238) );
XOR2_X1 U952 ( .A(n1239), .B(n1064), .Z(n1048) );
AND2_X1 U953 ( .A1(n1240), .A2(n1211), .ZN(n1064) );
XOR2_X1 U954 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U955 ( .A(n1136), .B(n1080), .ZN(n1242) );
XOR2_X1 U956 ( .A(n1215), .B(n1243), .Z(n1080) );
XNOR2_X1 U957 ( .A(KEYINPUT11), .B(n1244), .ZN(n1243) );
XOR2_X1 U958 ( .A(G128), .B(G146), .Z(n1215) );
XOR2_X1 U959 ( .A(n1245), .B(n1246), .Z(n1136) );
NAND2_X1 U960 ( .A1(KEYINPUT17), .A2(n1118), .ZN(n1245) );
XOR2_X1 U961 ( .A(n1128), .B(n1247), .Z(n1241) );
XOR2_X1 U962 ( .A(n1248), .B(KEYINPUT10), .Z(n1247) );
NAND2_X1 U963 ( .A1(KEYINPUT49), .A2(n1129), .ZN(n1248) );
XNOR2_X1 U964 ( .A(n1249), .B(n1250), .ZN(n1129) );
XOR2_X1 U965 ( .A(G140), .B(G110), .Z(n1250) );
NAND2_X1 U966 ( .A1(G227), .A2(n1026), .ZN(n1249) );
XNOR2_X1 U967 ( .A(n1081), .B(KEYINPUT28), .ZN(n1128) );
XNOR2_X1 U968 ( .A(n1251), .B(n1252), .ZN(n1081) );
XOR2_X1 U969 ( .A(KEYINPUT14), .B(G137), .Z(n1252) );
XOR2_X1 U970 ( .A(n1179), .B(n1253), .Z(n1251) );
INV_X1 U971 ( .A(G134), .ZN(n1179) );
NAND2_X1 U972 ( .A1(KEYINPUT3), .A2(G469), .ZN(n1239) );
INV_X1 U973 ( .A(n1202), .ZN(n1166) );
NAND2_X1 U974 ( .A1(n1033), .A2(n1254), .ZN(n1202) );
NAND4_X1 U975 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1255), .ZN(n1254) );
INV_X1 U976 ( .A(G898), .ZN(n1255) );
NAND3_X1 U977 ( .A1(n1194), .A2(n1026), .A3(G952), .ZN(n1033) );
NAND2_X1 U978 ( .A1(G237), .A2(G234), .ZN(n1194) );
INV_X1 U979 ( .A(n1029), .ZN(n1174) );
NOR2_X1 U980 ( .A1(n1049), .A2(n1050), .ZN(n1029) );
AND2_X1 U981 ( .A1(G214), .A2(n1256), .ZN(n1050) );
INV_X1 U982 ( .A(n1184), .ZN(n1049) );
NAND3_X1 U983 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1184) );
INV_X1 U984 ( .A(n1065), .ZN(n1259) );
NOR2_X1 U985 ( .A1(n1068), .A2(n1067), .ZN(n1065) );
OR2_X1 U986 ( .A1(n1067), .A2(KEYINPUT55), .ZN(n1258) );
NAND3_X1 U987 ( .A1(n1067), .A2(n1068), .A3(KEYINPUT55), .ZN(n1257) );
NAND2_X1 U988 ( .A1(n1138), .A2(n1211), .ZN(n1068) );
XNOR2_X1 U989 ( .A(n1260), .B(n1261), .ZN(n1138) );
XOR2_X1 U990 ( .A(n1262), .B(n1095), .Z(n1261) );
XNOR2_X1 U991 ( .A(n1263), .B(G122), .ZN(n1095) );
NAND2_X1 U992 ( .A1(n1264), .A2(KEYINPUT47), .ZN(n1263) );
XOR2_X1 U993 ( .A(n1205), .B(KEYINPUT15), .Z(n1264) );
INV_X1 U994 ( .A(n1123), .ZN(n1262) );
XOR2_X1 U995 ( .A(n1265), .B(G128), .Z(n1123) );
NAND2_X1 U996 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U997 ( .A1(n1244), .A2(n1268), .ZN(n1267) );
XOR2_X1 U998 ( .A(KEYINPUT9), .B(n1269), .Z(n1266) );
NOR2_X1 U999 ( .A1(n1244), .A2(n1268), .ZN(n1269) );
XNOR2_X1 U1000 ( .A(G143), .B(KEYINPUT22), .ZN(n1244) );
XOR2_X1 U1001 ( .A(n1270), .B(n1271), .Z(n1260) );
AND2_X1 U1002 ( .A1(n1026), .A2(G224), .ZN(n1271) );
XOR2_X1 U1003 ( .A(n1272), .B(G125), .Z(n1270) );
NAND3_X1 U1004 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1272) );
NAND2_X1 U1005 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U1006 ( .A1(n1278), .A2(n1279), .ZN(n1274) );
INV_X1 U1007 ( .A(KEYINPUT63), .ZN(n1279) );
NAND2_X1 U1008 ( .A1(n1097), .A2(n1280), .ZN(n1278) );
XOR2_X1 U1009 ( .A(KEYINPUT37), .B(n1098), .Z(n1280) );
INV_X1 U1010 ( .A(n1276), .ZN(n1098) );
NAND2_X1 U1011 ( .A1(KEYINPUT63), .A2(n1281), .ZN(n1273) );
NAND2_X1 U1012 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
OR3_X1 U1013 ( .A1(n1276), .A2(n1277), .A3(KEYINPUT37), .ZN(n1283) );
INV_X1 U1014 ( .A(n1097), .ZN(n1277) );
XOR2_X1 U1015 ( .A(n1284), .B(n1232), .Z(n1097) );
INV_X1 U1016 ( .A(n1285), .ZN(n1232) );
XOR2_X1 U1017 ( .A(n1286), .B(G113), .Z(n1284) );
NAND2_X1 U1018 ( .A1(KEYINPUT30), .A2(n1218), .ZN(n1286) );
XOR2_X1 U1019 ( .A(G119), .B(KEYINPUT48), .Z(n1218) );
NAND2_X1 U1020 ( .A1(KEYINPUT37), .A2(n1276), .ZN(n1282) );
XNOR2_X1 U1021 ( .A(n1246), .B(n1287), .ZN(n1276) );
XNOR2_X1 U1022 ( .A(n1288), .B(KEYINPUT35), .ZN(n1287) );
NAND2_X1 U1023 ( .A1(KEYINPUT18), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1024 ( .A(KEYINPUT51), .B(G104), .Z(n1289) );
XOR2_X1 U1025 ( .A(G101), .B(n1290), .Z(n1246) );
XOR2_X1 U1026 ( .A(KEYINPUT21), .B(G107), .Z(n1290) );
INV_X1 U1027 ( .A(n1140), .ZN(n1067) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1256), .ZN(n1140) );
NAND2_X1 U1029 ( .A1(n1291), .A2(n1211), .ZN(n1256) );
INV_X1 U1030 ( .A(G237), .ZN(n1291) );
INV_X1 U1031 ( .A(n1058), .ZN(n1021) );
NAND2_X1 U1032 ( .A1(n1175), .A2(n1176), .ZN(n1058) );
XOR2_X1 U1033 ( .A(n1292), .B(G475), .Z(n1176) );
NAND2_X1 U1034 ( .A1(n1211), .A2(n1114), .ZN(n1292) );
NAND2_X1 U1035 ( .A1(n1293), .A2(n1294), .ZN(n1114) );
NAND3_X1 U1036 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
XOR2_X1 U1037 ( .A(n1118), .B(n1298), .Z(n1295) );
INV_X1 U1038 ( .A(G104), .ZN(n1118) );
NAND2_X1 U1039 ( .A1(n1299), .A2(n1300), .ZN(n1293) );
NAND2_X1 U1040 ( .A1(n1297), .A2(n1296), .ZN(n1300) );
NAND2_X1 U1041 ( .A1(n1301), .A2(n1302), .ZN(n1296) );
XOR2_X1 U1042 ( .A(n1303), .B(n1253), .Z(n1301) );
XOR2_X1 U1043 ( .A(KEYINPUT25), .B(n1304), .Z(n1297) );
AND2_X1 U1044 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XNOR2_X1 U1045 ( .A(n1303), .B(n1253), .ZN(n1306) );
XOR2_X1 U1046 ( .A(G131), .B(KEYINPUT36), .Z(n1253) );
NAND3_X1 U1047 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1303) );
NAND2_X1 U1048 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
OR4_X1 U1049 ( .A1(n1310), .A2(KEYINPUT19), .A3(n1311), .A4(n1312), .ZN(n1308) );
INV_X1 U1050 ( .A(KEYINPUT5), .ZN(n1311) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1235), .ZN(n1310) );
NAND2_X1 U1052 ( .A1(n1312), .A2(n1313), .ZN(n1307) );
NAND3_X1 U1053 ( .A1(n1235), .A2(n1314), .A3(G214), .ZN(n1313) );
INV_X1 U1054 ( .A(KEYINPUT19), .ZN(n1314) );
NOR2_X1 U1055 ( .A1(G953), .A2(G237), .ZN(n1235) );
XNOR2_X1 U1056 ( .A(G143), .B(KEYINPUT24), .ZN(n1312) );
XOR2_X1 U1057 ( .A(n1302), .B(KEYINPUT45), .Z(n1305) );
XOR2_X1 U1058 ( .A(n1268), .B(n1079), .Z(n1302) );
XOR2_X1 U1059 ( .A(G125), .B(G140), .Z(n1079) );
INV_X1 U1060 ( .A(G146), .ZN(n1268) );
XOR2_X1 U1061 ( .A(n1298), .B(G104), .Z(n1299) );
NAND2_X1 U1062 ( .A1(n1315), .A2(KEYINPUT26), .ZN(n1298) );
XOR2_X1 U1063 ( .A(n1316), .B(G122), .Z(n1315) );
INV_X1 U1064 ( .A(G113), .ZN(n1316) );
INV_X1 U1065 ( .A(G902), .ZN(n1211) );
XOR2_X1 U1066 ( .A(n1317), .B(G478), .Z(n1175) );
OR2_X1 U1067 ( .A1(n1107), .A2(G902), .ZN(n1317) );
XNOR2_X1 U1068 ( .A(n1318), .B(n1319), .ZN(n1107) );
XOR2_X1 U1069 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1070 ( .A(G107), .B(n1322), .Z(n1321) );
AND3_X1 U1071 ( .A1(G234), .A2(n1026), .A3(G217), .ZN(n1322) );
INV_X1 U1072 ( .A(G953), .ZN(n1026) );
XOR2_X1 U1073 ( .A(G143), .B(G134), .Z(n1320) );
XOR2_X1 U1074 ( .A(n1285), .B(n1323), .Z(n1318) );
XNOR2_X1 U1075 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1076 ( .A1(G128), .A2(KEYINPUT52), .ZN(n1325) );
NAND2_X1 U1077 ( .A1(KEYINPUT42), .A2(n1326), .ZN(n1324) );
INV_X1 U1078 ( .A(G122), .ZN(n1326) );
XNOR2_X1 U1079 ( .A(G116), .B(KEYINPUT0), .ZN(n1285) );
INV_X1 U1080 ( .A(G110), .ZN(n1205) );
endmodule


