//Key = 0101100010111111110100000001011000111100001100010111101010011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319;

XNOR2_X1 U729 ( .A(G107), .B(n1003), .ZN(G9) );
NOR2_X1 U730 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1006), .A2(n1007), .A3(G953), .A4(n1008), .ZN(n1005) );
NOR2_X1 U732 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U733 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR3_X1 U734 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR3_X1 U735 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR2_X1 U736 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U739 ( .A1(n1025), .A2(n1026), .ZN(n1017) );
NOR2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U741 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
XOR2_X1 U742 ( .A(KEYINPUT52), .B(n1031), .Z(n1030) );
NOR2_X1 U743 ( .A1(n1032), .A2(n1033), .ZN(n1014) );
NOR3_X1 U744 ( .A1(n1020), .A2(n1034), .A3(n1026), .ZN(n1033) );
NOR4_X1 U745 ( .A1(n1035), .A2(n1016), .A3(n1026), .A4(n1020), .ZN(n1011) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1006) );
XNOR2_X1 U748 ( .A(n1040), .B(KEYINPUT60), .ZN(n1038) );
NOR3_X1 U749 ( .A1(n1008), .A2(G953), .A3(G952), .ZN(n1004) );
AND4_X1 U750 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1008) );
NOR3_X1 U751 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NAND3_X1 U753 ( .A1(n1024), .A2(n1050), .A3(n1029), .ZN(n1045) );
NOR3_X1 U754 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U756 ( .A(n1056), .B(KEYINPUT50), .Z(n1055) );
INV_X1 U757 ( .A(G472), .ZN(n1054) );
NOR2_X1 U758 ( .A1(G472), .A2(n1056), .ZN(n1052) );
XNOR2_X1 U759 ( .A(G469), .B(n1057), .ZN(n1051) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(G72) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
XOR2_X1 U762 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U763 ( .A(KEYINPUT19), .B(n1064), .Z(n1063) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(n1062) );
NAND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1058) );
NAND2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U767 ( .A(n1039), .B(KEYINPUT6), .ZN(n1069) );
NAND2_X1 U768 ( .A1(G953), .A2(n1071), .ZN(n1067) );
NAND2_X1 U769 ( .A1(n1072), .A2(G900), .ZN(n1071) );
XNOR2_X1 U770 ( .A(G227), .B(KEYINPUT54), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(G69) );
NAND2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U773 ( .A1(G953), .A2(n1077), .ZN(n1076) );
NAND3_X1 U774 ( .A1(G953), .A2(n1078), .A3(n1079), .ZN(n1073) );
XNOR2_X1 U775 ( .A(n1075), .B(KEYINPUT22), .ZN(n1079) );
XNOR2_X1 U776 ( .A(n1080), .B(n1081), .ZN(n1075) );
NOR3_X1 U777 ( .A1(n1082), .A2(KEYINPUT31), .A3(n1083), .ZN(n1081) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(n1082) );
XNOR2_X1 U779 ( .A(n1086), .B(KEYINPUT10), .ZN(n1085) );
NAND2_X1 U780 ( .A1(KEYINPUT1), .A2(n1087), .ZN(n1086) );
NAND2_X1 U781 ( .A1(n1070), .A2(n1088), .ZN(n1080) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1078) );
NOR2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XOR2_X1 U785 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND3_X1 U786 ( .A1(n1095), .A2(n1096), .A3(KEYINPUT17), .ZN(n1093) );
NOR2_X1 U787 ( .A1(n1091), .A2(n1097), .ZN(G63) );
XOR2_X1 U788 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U789 ( .A1(n1095), .A2(G478), .ZN(n1098) );
NOR3_X1 U790 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(G60) );
AND2_X1 U791 ( .A1(KEYINPUT36), .A2(n1091), .ZN(n1102) );
NOR3_X1 U792 ( .A1(KEYINPUT36), .A2(n1070), .A3(n1103), .ZN(n1101) );
INV_X1 U793 ( .A(G952), .ZN(n1103) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1100) );
NAND2_X1 U795 ( .A1(n1095), .A2(G475), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(G6) );
NAND2_X1 U797 ( .A1(G104), .A2(n1108), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1109), .B(KEYINPUT25), .Z(n1106) );
OR2_X1 U799 ( .A1(n1108), .A2(G104), .ZN(n1109) );
NOR3_X1 U800 ( .A1(n1091), .A2(n1110), .A3(n1111), .ZN(G57) );
NOR2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NOR2_X1 U805 ( .A1(G101), .A2(n1120), .ZN(n1110) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U807 ( .A1(n1118), .A2(n1116), .ZN(n1122) );
XNOR2_X1 U808 ( .A(n1123), .B(n1119), .ZN(n1116) );
XNOR2_X1 U809 ( .A(KEYINPUT40), .B(KEYINPUT37), .ZN(n1123) );
INV_X1 U810 ( .A(n1117), .ZN(n1118) );
NOR2_X1 U811 ( .A1(n1119), .A2(n1117), .ZN(n1121) );
XNOR2_X1 U812 ( .A(n1124), .B(n1125), .ZN(n1119) );
NAND2_X1 U813 ( .A1(n1095), .A2(G472), .ZN(n1124) );
NOR2_X1 U814 ( .A1(n1091), .A2(n1126), .ZN(G54) );
XOR2_X1 U815 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1129) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1127) );
XNOR2_X1 U819 ( .A(KEYINPUT34), .B(n1135), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1133) );
NOR2_X1 U821 ( .A1(KEYINPUT39), .A2(n1138), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1095), .A2(G469), .ZN(n1136) );
NOR2_X1 U823 ( .A1(n1091), .A2(n1139), .ZN(G51) );
XOR2_X1 U824 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U825 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U827 ( .A(KEYINPUT62), .B(n1146), .Z(n1144) );
AND2_X1 U828 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
XOR2_X1 U829 ( .A(n1147), .B(n1148), .Z(n1140) );
NAND2_X1 U830 ( .A1(n1095), .A2(n1048), .ZN(n1147) );
AND2_X1 U831 ( .A1(G902), .A2(n1149), .ZN(n1095) );
NAND2_X1 U832 ( .A1(n1039), .A2(n1040), .ZN(n1149) );
AND2_X1 U833 ( .A1(n1150), .A2(n1089), .ZN(n1040) );
AND4_X1 U834 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1089) );
NAND4_X1 U835 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1151) );
XOR2_X1 U836 ( .A(KEYINPUT26), .B(n1022), .Z(n1157) );
XNOR2_X1 U837 ( .A(n1090), .B(KEYINPUT30), .ZN(n1150) );
AND4_X1 U838 ( .A1(n1108), .A2(n1159), .A3(n1160), .A4(n1003), .ZN(n1090) );
NAND3_X1 U839 ( .A1(n1032), .A2(n1036), .A3(n1161), .ZN(n1003) );
NAND3_X1 U840 ( .A1(n1032), .A2(n1037), .A3(n1161), .ZN(n1108) );
AND4_X1 U841 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1039) );
NOR4_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NOR3_X1 U843 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
AND3_X1 U844 ( .A1(n1173), .A2(n1037), .A3(n1022), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1164) );
NOR2_X1 U846 ( .A1(n1070), .A2(G952), .ZN(n1091) );
XOR2_X1 U847 ( .A(n1176), .B(n1177), .Z(G48) );
NAND2_X1 U848 ( .A1(KEYINPUT29), .A2(G146), .ZN(n1177) );
NAND3_X1 U849 ( .A1(n1173), .A2(n1037), .A3(n1178), .ZN(n1176) );
XOR2_X1 U850 ( .A(n1171), .B(KEYINPUT35), .Z(n1178) );
INV_X1 U851 ( .A(n1170), .ZN(n1173) );
XOR2_X1 U852 ( .A(G143), .B(n1167), .Z(G45) );
AND3_X1 U853 ( .A1(n1179), .A2(n1022), .A3(n1180), .ZN(n1167) );
XNOR2_X1 U854 ( .A(n1166), .B(n1181), .ZN(G42) );
NAND2_X1 U855 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1181) );
AND3_X1 U856 ( .A1(n1182), .A2(n1028), .A3(n1183), .ZN(n1166) );
XOR2_X1 U857 ( .A(G137), .B(n1175), .Z(G39) );
NOR3_X1 U858 ( .A1(n1170), .A2(n1026), .A3(n1013), .ZN(n1175) );
XOR2_X1 U859 ( .A(G134), .B(n1174), .Z(G36) );
AND3_X1 U860 ( .A1(n1179), .A2(n1036), .A3(n1182), .ZN(n1174) );
XOR2_X1 U861 ( .A(G131), .B(n1184), .Z(G33) );
NOR2_X1 U862 ( .A1(KEYINPUT21), .A2(n1162), .ZN(n1184) );
NAND3_X1 U863 ( .A1(n1179), .A2(n1037), .A3(n1182), .ZN(n1162) );
INV_X1 U864 ( .A(n1026), .ZN(n1182) );
NAND2_X1 U865 ( .A1(n1185), .A2(n1024), .ZN(n1026) );
INV_X1 U866 ( .A(n1023), .ZN(n1185) );
AND3_X1 U867 ( .A1(n1028), .A2(n1186), .A3(n1187), .ZN(n1179) );
XOR2_X1 U868 ( .A(G128), .B(n1188), .Z(G30) );
NOR3_X1 U869 ( .A1(n1189), .A2(n1172), .A3(n1170), .ZN(n1188) );
NAND3_X1 U870 ( .A1(n1028), .A2(n1186), .A3(n1034), .ZN(n1170) );
XOR2_X1 U871 ( .A(KEYINPUT42), .B(n1022), .Z(n1189) );
XOR2_X1 U872 ( .A(n1113), .B(n1159), .Z(G3) );
NAND3_X1 U873 ( .A1(n1187), .A2(n1161), .A3(n1190), .ZN(n1159) );
XOR2_X1 U874 ( .A(n1191), .B(n1163), .Z(G27) );
NAND3_X1 U875 ( .A1(n1183), .A2(n1022), .A3(n1156), .ZN(n1163) );
AND4_X1 U876 ( .A1(n1192), .A2(n1037), .A3(n1047), .A4(n1186), .ZN(n1183) );
NAND2_X1 U877 ( .A1(n1010), .A2(n1193), .ZN(n1186) );
NAND3_X1 U878 ( .A1(G902), .A2(n1194), .A3(n1060), .ZN(n1193) );
NOR2_X1 U879 ( .A1(n1070), .A2(G900), .ZN(n1060) );
XOR2_X1 U880 ( .A(n1195), .B(G122), .Z(G24) );
NAND2_X1 U881 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND4_X1 U882 ( .A1(n1156), .A2(n1180), .A3(n1198), .A4(n1199), .ZN(n1197) );
NOR3_X1 U883 ( .A1(n1016), .A2(n1022), .A3(n1200), .ZN(n1198) );
INV_X1 U884 ( .A(n1032), .ZN(n1016) );
INV_X1 U885 ( .A(n1020), .ZN(n1156) );
OR2_X1 U886 ( .A1(n1152), .A2(n1199), .ZN(n1196) );
INV_X1 U887 ( .A(KEYINPUT3), .ZN(n1199) );
NAND3_X1 U888 ( .A1(n1180), .A2(n1032), .A3(n1201), .ZN(n1152) );
NOR2_X1 U889 ( .A1(n1202), .A2(n1047), .ZN(n1032) );
XOR2_X1 U890 ( .A(G119), .B(n1203), .Z(G21) );
AND2_X1 U891 ( .A1(n1201), .A2(n1155), .ZN(n1203) );
AND2_X1 U892 ( .A1(n1190), .A2(n1034), .ZN(n1155) );
AND2_X1 U893 ( .A1(n1047), .A2(n1202), .ZN(n1034) );
INV_X1 U894 ( .A(n1192), .ZN(n1202) );
XNOR2_X1 U895 ( .A(G116), .B(n1153), .ZN(G18) );
NAND3_X1 U896 ( .A1(n1187), .A2(n1036), .A3(n1201), .ZN(n1153) );
INV_X1 U897 ( .A(n1172), .ZN(n1036) );
NAND2_X1 U898 ( .A1(n1204), .A2(n1205), .ZN(n1172) );
XOR2_X1 U899 ( .A(n1206), .B(n1154), .Z(G15) );
NAND3_X1 U900 ( .A1(n1187), .A2(n1037), .A3(n1201), .ZN(n1154) );
NOR3_X1 U901 ( .A1(n1171), .A2(n1200), .A3(n1020), .ZN(n1201) );
NAND2_X1 U902 ( .A1(n1207), .A2(n1031), .ZN(n1020) );
XNOR2_X1 U903 ( .A(n1208), .B(KEYINPUT41), .ZN(n1031) );
XOR2_X1 U904 ( .A(n1029), .B(KEYINPUT32), .Z(n1207) );
INV_X1 U905 ( .A(n1158), .ZN(n1200) );
NAND2_X1 U906 ( .A1(n1209), .A2(n1210), .ZN(n1037) );
NAND3_X1 U907 ( .A1(n1211), .A2(n1041), .A3(n1212), .ZN(n1210) );
INV_X1 U908 ( .A(KEYINPUT28), .ZN(n1212) );
NAND2_X1 U909 ( .A1(KEYINPUT28), .A2(n1180), .ZN(n1209) );
AND2_X1 U910 ( .A1(n1211), .A2(n1204), .ZN(n1180) );
INV_X1 U911 ( .A(n1041), .ZN(n1204) );
XNOR2_X1 U912 ( .A(n1042), .B(KEYINPUT5), .ZN(n1211) );
NOR2_X1 U913 ( .A1(n1047), .A2(n1192), .ZN(n1187) );
XOR2_X1 U914 ( .A(n1213), .B(n1160), .Z(G12) );
NAND4_X1 U915 ( .A1(n1190), .A2(n1161), .A3(n1192), .A4(n1047), .ZN(n1160) );
XNOR2_X1 U916 ( .A(n1214), .B(n1096), .ZN(n1047) );
AND2_X1 U917 ( .A1(G217), .A2(n1215), .ZN(n1096) );
NAND2_X1 U918 ( .A1(n1094), .A2(n1216), .ZN(n1214) );
XOR2_X1 U919 ( .A(n1217), .B(n1218), .Z(n1094) );
XOR2_X1 U920 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U921 ( .A1(G137), .A2(KEYINPUT9), .ZN(n1220) );
NOR2_X1 U922 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
INV_X1 U923 ( .A(G221), .ZN(n1221) );
XOR2_X1 U924 ( .A(n1223), .B(n1224), .Z(n1217) );
NOR3_X1 U925 ( .A1(KEYINPUT44), .A2(n1225), .A3(n1226), .ZN(n1224) );
NOR3_X1 U926 ( .A1(G110), .A2(n1227), .A3(n1228), .ZN(n1226) );
NOR2_X1 U927 ( .A1(n1229), .A2(n1213), .ZN(n1225) );
NOR2_X1 U928 ( .A1(n1227), .A2(n1228), .ZN(n1229) );
XNOR2_X1 U929 ( .A(n1230), .B(KEYINPUT55), .ZN(n1228) );
NAND2_X1 U930 ( .A1(G128), .A2(n1231), .ZN(n1230) );
AND2_X1 U931 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
XOR2_X1 U932 ( .A(KEYINPUT53), .B(G119), .Z(n1232) );
NAND2_X1 U933 ( .A1(n1234), .A2(n1235), .ZN(n1223) );
NAND2_X1 U934 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XOR2_X1 U935 ( .A(KEYINPUT43), .B(n1238), .Z(n1234) );
NOR2_X1 U936 ( .A1(n1239), .A2(n1237), .ZN(n1238) );
XOR2_X1 U937 ( .A(n1064), .B(KEYINPUT13), .Z(n1237) );
INV_X1 U938 ( .A(n1240), .ZN(n1064) );
XOR2_X1 U939 ( .A(n1236), .B(KEYINPUT24), .Z(n1239) );
XOR2_X1 U940 ( .A(n1241), .B(KEYINPUT48), .Z(n1236) );
XOR2_X1 U941 ( .A(n1056), .B(G472), .Z(n1192) );
NAND2_X1 U942 ( .A1(n1242), .A2(n1216), .ZN(n1056) );
XOR2_X1 U943 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U944 ( .A(KEYINPUT18), .B(G101), .Z(n1244) );
XOR2_X1 U945 ( .A(n1125), .B(n1117), .Z(n1243) );
NAND2_X1 U946 ( .A1(n1245), .A2(G210), .ZN(n1117) );
XNOR2_X1 U947 ( .A(n1246), .B(n1247), .ZN(n1125) );
XOR2_X1 U948 ( .A(n1206), .B(n1248), .Z(n1247) );
XOR2_X1 U949 ( .A(n1249), .B(n1250), .Z(n1246) );
AND3_X1 U950 ( .A1(n1022), .A2(n1158), .A3(n1028), .ZN(n1161) );
AND2_X1 U951 ( .A1(n1208), .A2(n1029), .ZN(n1028) );
NAND2_X1 U952 ( .A1(G221), .A2(n1215), .ZN(n1029) );
NAND2_X1 U953 ( .A1(G234), .A2(n1251), .ZN(n1215) );
XNOR2_X1 U954 ( .A(G469), .B(n1252), .ZN(n1208) );
NOR2_X1 U955 ( .A1(KEYINPUT2), .A2(n1253), .ZN(n1252) );
XOR2_X1 U956 ( .A(n1057), .B(KEYINPUT15), .Z(n1253) );
NAND2_X1 U957 ( .A1(n1216), .A2(n1254), .ZN(n1057) );
XNOR2_X1 U958 ( .A(n1138), .B(n1255), .ZN(n1254) );
XOR2_X1 U959 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U960 ( .A1(KEYINPUT46), .A2(n1135), .ZN(n1257) );
NAND2_X1 U961 ( .A1(G227), .A2(n1070), .ZN(n1135) );
NOR2_X1 U962 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
XOR2_X1 U963 ( .A(n1260), .B(KEYINPUT8), .Z(n1259) );
NAND2_X1 U964 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U965 ( .A(KEYINPUT4), .B(n1263), .Z(n1262) );
INV_X1 U966 ( .A(n1131), .ZN(n1263) );
NOR2_X1 U967 ( .A1(n1131), .A2(n1261), .ZN(n1258) );
XOR2_X1 U968 ( .A(n1264), .B(n1132), .Z(n1261) );
INV_X1 U969 ( .A(n1065), .ZN(n1132) );
XOR2_X1 U970 ( .A(n1233), .B(n1265), .Z(n1065) );
XOR2_X1 U971 ( .A(G146), .B(G143), .Z(n1265) );
NAND2_X1 U972 ( .A1(KEYINPUT12), .A2(n1130), .ZN(n1264) );
XNOR2_X1 U973 ( .A(n1266), .B(n1267), .ZN(n1130) );
XOR2_X1 U974 ( .A(n1113), .B(KEYINPUT63), .Z(n1266) );
INV_X1 U975 ( .A(G101), .ZN(n1113) );
XOR2_X1 U976 ( .A(n1249), .B(KEYINPUT56), .Z(n1131) );
XNOR2_X1 U977 ( .A(n1066), .B(KEYINPUT47), .ZN(n1249) );
XOR2_X1 U978 ( .A(G131), .B(n1268), .Z(n1066) );
XOR2_X1 U979 ( .A(G137), .B(G134), .Z(n1268) );
XOR2_X1 U980 ( .A(G140), .B(n1213), .Z(n1138) );
NAND2_X1 U981 ( .A1(n1010), .A2(n1269), .ZN(n1158) );
NAND3_X1 U982 ( .A1(G902), .A2(n1194), .A3(n1083), .ZN(n1269) );
NOR2_X1 U983 ( .A1(n1070), .A2(G898), .ZN(n1083) );
NAND3_X1 U984 ( .A1(n1194), .A2(n1070), .A3(G952), .ZN(n1010) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1194) );
INV_X1 U986 ( .A(n1171), .ZN(n1022) );
NAND2_X1 U987 ( .A1(n1023), .A2(n1024), .ZN(n1171) );
NAND2_X1 U988 ( .A1(G214), .A2(n1270), .ZN(n1024) );
NAND2_X1 U989 ( .A1(n1271), .A2(n1272), .ZN(n1023) );
NAND2_X1 U990 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U991 ( .A1(KEYINPUT51), .A2(n1049), .ZN(n1273) );
NAND2_X1 U992 ( .A1(n1275), .A2(KEYINPUT51), .ZN(n1271) );
INV_X1 U993 ( .A(n1050), .ZN(n1275) );
NAND2_X1 U994 ( .A1(n1048), .A2(n1049), .ZN(n1050) );
NAND2_X1 U995 ( .A1(n1276), .A2(n1216), .ZN(n1049) );
XOR2_X1 U996 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U997 ( .A(n1148), .B(n1145), .Z(n1278) );
XOR2_X1 U998 ( .A(n1248), .B(G125), .Z(n1145) );
NAND2_X1 U999 ( .A1(n1279), .A2(n1280), .ZN(n1248) );
NAND2_X1 U1000 ( .A1(n1281), .A2(n1233), .ZN(n1280) );
XOR2_X1 U1001 ( .A(n1282), .B(KEYINPUT61), .Z(n1279) );
OR2_X1 U1002 ( .A1(n1281), .A2(n1233), .ZN(n1282) );
INV_X1 U1003 ( .A(G128), .ZN(n1233) );
XNOR2_X1 U1004 ( .A(n1283), .B(G143), .ZN(n1281) );
NAND2_X1 U1005 ( .A1(KEYINPUT11), .A2(n1241), .ZN(n1283) );
INV_X1 U1006 ( .A(G146), .ZN(n1241) );
XOR2_X1 U1007 ( .A(n1084), .B(n1087), .Z(n1148) );
XNOR2_X1 U1008 ( .A(G113), .B(n1284), .ZN(n1087) );
NOR2_X1 U1009 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
AND3_X1 U1010 ( .A1(KEYINPUT23), .A2(n1231), .A3(G116), .ZN(n1286) );
INV_X1 U1011 ( .A(G119), .ZN(n1231) );
NOR2_X1 U1012 ( .A1(KEYINPUT23), .A2(n1250), .ZN(n1285) );
XOR2_X1 U1013 ( .A(G116), .B(G119), .Z(n1250) );
XOR2_X1 U1014 ( .A(n1287), .B(n1288), .Z(n1084) );
XOR2_X1 U1015 ( .A(n1289), .B(n1267), .Z(n1288) );
XOR2_X1 U1016 ( .A(G104), .B(G107), .Z(n1267) );
NOR2_X1 U1017 ( .A1(G101), .A2(KEYINPUT0), .ZN(n1289) );
XOR2_X1 U1018 ( .A(n1213), .B(G122), .Z(n1287) );
XNOR2_X1 U1019 ( .A(n1146), .B(KEYINPUT14), .ZN(n1277) );
NOR2_X1 U1020 ( .A1(n1077), .A2(G953), .ZN(n1146) );
INV_X1 U1021 ( .A(G224), .ZN(n1077) );
INV_X1 U1022 ( .A(n1274), .ZN(n1048) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1270), .ZN(n1274) );
NAND2_X1 U1024 ( .A1(n1290), .A2(n1251), .ZN(n1270) );
INV_X1 U1025 ( .A(G237), .ZN(n1290) );
INV_X1 U1026 ( .A(n1013), .ZN(n1190) );
NAND2_X1 U1027 ( .A1(n1291), .A2(n1205), .ZN(n1013) );
XNOR2_X1 U1028 ( .A(n1042), .B(KEYINPUT59), .ZN(n1205) );
XOR2_X1 U1029 ( .A(n1292), .B(G475), .Z(n1042) );
NAND2_X1 U1030 ( .A1(n1105), .A2(n1216), .ZN(n1292) );
XOR2_X1 U1031 ( .A(n1293), .B(n1294), .Z(n1105) );
XOR2_X1 U1032 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1033 ( .A(G131), .B(G104), .Z(n1296) );
XOR2_X1 U1034 ( .A(KEYINPUT45), .B(G146), .Z(n1295) );
XOR2_X1 U1035 ( .A(n1297), .B(n1298), .Z(n1293) );
XOR2_X1 U1036 ( .A(n1299), .B(n1240), .Z(n1298) );
XOR2_X1 U1037 ( .A(n1191), .B(G140), .Z(n1240) );
INV_X1 U1038 ( .A(G125), .ZN(n1191) );
NAND2_X1 U1039 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U1040 ( .A1(G122), .A2(n1206), .ZN(n1301) );
XOR2_X1 U1041 ( .A(n1302), .B(KEYINPUT38), .Z(n1300) );
OR2_X1 U1042 ( .A1(n1206), .A2(G122), .ZN(n1302) );
INV_X1 U1043 ( .A(G113), .ZN(n1206) );
XOR2_X1 U1044 ( .A(n1303), .B(n1304), .Z(n1297) );
NOR2_X1 U1045 ( .A1(KEYINPUT58), .A2(n1305), .ZN(n1304) );
INV_X1 U1046 ( .A(G143), .ZN(n1305) );
NAND2_X1 U1047 ( .A1(n1245), .A2(G214), .ZN(n1303) );
NOR2_X1 U1048 ( .A1(G953), .A2(G237), .ZN(n1245) );
XOR2_X1 U1049 ( .A(n1041), .B(KEYINPUT33), .Z(n1291) );
XOR2_X1 U1050 ( .A(n1306), .B(G478), .Z(n1041) );
NAND2_X1 U1051 ( .A1(n1099), .A2(n1216), .ZN(n1306) );
XOR2_X1 U1052 ( .A(n1251), .B(KEYINPUT20), .Z(n1216) );
INV_X1 U1053 ( .A(G902), .ZN(n1251) );
XOR2_X1 U1054 ( .A(n1307), .B(n1308), .Z(n1099) );
NOR2_X1 U1055 ( .A1(n1309), .A2(n1222), .ZN(n1308) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1070), .ZN(n1222) );
INV_X1 U1057 ( .A(G953), .ZN(n1070) );
INV_X1 U1058 ( .A(G217), .ZN(n1309) );
NAND2_X1 U1059 ( .A1(n1310), .A2(n1311), .ZN(n1307) );
NAND2_X1 U1060 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1061 ( .A(KEYINPUT16), .B(n1314), .Z(n1310) );
NOR2_X1 U1062 ( .A1(n1313), .A2(n1312), .ZN(n1314) );
XOR2_X1 U1063 ( .A(G107), .B(n1315), .Z(n1312) );
NOR2_X1 U1064 ( .A1(KEYINPUT7), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1065 ( .A(G116), .B(G122), .ZN(n1316) );
XNOR2_X1 U1066 ( .A(n1317), .B(n1318), .ZN(n1313) );
NOR2_X1 U1067 ( .A1(G134), .A2(KEYINPUT57), .ZN(n1318) );
XOR2_X1 U1068 ( .A(n1319), .B(G143), .Z(n1317) );
NAND2_X1 U1069 ( .A1(KEYINPUT27), .A2(G128), .ZN(n1319) );
INV_X1 U1070 ( .A(G110), .ZN(n1213) );
endmodule


