//Key = 0010001111011010111011111011110100001100100111101010000100111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363;

XNOR2_X1 U757 ( .A(G107), .B(n1047), .ZN(G9) );
NOR2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
XOR2_X1 U760 ( .A(KEYINPUT29), .B(n1053), .Z(n1052) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR4_X1 U762 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1056) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U767 ( .A(n1068), .B(KEYINPUT34), .Z(n1066) );
NOR2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1060) );
NOR4_X1 U769 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1069) );
NOR2_X1 U770 ( .A1(n1075), .A2(n1068), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1063), .ZN(n1073) );
NOR2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1077) );
INV_X1 U775 ( .A(KEYINPUT30), .ZN(n1082) );
NOR4_X1 U776 ( .A1(KEYINPUT30), .A2(n1081), .A3(n1083), .A4(n1084), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1068), .B(KEYINPUT39), .Z(n1081) );
NOR4_X1 U778 ( .A1(n1085), .A2(n1068), .A3(n1086), .A4(n1070), .ZN(n1054) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1057), .ZN(n1087) );
OR2_X1 U781 ( .A1(n1058), .A2(n1063), .ZN(n1085) );
NAND3_X1 U782 ( .A1(n1090), .A2(n1091), .A3(G952), .ZN(n1050) );
NOR3_X1 U783 ( .A1(n1092), .A2(G953), .A3(n1093), .ZN(n1048) );
INV_X1 U784 ( .A(n1090), .ZN(n1093) );
NAND4_X1 U785 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1090) );
NOR4_X1 U786 ( .A1(n1098), .A2(n1099), .A3(n1070), .A4(n1057), .ZN(n1097) );
INV_X1 U787 ( .A(n1083), .ZN(n1099) );
INV_X1 U788 ( .A(n1080), .ZN(n1098) );
XOR2_X1 U789 ( .A(n1100), .B(n1101), .Z(n1096) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U791 ( .A1(KEYINPUT1), .A2(n1104), .ZN(n1103) );
NAND2_X1 U792 ( .A1(KEYINPUT40), .A2(n1105), .ZN(n1102) );
XOR2_X1 U793 ( .A(n1089), .B(KEYINPUT61), .Z(n1095) );
XNOR2_X1 U794 ( .A(n1106), .B(n1107), .ZN(n1094) );
NAND2_X1 U795 ( .A1(KEYINPUT6), .A2(G469), .ZN(n1106) );
XOR2_X1 U796 ( .A(KEYINPUT15), .B(G952), .Z(n1092) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1091), .ZN(n1109) );
AND2_X1 U799 ( .A1(G227), .A2(G900), .ZN(n1110) );
NAND2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U801 ( .A1(n1113), .A2(n1091), .ZN(n1112) );
XNOR2_X1 U802 ( .A(n1114), .B(n1115), .ZN(n1113) );
NAND3_X1 U803 ( .A1(G900), .A2(n1115), .A3(G953), .ZN(n1111) );
XNOR2_X1 U804 ( .A(n1116), .B(n1117), .ZN(n1115) );
XNOR2_X1 U805 ( .A(n1118), .B(KEYINPUT57), .ZN(n1117) );
NAND2_X1 U806 ( .A1(n1119), .A2(KEYINPUT45), .ZN(n1118) );
XNOR2_X1 U807 ( .A(G125), .B(n1120), .ZN(n1119) );
XOR2_X1 U808 ( .A(KEYINPUT5), .B(G140), .Z(n1120) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1116) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(G69) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1091), .ZN(n1124) );
AND2_X1 U812 ( .A1(G224), .A2(G898), .ZN(n1125) );
NAND2_X1 U813 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
NAND3_X1 U814 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
INV_X1 U815 ( .A(n1131), .ZN(n1129) );
OR2_X1 U816 ( .A1(n1130), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U817 ( .A(n1132), .B(n1133), .ZN(n1128) );
XNOR2_X1 U818 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U819 ( .A(n1136), .B(KEYINPUT22), .Z(n1132) );
NAND2_X1 U820 ( .A1(n1091), .A2(n1137), .ZN(n1130) );
NAND2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U823 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND3_X1 U824 ( .A1(n1144), .A2(n1145), .A3(KEYINPUT36), .ZN(n1142) );
NOR2_X1 U825 ( .A1(n1140), .A2(n1146), .ZN(G63) );
XNOR2_X1 U826 ( .A(n1147), .B(n1148), .ZN(n1146) );
AND2_X1 U827 ( .A1(G478), .A2(n1144), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1149), .ZN(G60) );
XOR2_X1 U829 ( .A(n1150), .B(n1151), .Z(n1149) );
AND2_X1 U830 ( .A1(G475), .A2(n1144), .ZN(n1150) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(G6) );
NOR2_X1 U832 ( .A1(n1140), .A2(n1154), .ZN(G57) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U834 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U835 ( .A1(KEYINPUT37), .A2(n1159), .ZN(n1155) );
XOR2_X1 U836 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U837 ( .A(n1162), .B(n1163), .ZN(n1161) );
XNOR2_X1 U838 ( .A(n1164), .B(n1165), .ZN(n1160) );
NAND2_X1 U839 ( .A1(KEYINPUT48), .A2(n1166), .ZN(n1164) );
NAND2_X1 U840 ( .A1(n1144), .A2(G472), .ZN(n1166) );
INV_X1 U841 ( .A(n1167), .ZN(n1144) );
NOR2_X1 U842 ( .A1(n1140), .A2(n1168), .ZN(G54) );
XOR2_X1 U843 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U844 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U845 ( .A1(KEYINPUT27), .A2(n1173), .ZN(n1171) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1169) );
NAND3_X1 U847 ( .A1(G469), .A2(n1051), .A3(n1176), .ZN(n1175) );
XOR2_X1 U848 ( .A(n1177), .B(KEYINPUT2), .Z(n1176) );
NOR2_X1 U849 ( .A1(n1140), .A2(n1178), .ZN(G51) );
XOR2_X1 U850 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U851 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U852 ( .A1(n1104), .A2(n1167), .ZN(n1182) );
NAND2_X1 U853 ( .A1(G902), .A2(n1051), .ZN(n1167) );
NAND3_X1 U854 ( .A1(n1114), .A2(n1138), .A3(n1183), .ZN(n1051) );
XNOR2_X1 U855 ( .A(n1139), .B(KEYINPUT20), .ZN(n1183) );
AND4_X1 U856 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1139) );
NAND4_X1 U857 ( .A1(n1188), .A2(n1189), .A3(n1088), .A4(n1190), .ZN(n1184) );
AND2_X1 U858 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
OR2_X1 U859 ( .A1(n1071), .A2(KEYINPUT19), .ZN(n1189) );
NAND2_X1 U860 ( .A1(KEYINPUT19), .A2(n1193), .ZN(n1188) );
NAND2_X1 U861 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
AND4_X1 U862 ( .A1(n1153), .A2(n1196), .A3(n1197), .A4(n1047), .ZN(n1138) );
NAND3_X1 U863 ( .A1(n1089), .A2(n1192), .A3(n1198), .ZN(n1047) );
NAND3_X1 U864 ( .A1(n1089), .A2(n1198), .A3(n1199), .ZN(n1153) );
AND4_X1 U865 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1114) );
AND3_X1 U866 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NAND2_X1 U867 ( .A1(n1207), .A2(n1208), .ZN(n1202) );
NAND2_X1 U868 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
XOR2_X1 U870 ( .A(KEYINPUT35), .B(n1194), .Z(n1212) );
INV_X1 U871 ( .A(n1063), .ZN(n1194) );
NAND3_X1 U872 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1200) );
NAND2_X1 U873 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NOR2_X1 U875 ( .A1(KEYINPUT32), .A2(n1220), .ZN(n1181) );
XOR2_X1 U876 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U877 ( .A(n1165), .B(n1223), .ZN(n1221) );
NOR2_X1 U878 ( .A1(n1091), .A2(G952), .ZN(n1140) );
XOR2_X1 U879 ( .A(n1201), .B(n1224), .Z(G48) );
NAND2_X1 U880 ( .A1(G146), .A2(n1225), .ZN(n1224) );
XOR2_X1 U881 ( .A(KEYINPUT54), .B(KEYINPUT44), .Z(n1225) );
NAND3_X1 U882 ( .A1(n1218), .A2(n1226), .A3(n1199), .ZN(n1201) );
XOR2_X1 U883 ( .A(n1227), .B(n1228), .Z(G45) );
NAND2_X1 U884 ( .A1(n1229), .A2(n1207), .ZN(n1228) );
INV_X1 U885 ( .A(n1195), .ZN(n1207) );
XOR2_X1 U886 ( .A(n1210), .B(KEYINPUT50), .Z(n1229) );
NAND3_X1 U887 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1210) );
INV_X1 U888 ( .A(n1233), .ZN(n1230) );
XOR2_X1 U889 ( .A(G140), .B(n1234), .Z(G42) );
NOR3_X1 U890 ( .A1(n1235), .A2(n1068), .A3(n1217), .ZN(n1234) );
XOR2_X1 U891 ( .A(KEYINPUT23), .B(n1213), .Z(n1235) );
XNOR2_X1 U892 ( .A(G137), .B(n1236), .ZN(G39) );
NOR2_X1 U893 ( .A1(KEYINPUT56), .A2(n1237), .ZN(n1236) );
NOR4_X1 U894 ( .A1(n1238), .A2(n1070), .A3(n1068), .A4(n1239), .ZN(n1237) );
XOR2_X1 U895 ( .A(n1075), .B(KEYINPUT52), .Z(n1238) );
XNOR2_X1 U896 ( .A(G134), .B(n1205), .ZN(G36) );
NAND2_X1 U897 ( .A1(n1064), .A2(n1232), .ZN(n1205) );
AND2_X1 U898 ( .A1(n1215), .A2(n1192), .ZN(n1064) );
NAND2_X1 U899 ( .A1(n1240), .A2(n1241), .ZN(G33) );
OR2_X1 U900 ( .A1(n1204), .A2(G131), .ZN(n1241) );
XOR2_X1 U901 ( .A(n1242), .B(KEYINPUT10), .Z(n1240) );
NAND2_X1 U902 ( .A1(G131), .A2(n1204), .ZN(n1242) );
NAND3_X1 U903 ( .A1(n1232), .A2(n1215), .A3(n1199), .ZN(n1204) );
INV_X1 U904 ( .A(n1068), .ZN(n1215) );
NAND2_X1 U905 ( .A1(n1243), .A2(n1080), .ZN(n1068) );
AND3_X1 U906 ( .A1(n1213), .A2(n1244), .A3(n1088), .ZN(n1232) );
INV_X1 U907 ( .A(n1075), .ZN(n1213) );
NAND2_X1 U908 ( .A1(n1245), .A2(n1246), .ZN(G30) );
NAND2_X1 U909 ( .A1(n1247), .A2(n1206), .ZN(n1246) );
NAND2_X1 U910 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U911 ( .A1(KEYINPUT11), .A2(n1250), .ZN(n1249) );
INV_X1 U912 ( .A(KEYINPUT24), .ZN(n1250) );
NAND3_X1 U913 ( .A1(n1251), .A2(n1252), .A3(KEYINPUT24), .ZN(n1245) );
OR2_X1 U914 ( .A1(G128), .A2(KEYINPUT11), .ZN(n1252) );
NAND2_X1 U915 ( .A1(KEYINPUT11), .A2(n1253), .ZN(n1251) );
OR2_X1 U916 ( .A1(n1206), .A2(G128), .ZN(n1253) );
NAND3_X1 U917 ( .A1(n1192), .A2(n1226), .A3(n1218), .ZN(n1206) );
INV_X1 U918 ( .A(n1239), .ZN(n1218) );
NAND3_X1 U919 ( .A1(n1057), .A2(n1244), .A3(n1059), .ZN(n1239) );
XOR2_X1 U920 ( .A(G101), .B(n1254), .Z(G3) );
NOR2_X1 U921 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
AND2_X1 U922 ( .A1(KEYINPUT26), .A2(n1196), .ZN(n1256) );
NOR2_X1 U923 ( .A1(KEYINPUT59), .A2(n1196), .ZN(n1255) );
NAND4_X1 U924 ( .A1(n1088), .A2(n1219), .A3(n1226), .A4(n1191), .ZN(n1196) );
NAND2_X1 U925 ( .A1(n1257), .A2(n1258), .ZN(G27) );
OR2_X1 U926 ( .A1(G125), .A2(KEYINPUT58), .ZN(n1258) );
XOR2_X1 U927 ( .A(n1259), .B(n1260), .Z(n1257) );
AND2_X1 U928 ( .A1(n1211), .A2(n1071), .ZN(n1260) );
INV_X1 U929 ( .A(n1217), .ZN(n1211) );
NAND4_X1 U930 ( .A1(n1261), .A2(n1199), .A3(n1059), .A4(n1244), .ZN(n1217) );
NAND2_X1 U931 ( .A1(n1058), .A2(n1262), .ZN(n1244) );
NAND4_X1 U932 ( .A1(G902), .A2(G953), .A3(n1263), .A4(n1264), .ZN(n1262) );
INV_X1 U933 ( .A(G900), .ZN(n1264) );
NAND2_X1 U934 ( .A1(KEYINPUT58), .A2(G125), .ZN(n1259) );
XNOR2_X1 U935 ( .A(G122), .B(n1185), .ZN(G24) );
NAND3_X1 U936 ( .A1(n1089), .A2(n1265), .A3(n1266), .ZN(n1185) );
NOR3_X1 U937 ( .A1(n1057), .A2(n1267), .A3(n1233), .ZN(n1266) );
XOR2_X1 U938 ( .A(n1268), .B(n1186), .Z(G21) );
NAND4_X1 U939 ( .A1(n1265), .A2(n1219), .A3(n1059), .A4(n1057), .ZN(n1186) );
INV_X1 U940 ( .A(n1261), .ZN(n1057) );
XNOR2_X1 U941 ( .A(G116), .B(n1269), .ZN(G18) );
NAND2_X1 U942 ( .A1(n1270), .A2(n1192), .ZN(n1269) );
NOR2_X1 U943 ( .A1(n1231), .A2(n1233), .ZN(n1192) );
XOR2_X1 U944 ( .A(n1187), .B(n1271), .Z(G15) );
NAND2_X1 U945 ( .A1(KEYINPUT8), .A2(G113), .ZN(n1271) );
NAND2_X1 U946 ( .A1(n1270), .A2(n1199), .ZN(n1187) );
INV_X1 U947 ( .A(n1067), .ZN(n1199) );
NAND2_X1 U948 ( .A1(n1233), .A2(n1231), .ZN(n1067) );
INV_X1 U949 ( .A(n1267), .ZN(n1231) );
AND2_X1 U950 ( .A1(n1265), .A2(n1088), .ZN(n1270) );
NOR2_X1 U951 ( .A1(n1059), .A2(n1261), .ZN(n1088) );
AND2_X1 U952 ( .A1(n1071), .A2(n1191), .ZN(n1265) );
NOR2_X1 U953 ( .A1(n1063), .A2(n1195), .ZN(n1071) );
NAND2_X1 U954 ( .A1(n1272), .A2(n1083), .ZN(n1063) );
NAND2_X1 U955 ( .A1(n1273), .A2(n1274), .ZN(G12) );
NAND2_X1 U956 ( .A1(G110), .A2(n1197), .ZN(n1274) );
XOR2_X1 U957 ( .A(KEYINPUT16), .B(n1275), .Z(n1273) );
NOR2_X1 U958 ( .A1(G110), .A2(n1197), .ZN(n1275) );
NAND3_X1 U959 ( .A1(n1198), .A2(n1059), .A3(n1219), .ZN(n1197) );
INV_X1 U960 ( .A(n1070), .ZN(n1219) );
NAND2_X1 U961 ( .A1(n1233), .A2(n1267), .ZN(n1070) );
XOR2_X1 U962 ( .A(n1276), .B(G475), .Z(n1267) );
OR2_X1 U963 ( .A1(n1151), .A2(G902), .ZN(n1276) );
XNOR2_X1 U964 ( .A(n1277), .B(n1278), .ZN(n1151) );
XNOR2_X1 U965 ( .A(n1279), .B(n1280), .ZN(n1278) );
XOR2_X1 U966 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U967 ( .A1(n1283), .A2(G214), .ZN(n1281) );
XOR2_X1 U968 ( .A(n1284), .B(n1285), .Z(n1277) );
XOR2_X1 U969 ( .A(KEYINPUT41), .B(G131), .Z(n1285) );
XOR2_X1 U970 ( .A(n1286), .B(n1287), .Z(n1284) );
NOR2_X1 U971 ( .A1(G140), .A2(KEYINPUT38), .ZN(n1287) );
NAND3_X1 U972 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1286) );
NAND2_X1 U973 ( .A1(KEYINPUT4), .A2(n1291), .ZN(n1290) );
OR3_X1 U974 ( .A1(n1291), .A2(KEYINPUT4), .A3(n1152), .ZN(n1289) );
NAND2_X1 U975 ( .A1(n1292), .A2(n1152), .ZN(n1288) );
INV_X1 U976 ( .A(G104), .ZN(n1152) );
NAND2_X1 U977 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
INV_X1 U978 ( .A(KEYINPUT4), .ZN(n1294) );
XOR2_X1 U979 ( .A(KEYINPUT46), .B(n1291), .Z(n1293) );
XOR2_X1 U980 ( .A(G113), .B(n1295), .Z(n1291) );
XOR2_X1 U981 ( .A(n1296), .B(G478), .Z(n1233) );
NAND2_X1 U982 ( .A1(n1297), .A2(n1147), .ZN(n1296) );
XNOR2_X1 U983 ( .A(n1298), .B(n1299), .ZN(n1147) );
XOR2_X1 U984 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U985 ( .A(n1302), .B(n1303), .Z(n1301) );
AND3_X1 U986 ( .A1(G217), .A2(n1091), .A3(G234), .ZN(n1303) );
NAND2_X1 U987 ( .A1(n1304), .A2(KEYINPUT17), .ZN(n1302) );
XOR2_X1 U988 ( .A(n1248), .B(n1305), .Z(n1304) );
XOR2_X1 U989 ( .A(G143), .B(G134), .Z(n1305) );
XNOR2_X1 U990 ( .A(G107), .B(n1306), .ZN(n1298) );
XOR2_X1 U991 ( .A(KEYINPUT51), .B(G116), .Z(n1306) );
XOR2_X1 U992 ( .A(n1177), .B(KEYINPUT49), .Z(n1297) );
INV_X1 U993 ( .A(n1089), .ZN(n1059) );
XOR2_X1 U994 ( .A(n1307), .B(n1145), .Z(n1089) );
AND2_X1 U995 ( .A1(G217), .A2(n1308), .ZN(n1145) );
NAND2_X1 U996 ( .A1(n1143), .A2(n1177), .ZN(n1307) );
XOR2_X1 U997 ( .A(n1309), .B(n1310), .Z(n1143) );
XOR2_X1 U998 ( .A(G137), .B(n1311), .Z(n1310) );
AND3_X1 U999 ( .A1(G221), .A2(n1091), .A3(G234), .ZN(n1311) );
NAND2_X1 U1000 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1001 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1002 ( .A(n1316), .B(KEYINPUT62), .Z(n1312) );
NAND2_X1 U1003 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1004 ( .A(KEYINPUT31), .B(n1315), .Z(n1318) );
XNOR2_X1 U1005 ( .A(n1319), .B(n1282), .ZN(n1315) );
XOR2_X1 U1006 ( .A(G125), .B(KEYINPUT25), .Z(n1282) );
XOR2_X1 U1007 ( .A(G146), .B(n1174), .Z(n1319) );
XOR2_X1 U1008 ( .A(n1314), .B(KEYINPUT28), .Z(n1317) );
XNOR2_X1 U1009 ( .A(G110), .B(n1320), .ZN(n1314) );
XOR2_X1 U1010 ( .A(G128), .B(G119), .Z(n1320) );
AND3_X1 U1011 ( .A1(n1261), .A2(n1191), .A3(n1226), .ZN(n1198) );
NOR2_X1 U1012 ( .A1(n1195), .A2(n1075), .ZN(n1226) );
NAND2_X1 U1013 ( .A1(n1084), .A2(n1083), .ZN(n1075) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1308), .ZN(n1083) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1177), .ZN(n1308) );
INV_X1 U1016 ( .A(n1272), .ZN(n1084) );
XOR2_X1 U1017 ( .A(n1107), .B(G469), .Z(n1272) );
NAND2_X1 U1018 ( .A1(n1321), .A2(n1177), .ZN(n1107) );
XNOR2_X1 U1019 ( .A(n1173), .B(n1322), .ZN(n1321) );
NOR2_X1 U1020 ( .A1(KEYINPUT63), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1021 ( .A(n1324), .B(n1172), .Z(n1323) );
XOR2_X1 U1022 ( .A(n1325), .B(G110), .Z(n1172) );
NAND2_X1 U1023 ( .A1(n1326), .A2(n1091), .ZN(n1325) );
XOR2_X1 U1024 ( .A(KEYINPUT47), .B(G227), .Z(n1326) );
NAND2_X1 U1025 ( .A1(KEYINPUT14), .A2(n1174), .ZN(n1324) );
INV_X1 U1026 ( .A(G140), .ZN(n1174) );
XNOR2_X1 U1027 ( .A(n1327), .B(n1328), .ZN(n1173) );
XNOR2_X1 U1028 ( .A(n1121), .B(n1329), .ZN(n1328) );
XOR2_X1 U1029 ( .A(n1330), .B(G128), .Z(n1121) );
NAND2_X1 U1030 ( .A1(KEYINPUT43), .A2(n1279), .ZN(n1330) );
XOR2_X1 U1031 ( .A(n1162), .B(G101), .Z(n1327) );
NAND2_X1 U1032 ( .A1(n1079), .A2(n1080), .ZN(n1195) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1331), .ZN(n1080) );
INV_X1 U1034 ( .A(n1243), .ZN(n1079) );
XOR2_X1 U1035 ( .A(n1100), .B(n1105), .Z(n1243) );
INV_X1 U1036 ( .A(n1104), .ZN(n1105) );
NAND2_X1 U1037 ( .A1(G210), .A2(n1331), .ZN(n1104) );
NAND2_X1 U1038 ( .A1(n1332), .A2(n1177), .ZN(n1331) );
INV_X1 U1039 ( .A(G237), .ZN(n1332) );
NAND2_X1 U1040 ( .A1(n1333), .A2(n1177), .ZN(n1100) );
XOR2_X1 U1041 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1042 ( .A(n1222), .B(n1179), .Z(n1335) );
XOR2_X1 U1043 ( .A(n1336), .B(n1136), .Z(n1179) );
NAND2_X1 U1044 ( .A1(n1337), .A2(n1338), .ZN(n1136) );
NAND2_X1 U1045 ( .A1(G110), .A2(n1295), .ZN(n1338) );
XOR2_X1 U1046 ( .A(n1339), .B(KEYINPUT42), .Z(n1337) );
OR2_X1 U1047 ( .A1(n1295), .A2(G110), .ZN(n1339) );
INV_X1 U1048 ( .A(n1300), .ZN(n1295) );
XNOR2_X1 U1049 ( .A(G122), .B(KEYINPUT18), .ZN(n1300) );
NAND2_X1 U1050 ( .A1(n1340), .A2(n1341), .ZN(n1336) );
NAND2_X1 U1051 ( .A1(n1135), .A2(n1134), .ZN(n1341) );
XOR2_X1 U1052 ( .A(KEYINPUT55), .B(n1342), .Z(n1340) );
NOR2_X1 U1053 ( .A1(n1135), .A2(n1134), .ZN(n1342) );
XOR2_X1 U1054 ( .A(G101), .B(n1343), .Z(n1134) );
NOR2_X1 U1055 ( .A1(KEYINPUT13), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1056 ( .A(KEYINPUT21), .B(n1329), .Z(n1344) );
XOR2_X1 U1057 ( .A(G107), .B(G104), .Z(n1329) );
XOR2_X1 U1058 ( .A(n1345), .B(n1346), .Z(n1135) );
NAND2_X1 U1059 ( .A1(KEYINPUT9), .A2(n1268), .ZN(n1345) );
XOR2_X1 U1060 ( .A(G125), .B(KEYINPUT33), .Z(n1222) );
XOR2_X1 U1061 ( .A(n1347), .B(n1223), .Z(n1334) );
AND2_X1 U1062 ( .A1(G224), .A2(n1091), .ZN(n1223) );
NAND2_X1 U1063 ( .A1(KEYINPUT60), .A2(n1165), .ZN(n1347) );
NAND2_X1 U1064 ( .A1(n1058), .A2(n1348), .ZN(n1191) );
NAND3_X1 U1065 ( .A1(n1131), .A2(n1263), .A3(G902), .ZN(n1348) );
NOR2_X1 U1066 ( .A1(n1091), .A2(G898), .ZN(n1131) );
NAND3_X1 U1067 ( .A1(n1263), .A2(n1091), .A3(G952), .ZN(n1058) );
INV_X1 U1068 ( .A(G953), .ZN(n1091) );
NAND2_X1 U1069 ( .A1(G237), .A2(G234), .ZN(n1263) );
XOR2_X1 U1070 ( .A(n1349), .B(G472), .Z(n1261) );
NAND2_X1 U1071 ( .A1(n1350), .A2(n1177), .ZN(n1349) );
INV_X1 U1072 ( .A(G902), .ZN(n1177) );
XOR2_X1 U1073 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1074 ( .A1(n1158), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1075 ( .A(KEYINPUT3), .B(n1157), .Z(n1353) );
NOR2_X1 U1076 ( .A1(n1354), .A2(G101), .ZN(n1157) );
AND2_X1 U1077 ( .A1(n1283), .A2(G210), .ZN(n1354) );
AND3_X1 U1078 ( .A1(G210), .A2(G101), .A3(n1283), .ZN(n1158) );
NOR2_X1 U1079 ( .A1(G953), .A2(G237), .ZN(n1283) );
NOR2_X1 U1080 ( .A1(n1355), .A2(n1356), .ZN(n1351) );
XOR2_X1 U1081 ( .A(n1357), .B(KEYINPUT7), .Z(n1356) );
NAND3_X1 U1082 ( .A1(n1358), .A2(n1359), .A3(n1163), .ZN(n1357) );
NOR2_X1 U1083 ( .A1(n1360), .A2(n1163), .ZN(n1355) );
XOR2_X1 U1084 ( .A(n1346), .B(n1361), .Z(n1163) );
NOR2_X1 U1085 ( .A1(KEYINPUT0), .A2(n1268), .ZN(n1361) );
INV_X1 U1086 ( .A(G119), .ZN(n1268) );
XOR2_X1 U1087 ( .A(G113), .B(G116), .Z(n1346) );
AND2_X1 U1088 ( .A1(n1359), .A2(n1358), .ZN(n1360) );
OR2_X1 U1089 ( .A1(n1165), .A2(n1162), .ZN(n1358) );
NAND2_X1 U1090 ( .A1(n1362), .A2(n1165), .ZN(n1359) );
XNOR2_X1 U1091 ( .A(n1248), .B(n1279), .ZN(n1165) );
XNOR2_X1 U1092 ( .A(n1227), .B(G146), .ZN(n1279) );
INV_X1 U1093 ( .A(G143), .ZN(n1227) );
INV_X1 U1094 ( .A(G128), .ZN(n1248) );
XOR2_X1 U1095 ( .A(n1162), .B(KEYINPUT53), .Z(n1362) );
XNOR2_X1 U1096 ( .A(n1122), .B(KEYINPUT12), .ZN(n1162) );
XOR2_X1 U1097 ( .A(G131), .B(n1363), .Z(n1122) );
XOR2_X1 U1098 ( .A(G137), .B(G134), .Z(n1363) );
endmodule


