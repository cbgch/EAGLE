//Key = 1000111101110000010001011000000001010000000101011110001100011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333;

XOR2_X1 U738 ( .A(n1018), .B(n1019), .Z(G9) );
NAND2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR3_X1 U741 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR3_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
NOR3_X1 U743 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
AND4_X1 U745 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(KEYINPUT54), .ZN(n1031) );
OR2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
INV_X1 U750 ( .A(n1046), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
AND2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
XOR2_X1 U753 ( .A(KEYINPUT62), .B(n1051), .Z(n1030) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1034), .ZN(n1051) );
XNOR2_X1 U755 ( .A(n1020), .B(KEYINPUT27), .ZN(n1052) );
NAND3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1024) );
NAND3_X1 U757 ( .A1(n1037), .A2(n1056), .A3(n1057), .ZN(n1055) );
INV_X1 U758 ( .A(n1034), .ZN(n1057) );
NAND4_X1 U759 ( .A1(KEYINPUT54), .A2(n1058), .A3(n1046), .A4(n1036), .ZN(n1034) );
NAND2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1028), .A2(n1061), .ZN(n1060) );
NOR3_X1 U762 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U763 ( .A(n1053), .ZN(n1062) );
NAND4_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1053) );
NOR4_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XNOR2_X1 U766 ( .A(G469), .B(n1071), .ZN(n1070) );
XOR2_X1 U767 ( .A(G478), .B(n1072), .Z(n1069) );
NOR2_X1 U768 ( .A1(KEYINPUT15), .A2(n1073), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1074), .B(KEYINPUT26), .Z(n1073) );
XOR2_X1 U770 ( .A(n1061), .B(KEYINPUT43), .Z(n1067) );
NOR3_X1 U771 ( .A1(n1050), .A2(n1075), .A3(n1028), .ZN(n1065) );
INV_X1 U772 ( .A(n1076), .ZN(n1028) );
XOR2_X1 U773 ( .A(G472), .B(n1077), .Z(n1063) );
NOR2_X1 U774 ( .A1(n1078), .A2(KEYINPUT51), .ZN(n1077) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U776 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U778 ( .A1(G953), .A2(n1085), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1083) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U781 ( .A(G140), .B(G131), .Z(n1089) );
XOR2_X1 U782 ( .A(KEYINPUT21), .B(KEYINPUT10), .Z(n1088) );
XOR2_X1 U783 ( .A(n1090), .B(n1091), .Z(n1086) );
XOR2_X1 U784 ( .A(G125), .B(n1092), .Z(n1091) );
NAND2_X1 U785 ( .A1(n1054), .A2(n1093), .ZN(n1081) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XNOR2_X1 U787 ( .A(KEYINPUT33), .B(n1096), .ZN(n1095) );
NOR3_X1 U788 ( .A1(n1054), .A2(KEYINPUT34), .A3(n1097), .ZN(n1079) );
AND2_X1 U789 ( .A1(G227), .A2(G900), .ZN(n1097) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(G69) );
XOR2_X1 U791 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U792 ( .A1(n1102), .A2(n1054), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
NAND2_X1 U795 ( .A1(G953), .A2(n1104), .ZN(n1106) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(n1105) );
NAND2_X1 U797 ( .A1(n1054), .A2(n1109), .ZN(n1098) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XNOR2_X1 U799 ( .A(n1112), .B(n1113), .ZN(n1111) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1110), .A2(n1116), .ZN(G63) );
NOR3_X1 U802 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR3_X1 U804 ( .A1(n1122), .A2(KEYINPUT18), .A3(n1123), .ZN(n1120) );
INV_X1 U805 ( .A(n1026), .ZN(n1123) );
NOR4_X1 U806 ( .A1(n1124), .A2(n1115), .A3(KEYINPUT18), .A4(n1122), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1110), .A2(n1125), .ZN(G60) );
XNOR2_X1 U808 ( .A(n1126), .B(n1127), .ZN(n1125) );
AND2_X1 U809 ( .A1(G475), .A2(n1128), .ZN(n1127) );
XNOR2_X1 U810 ( .A(G104), .B(n1129), .ZN(G6) );
NOR2_X1 U811 ( .A1(n1110), .A2(n1130), .ZN(G57) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U814 ( .A1(KEYINPUT60), .A2(n1090), .ZN(n1133) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1131) );
AND2_X1 U816 ( .A1(G472), .A2(n1128), .ZN(n1136) );
XNOR2_X1 U817 ( .A(n1137), .B(KEYINPUT16), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1110), .A2(n1138), .ZN(G54) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U820 ( .A(KEYINPUT20), .B(n1141), .Z(n1140) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
AND2_X1 U822 ( .A1(n1143), .A2(n1142), .ZN(n1139) );
XNOR2_X1 U823 ( .A(n1144), .B(n1145), .ZN(n1142) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U825 ( .A1(KEYINPUT1), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U826 ( .A(n1149), .B(n1150), .ZN(n1144) );
NAND2_X1 U827 ( .A1(n1128), .A2(G469), .ZN(n1143) );
INV_X1 U828 ( .A(n1115), .ZN(n1128) );
NOR2_X1 U829 ( .A1(n1110), .A2(n1151), .ZN(G51) );
XOR2_X1 U830 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U831 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U832 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U833 ( .A1(n1158), .A2(n1115), .ZN(n1157) );
NAND2_X1 U834 ( .A1(G902), .A2(n1026), .ZN(n1115) );
NAND3_X1 U835 ( .A1(n1159), .A2(n1096), .A3(n1094), .ZN(n1026) );
AND4_X1 U836 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1094) );
AND4_X1 U837 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NAND3_X1 U838 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1162) );
XOR2_X1 U839 ( .A(n1171), .B(KEYINPUT40), .Z(n1168) );
INV_X1 U840 ( .A(n1109), .ZN(n1159) );
NAND4_X1 U841 ( .A1(n1129), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1109) );
NOR4_X1 U842 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
INV_X1 U843 ( .A(n1179), .ZN(n1178) );
NAND2_X1 U844 ( .A1(n1020), .A2(n1180), .ZN(n1173) );
NAND2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND3_X1 U846 ( .A1(n1046), .A2(n1183), .A3(n1184), .ZN(n1182) );
XOR2_X1 U847 ( .A(KEYINPUT3), .B(n1048), .Z(n1183) );
NAND2_X1 U848 ( .A1(n1185), .A2(n1042), .ZN(n1181) );
NAND2_X1 U849 ( .A1(n1169), .A2(n1021), .ZN(n1129) );
AND3_X1 U850 ( .A1(n1046), .A2(n1048), .A3(n1184), .ZN(n1021) );
NAND2_X1 U851 ( .A1(KEYINPUT0), .A2(G125), .ZN(n1156) );
NOR2_X1 U852 ( .A1(n1054), .A2(G952), .ZN(n1110) );
XOR2_X1 U853 ( .A(n1186), .B(n1187), .Z(G48) );
NAND3_X1 U854 ( .A1(n1188), .A2(n1171), .A3(n1189), .ZN(n1187) );
XOR2_X1 U855 ( .A(KEYINPUT37), .B(n1048), .Z(n1188) );
XNOR2_X1 U856 ( .A(G143), .B(n1160), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1170), .A2(n1042), .A3(n1190), .A4(n1191), .ZN(n1160) );
XOR2_X1 U858 ( .A(n1161), .B(n1192), .Z(G42) );
NAND2_X1 U859 ( .A1(KEYINPUT47), .A2(G140), .ZN(n1192) );
NAND3_X1 U860 ( .A1(n1169), .A2(n1043), .A3(n1193), .ZN(n1161) );
XNOR2_X1 U861 ( .A(G137), .B(n1167), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1193), .A2(n1171), .A3(n1037), .ZN(n1167) );
NAND2_X1 U863 ( .A1(n1194), .A2(n1195), .ZN(G36) );
OR2_X1 U864 ( .A1(n1096), .A2(G134), .ZN(n1195) );
XOR2_X1 U865 ( .A(n1196), .B(KEYINPUT56), .Z(n1194) );
NAND2_X1 U866 ( .A1(G134), .A2(n1096), .ZN(n1196) );
NAND3_X1 U867 ( .A1(n1042), .A2(n1020), .A3(n1193), .ZN(n1096) );
NAND2_X1 U868 ( .A1(n1197), .A2(n1198), .ZN(G33) );
NAND2_X1 U869 ( .A1(G131), .A2(n1166), .ZN(n1198) );
XOR2_X1 U870 ( .A(n1199), .B(KEYINPUT19), .Z(n1197) );
OR2_X1 U871 ( .A1(n1166), .A2(G131), .ZN(n1199) );
NAND3_X1 U872 ( .A1(n1042), .A2(n1169), .A3(n1193), .ZN(n1166) );
AND4_X1 U873 ( .A1(n1061), .A2(n1048), .A3(n1200), .A4(n1076), .ZN(n1193) );
XOR2_X1 U874 ( .A(n1201), .B(n1165), .Z(G30) );
NAND3_X1 U875 ( .A1(n1020), .A2(n1171), .A3(n1170), .ZN(n1165) );
AND3_X1 U876 ( .A1(n1202), .A2(n1200), .A3(n1048), .ZN(n1170) );
XOR2_X1 U877 ( .A(n1177), .B(n1203), .Z(G3) );
XOR2_X1 U878 ( .A(KEYINPUT25), .B(G101), .Z(n1203) );
AND2_X1 U879 ( .A1(n1204), .A2(n1042), .ZN(n1177) );
XOR2_X1 U880 ( .A(n1205), .B(n1164), .Z(G27) );
NAND3_X1 U881 ( .A1(n1189), .A2(n1043), .A3(n1058), .ZN(n1164) );
AND3_X1 U882 ( .A1(n1202), .A2(n1200), .A3(n1169), .ZN(n1189) );
NAND2_X1 U883 ( .A1(n1206), .A2(n1207), .ZN(n1200) );
NAND2_X1 U884 ( .A1(n1208), .A2(n1085), .ZN(n1207) );
INV_X1 U885 ( .A(G900), .ZN(n1085) );
XNOR2_X1 U886 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U887 ( .A1(n1185), .A2(n1046), .A3(n1190), .A4(n1191), .ZN(n1172) );
XOR2_X1 U888 ( .A(n1209), .B(n1179), .Z(G21) );
NAND3_X1 U889 ( .A1(n1037), .A2(n1171), .A3(n1185), .ZN(n1179) );
NAND2_X1 U890 ( .A1(n1210), .A2(n1211), .ZN(n1171) );
NAND2_X1 U891 ( .A1(n1042), .A2(n1212), .ZN(n1211) );
NAND3_X1 U892 ( .A1(n1213), .A2(n1068), .A3(KEYINPUT63), .ZN(n1210) );
XNOR2_X1 U893 ( .A(G116), .B(n1214), .ZN(G18) );
NAND4_X1 U894 ( .A1(n1215), .A2(KEYINPUT17), .A3(n1185), .A4(n1042), .ZN(n1214) );
XNOR2_X1 U895 ( .A(n1020), .B(KEYINPUT23), .ZN(n1215) );
NOR2_X1 U896 ( .A1(n1191), .A2(n1216), .ZN(n1020) );
XOR2_X1 U897 ( .A(n1176), .B(n1217), .Z(G15) );
NOR2_X1 U898 ( .A1(KEYINPUT58), .A2(n1218), .ZN(n1217) );
AND3_X1 U899 ( .A1(n1042), .A2(n1169), .A3(n1185), .ZN(n1176) );
AND2_X1 U900 ( .A1(n1058), .A2(n1184), .ZN(n1185) );
INV_X1 U901 ( .A(n1041), .ZN(n1058) );
NAND2_X1 U902 ( .A1(n1049), .A2(n1219), .ZN(n1041) );
INV_X1 U903 ( .A(n1050), .ZN(n1219) );
INV_X1 U904 ( .A(n1033), .ZN(n1169) );
NAND2_X1 U905 ( .A1(n1216), .A2(n1191), .ZN(n1033) );
INV_X1 U906 ( .A(n1190), .ZN(n1216) );
NOR2_X1 U907 ( .A1(n1068), .A2(n1220), .ZN(n1042) );
NAND2_X1 U908 ( .A1(n1221), .A2(n1222), .ZN(G12) );
NAND2_X1 U909 ( .A1(n1175), .A2(n1148), .ZN(n1222) );
XOR2_X1 U910 ( .A(KEYINPUT61), .B(n1223), .Z(n1221) );
NOR2_X1 U911 ( .A1(n1175), .A2(n1148), .ZN(n1223) );
AND2_X1 U912 ( .A1(n1204), .A2(n1043), .ZN(n1175) );
NAND2_X1 U913 ( .A1(n1224), .A2(n1225), .ZN(n1043) );
NAND2_X1 U914 ( .A1(n1046), .A2(n1212), .ZN(n1225) );
INV_X1 U915 ( .A(KEYINPUT63), .ZN(n1212) );
NOR2_X1 U916 ( .A1(n1068), .A2(n1213), .ZN(n1046) );
NAND3_X1 U917 ( .A1(n1068), .A2(n1220), .A3(KEYINPUT63), .ZN(n1224) );
INV_X1 U918 ( .A(n1213), .ZN(n1220) );
XOR2_X1 U919 ( .A(n1078), .B(G472), .Z(n1213) );
AND2_X1 U920 ( .A1(n1226), .A2(n1227), .ZN(n1078) );
XNOR2_X1 U921 ( .A(n1134), .B(n1228), .ZN(n1226) );
XOR2_X1 U922 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U923 ( .A1(KEYINPUT55), .A2(n1137), .ZN(n1229) );
AND3_X1 U924 ( .A1(n1231), .A2(n1054), .A3(G210), .ZN(n1137) );
XNOR2_X1 U925 ( .A(n1232), .B(n1233), .ZN(n1134) );
XOR2_X1 U926 ( .A(G101), .B(n1234), .Z(n1233) );
XOR2_X1 U927 ( .A(KEYINPUT14), .B(G113), .Z(n1234) );
XOR2_X1 U928 ( .A(n1235), .B(n1236), .Z(n1232) );
NOR2_X1 U929 ( .A1(KEYINPUT8), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U930 ( .A(G116), .B(n1238), .ZN(n1237) );
NAND2_X1 U931 ( .A1(KEYINPUT5), .A2(n1209), .ZN(n1238) );
XNOR2_X1 U932 ( .A(n1239), .B(n1240), .ZN(n1068) );
NOR2_X1 U933 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U934 ( .A(KEYINPUT9), .B(G217), .Z(n1242) );
NAND2_X1 U935 ( .A1(n1112), .A2(n1227), .ZN(n1239) );
XNOR2_X1 U936 ( .A(n1243), .B(n1244), .ZN(n1112) );
XOR2_X1 U937 ( .A(G137), .B(n1245), .Z(n1244) );
NOR2_X1 U938 ( .A1(KEYINPUT36), .A2(n1246), .ZN(n1245) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U940 ( .A(G146), .B(G125), .Z(n1248) );
NOR2_X1 U941 ( .A1(G140), .A2(KEYINPUT28), .ZN(n1247) );
XOR2_X1 U942 ( .A(n1249), .B(n1250), .Z(n1243) );
NOR4_X1 U943 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
XNOR2_X1 U944 ( .A(KEYINPUT39), .B(KEYINPUT24), .ZN(n1252) );
XOR2_X1 U945 ( .A(n1054), .B(KEYINPUT49), .Z(n1251) );
NAND2_X1 U946 ( .A1(n1255), .A2(n1256), .ZN(n1249) );
OR2_X1 U947 ( .A1(n1257), .A2(G110), .ZN(n1256) );
XOR2_X1 U948 ( .A(n1258), .B(KEYINPUT30), .Z(n1255) );
NAND2_X1 U949 ( .A1(G110), .A2(n1257), .ZN(n1258) );
XNOR2_X1 U950 ( .A(n1209), .B(n1259), .ZN(n1257) );
XOR2_X1 U951 ( .A(KEYINPUT13), .B(G128), .Z(n1259) );
INV_X1 U952 ( .A(G119), .ZN(n1209) );
AND3_X1 U953 ( .A1(n1184), .A2(n1048), .A3(n1037), .ZN(n1204) );
NOR2_X1 U954 ( .A1(n1191), .A2(n1190), .ZN(n1037) );
XOR2_X1 U955 ( .A(n1260), .B(n1117), .Z(n1190) );
INV_X1 U956 ( .A(n1074), .ZN(n1117) );
NAND2_X1 U957 ( .A1(n1124), .A2(n1227), .ZN(n1074) );
INV_X1 U958 ( .A(n1121), .ZN(n1124) );
XOR2_X1 U959 ( .A(n1261), .B(n1262), .Z(n1121) );
XOR2_X1 U960 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U961 ( .A(n1018), .B(n1265), .Z(n1264) );
INV_X1 U962 ( .A(G107), .ZN(n1018) );
NAND2_X1 U963 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
NAND2_X1 U964 ( .A1(n1268), .A2(n1201), .ZN(n1267) );
XOR2_X1 U965 ( .A(KEYINPUT50), .B(n1269), .Z(n1268) );
NAND2_X1 U966 ( .A1(n1270), .A2(G128), .ZN(n1266) );
XOR2_X1 U967 ( .A(KEYINPUT12), .B(n1269), .Z(n1270) );
NOR3_X1 U968 ( .A1(n1114), .A2(G953), .A3(n1253), .ZN(n1269) );
INV_X1 U969 ( .A(G217), .ZN(n1114) );
XNOR2_X1 U970 ( .A(G116), .B(n1271), .ZN(n1261) );
XOR2_X1 U971 ( .A(G143), .B(G134), .Z(n1271) );
NAND2_X1 U972 ( .A1(KEYINPUT6), .A2(n1122), .ZN(n1260) );
INV_X1 U973 ( .A(G478), .ZN(n1122) );
NAND2_X1 U974 ( .A1(n1272), .A2(n1064), .ZN(n1191) );
NAND2_X1 U975 ( .A1(G475), .A2(n1273), .ZN(n1064) );
XOR2_X1 U976 ( .A(KEYINPUT7), .B(n1075), .Z(n1272) );
NOR2_X1 U977 ( .A1(n1273), .A2(G475), .ZN(n1075) );
NAND2_X1 U978 ( .A1(n1126), .A2(n1227), .ZN(n1273) );
XNOR2_X1 U979 ( .A(n1274), .B(n1275), .ZN(n1126) );
NOR2_X1 U980 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U981 ( .A(KEYINPUT53), .B(n1278), .Z(n1277) );
NOR2_X1 U982 ( .A1(n1186), .A2(n1279), .ZN(n1278) );
XOR2_X1 U983 ( .A(KEYINPUT31), .B(n1280), .Z(n1279) );
AND2_X1 U984 ( .A1(n1186), .A2(n1280), .ZN(n1276) );
XNOR2_X1 U985 ( .A(n1281), .B(G125), .ZN(n1280) );
NAND2_X1 U986 ( .A1(KEYINPUT4), .A2(n1282), .ZN(n1281) );
INV_X1 U987 ( .A(G140), .ZN(n1282) );
INV_X1 U988 ( .A(G146), .ZN(n1186) );
XOR2_X1 U989 ( .A(n1283), .B(n1284), .Z(n1274) );
NOR2_X1 U990 ( .A1(KEYINPUT52), .A2(n1285), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U992 ( .A(G143), .B(G131), .Z(n1287) );
NAND3_X1 U993 ( .A1(G214), .A2(n1054), .A3(n1288), .ZN(n1286) );
XOR2_X1 U994 ( .A(n1231), .B(KEYINPUT22), .Z(n1288) );
NAND2_X1 U995 ( .A1(n1289), .A2(n1290), .ZN(n1283) );
NAND2_X1 U996 ( .A1(G104), .A2(n1291), .ZN(n1290) );
XOR2_X1 U997 ( .A(KEYINPUT35), .B(n1292), .Z(n1289) );
NOR2_X1 U998 ( .A1(G104), .A2(n1291), .ZN(n1292) );
XOR2_X1 U999 ( .A(n1218), .B(n1293), .Z(n1291) );
NOR2_X1 U1000 ( .A1(KEYINPUT44), .A2(n1265), .ZN(n1293) );
INV_X1 U1001 ( .A(G113), .ZN(n1218) );
NOR2_X1 U1002 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U1003 ( .A1(n1254), .A2(n1241), .ZN(n1050) );
NOR2_X1 U1004 ( .A1(n1253), .A2(G902), .ZN(n1241) );
INV_X1 U1005 ( .A(G234), .ZN(n1253) );
INV_X1 U1006 ( .A(G221), .ZN(n1254) );
XNOR2_X1 U1007 ( .A(n1071), .B(n1294), .ZN(n1049) );
NOR2_X1 U1008 ( .A1(G469), .A2(KEYINPUT41), .ZN(n1294) );
NAND3_X1 U1009 ( .A1(n1295), .A2(n1296), .A3(n1227), .ZN(n1071) );
OR3_X1 U1010 ( .A1(n1297), .A2(n1298), .A3(KEYINPUT48), .ZN(n1296) );
NAND2_X1 U1011 ( .A1(n1299), .A2(KEYINPUT48), .ZN(n1295) );
XOR2_X1 U1012 ( .A(n1297), .B(n1298), .Z(n1299) );
AND2_X1 U1013 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND2_X1 U1014 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U1015 ( .A(n1304), .B(n1150), .ZN(n1302) );
XOR2_X1 U1016 ( .A(n1305), .B(KEYINPUT2), .Z(n1300) );
NAND2_X1 U1017 ( .A1(n1146), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1018 ( .A(n1304), .B(n1150), .Z(n1306) );
XOR2_X1 U1019 ( .A(G140), .B(KEYINPUT42), .Z(n1150) );
NOR2_X1 U1020 ( .A1(G110), .A2(KEYINPUT46), .ZN(n1304) );
INV_X1 U1021 ( .A(n1303), .ZN(n1146) );
NAND2_X1 U1022 ( .A1(G227), .A2(n1054), .ZN(n1303) );
NAND2_X1 U1023 ( .A1(n1307), .A2(n1308), .ZN(n1297) );
NAND3_X1 U1024 ( .A1(n1309), .A2(n1235), .A3(n1310), .ZN(n1308) );
INV_X1 U1025 ( .A(KEYINPUT59), .ZN(n1310) );
NAND2_X1 U1026 ( .A1(n1149), .A2(KEYINPUT59), .ZN(n1307) );
XOR2_X1 U1027 ( .A(n1309), .B(n1235), .Z(n1149) );
XNOR2_X1 U1028 ( .A(G131), .B(n1092), .ZN(n1235) );
XOR2_X1 U1029 ( .A(G137), .B(G134), .Z(n1092) );
XOR2_X1 U1030 ( .A(n1311), .B(n1230), .Z(n1309) );
INV_X1 U1031 ( .A(n1090), .ZN(n1230) );
AND2_X1 U1032 ( .A1(n1202), .A2(n1312), .ZN(n1184) );
NAND2_X1 U1033 ( .A1(n1206), .A2(n1313), .ZN(n1312) );
NAND2_X1 U1034 ( .A1(n1208), .A2(n1104), .ZN(n1313) );
INV_X1 U1035 ( .A(G898), .ZN(n1104) );
AND3_X1 U1036 ( .A1(G902), .A2(n1036), .A3(G953), .ZN(n1208) );
NAND3_X1 U1037 ( .A1(n1036), .A2(n1054), .A3(G952), .ZN(n1206) );
INV_X1 U1038 ( .A(G953), .ZN(n1054) );
NAND2_X1 U1039 ( .A1(G234), .A2(G237), .ZN(n1036) );
INV_X1 U1040 ( .A(n1059), .ZN(n1202) );
NAND2_X1 U1041 ( .A1(n1027), .A2(n1076), .ZN(n1059) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1314), .ZN(n1076) );
INV_X1 U1043 ( .A(n1061), .ZN(n1027) );
XNOR2_X1 U1044 ( .A(n1315), .B(n1158), .ZN(n1061) );
NAND2_X1 U1045 ( .A1(G210), .A2(n1314), .ZN(n1158) );
NAND2_X1 U1046 ( .A1(n1231), .A2(n1227), .ZN(n1314) );
INV_X1 U1047 ( .A(G237), .ZN(n1231) );
NAND2_X1 U1048 ( .A1(n1316), .A2(n1227), .ZN(n1315) );
INV_X1 U1049 ( .A(G902), .ZN(n1227) );
XNOR2_X1 U1050 ( .A(n1317), .B(n1155), .ZN(n1316) );
NAND2_X1 U1051 ( .A1(n1318), .A2(n1319), .ZN(n1155) );
NAND2_X1 U1052 ( .A1(n1320), .A2(n1311), .ZN(n1319) );
XOR2_X1 U1053 ( .A(n1107), .B(KEYINPUT32), .Z(n1320) );
NAND2_X1 U1054 ( .A1(n1321), .A2(n1108), .ZN(n1318) );
INV_X1 U1055 ( .A(n1311), .ZN(n1108) );
XOR2_X1 U1056 ( .A(n1322), .B(n1323), .Z(n1311) );
XOR2_X1 U1057 ( .A(G107), .B(G104), .Z(n1323) );
INV_X1 U1058 ( .A(G101), .ZN(n1322) );
XOR2_X1 U1059 ( .A(KEYINPUT38), .B(n1324), .Z(n1321) );
INV_X1 U1060 ( .A(n1107), .ZN(n1324) );
XOR2_X1 U1061 ( .A(n1325), .B(n1326), .Z(n1107) );
XOR2_X1 U1062 ( .A(G113), .B(n1327), .Z(n1326) );
XOR2_X1 U1063 ( .A(G119), .B(G116), .Z(n1327) );
XOR2_X1 U1064 ( .A(n1148), .B(n1265), .Z(n1325) );
XOR2_X1 U1065 ( .A(G122), .B(KEYINPUT57), .Z(n1265) );
INV_X1 U1066 ( .A(G110), .ZN(n1148) );
NAND2_X1 U1067 ( .A1(KEYINPUT11), .A2(n1328), .ZN(n1317) );
XOR2_X1 U1068 ( .A(n1329), .B(n1330), .Z(n1328) );
INV_X1 U1069 ( .A(n1154), .ZN(n1330) );
XOR2_X1 U1070 ( .A(n1090), .B(n1331), .Z(n1154) );
NOR2_X1 U1071 ( .A1(G953), .A2(n1103), .ZN(n1331) );
INV_X1 U1072 ( .A(G224), .ZN(n1103) );
XOR2_X1 U1073 ( .A(n1201), .B(n1332), .Z(n1090) );
XOR2_X1 U1074 ( .A(G146), .B(G143), .Z(n1332) );
INV_X1 U1075 ( .A(G128), .ZN(n1201) );
NOR2_X1 U1076 ( .A1(KEYINPUT29), .A2(n1333), .ZN(n1329) );
XOR2_X1 U1077 ( .A(n1205), .B(KEYINPUT45), .Z(n1333) );
INV_X1 U1078 ( .A(G125), .ZN(n1205) );
endmodule


