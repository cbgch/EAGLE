//Key = 1110110000111010100010111100000001010000101000111111001001111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;

XOR2_X1 U721 ( .A(G107), .B(n1003), .Z(G9) );
NOR4_X1 U722 ( .A1(KEYINPUT3), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1003) );
NOR2_X1 U723 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR3_X1 U724 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
NOR2_X1 U725 ( .A1(n1012), .A2(n1004), .ZN(n1010) );
NOR2_X1 U726 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U727 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
INV_X1 U728 ( .A(n1017), .ZN(n1016) );
NOR2_X1 U729 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
XOR2_X1 U730 ( .A(KEYINPUT17), .B(n1020), .Z(n1019) );
NOR2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR3_X1 U732 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1013) );
NOR4_X1 U733 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025) );
AND2_X1 U734 ( .A1(n1030), .A2(KEYINPUT51), .ZN(n1029) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
NOR3_X1 U736 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1031) );
AND3_X1 U737 ( .A1(KEYINPUT2), .A2(n1036), .A3(n1037), .ZN(n1035) );
NOR2_X1 U738 ( .A1(KEYINPUT2), .A2(n1037), .ZN(n1034) );
AND2_X1 U739 ( .A1(n1038), .A2(n1039), .ZN(n1027) );
NOR2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1024) );
NOR2_X1 U741 ( .A1(KEYINPUT51), .A2(n1042), .ZN(n1041) );
INV_X1 U742 ( .A(n1030), .ZN(n1042) );
INV_X1 U743 ( .A(n1026), .ZN(n1040) );
NAND3_X1 U744 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1009) );
NAND3_X1 U745 ( .A1(n1046), .A2(n1047), .A3(n1017), .ZN(n1045) );
NOR3_X1 U746 ( .A1(n1048), .A2(n1032), .A3(n1026), .ZN(n1017) );
NAND2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U749 ( .A1(n1053), .A2(G953), .A3(G952), .ZN(n1007) );
INV_X1 U750 ( .A(n1043), .ZN(n1053) );
NAND4_X1 U751 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1043) );
NOR4_X1 U752 ( .A1(n1037), .A2(n1058), .A3(n1059), .A4(n1032), .ZN(n1057) );
XNOR2_X1 U753 ( .A(n1060), .B(KEYINPUT61), .ZN(n1059) );
XNOR2_X1 U754 ( .A(n1061), .B(KEYINPUT58), .ZN(n1056) );
XNOR2_X1 U755 ( .A(n1062), .B(n1063), .ZN(n1055) );
XOR2_X1 U756 ( .A(n1064), .B(n1065), .Z(n1054) );
XOR2_X1 U757 ( .A(KEYINPUT54), .B(G469), .Z(n1065) );
NAND2_X1 U758 ( .A1(KEYINPUT48), .A2(n1066), .ZN(n1064) );
XNOR2_X1 U759 ( .A(KEYINPUT50), .B(n1067), .ZN(n1066) );
NAND2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(G72) );
OR3_X1 U761 ( .A1(n1070), .A2(KEYINPUT7), .A3(n1071), .ZN(n1069) );
NAND2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
OR2_X1 U764 ( .A1(n1075), .A2(KEYINPUT34), .ZN(n1074) );
NAND2_X1 U765 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
OR2_X1 U766 ( .A1(KEYINPUT34), .A2(KEYINPUT7), .ZN(n1076) );
INV_X1 U767 ( .A(n1070), .ZN(n1075) );
NAND2_X1 U768 ( .A1(G953), .A2(n1077), .ZN(n1070) );
NAND2_X1 U769 ( .A1(G900), .A2(G227), .ZN(n1077) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1071) );
NAND2_X1 U771 ( .A1(n1080), .A2(n1044), .ZN(n1079) );
XNOR2_X1 U772 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U774 ( .A(n1085), .B(KEYINPUT53), .Z(n1083) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U776 ( .A1(G900), .A2(n1081), .A3(G953), .ZN(n1078) );
XNOR2_X1 U777 ( .A(n1088), .B(n1089), .ZN(n1081) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1089) );
XNOR2_X1 U779 ( .A(KEYINPUT60), .B(n1092), .ZN(n1088) );
NOR2_X1 U780 ( .A1(KEYINPUT13), .A2(n1093), .ZN(n1092) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(G69) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U784 ( .A1(G953), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U785 ( .A(n1101), .B(n1102), .ZN(n1098) );
XNOR2_X1 U786 ( .A(n1103), .B(n1104), .ZN(n1101) );
NOR2_X1 U787 ( .A1(KEYINPUT18), .A2(n1105), .ZN(n1104) );
NAND2_X1 U788 ( .A1(G953), .A2(n1106), .ZN(n1096) );
NAND2_X1 U789 ( .A1(G224), .A2(n1107), .ZN(n1106) );
XNOR2_X1 U790 ( .A(KEYINPUT21), .B(n1100), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1108), .A2(G953), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1115), .ZN(G63) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND3_X1 U797 ( .A1(n1118), .A2(G478), .A3(KEYINPUT49), .ZN(n1116) );
NOR2_X1 U798 ( .A1(n1109), .A2(n1119), .ZN(G60) );
XOR2_X1 U799 ( .A(n1120), .B(n1121), .Z(n1119) );
AND2_X1 U800 ( .A1(G475), .A2(n1118), .ZN(n1120) );
XOR2_X1 U801 ( .A(G104), .B(n1122), .Z(G6) );
NOR2_X1 U802 ( .A1(n1109), .A2(n1123), .ZN(G57) );
XOR2_X1 U803 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U804 ( .A(n1126), .B(n1127), .Z(n1124) );
NOR2_X1 U805 ( .A1(n1063), .A2(n1114), .ZN(n1127) );
NAND2_X1 U806 ( .A1(KEYINPUT42), .A2(n1128), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1109), .A2(n1129), .ZN(G54) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U809 ( .A(n1132), .B(n1133), .ZN(n1131) );
XNOR2_X1 U810 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U811 ( .A(n1136), .B(n1137), .Z(n1130) );
XNOR2_X1 U812 ( .A(n1138), .B(n1139), .ZN(n1137) );
AND2_X1 U813 ( .A1(G469), .A2(n1118), .ZN(n1139) );
NAND2_X1 U814 ( .A1(KEYINPUT33), .A2(n1140), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1109), .A2(n1141), .ZN(G51) );
XOR2_X1 U816 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U817 ( .A(n1144), .B(n1128), .Z(n1143) );
XOR2_X1 U818 ( .A(n1145), .B(n1146), .Z(n1142) );
XNOR2_X1 U819 ( .A(n1147), .B(KEYINPUT27), .ZN(n1146) );
NAND2_X1 U820 ( .A1(KEYINPUT35), .A2(n1148), .ZN(n1147) );
NAND3_X1 U821 ( .A1(n1118), .A2(G210), .A3(KEYINPUT16), .ZN(n1145) );
INV_X1 U822 ( .A(n1114), .ZN(n1118) );
NAND2_X1 U823 ( .A1(G902), .A2(n1011), .ZN(n1114) );
NAND4_X1 U824 ( .A1(n1149), .A2(n1108), .A3(n1150), .A4(n1086), .ZN(n1011) );
AND3_X1 U825 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1086) );
NAND2_X1 U826 ( .A1(n1018), .A2(n1154), .ZN(n1153) );
XOR2_X1 U827 ( .A(KEYINPUT19), .B(n1155), .Z(n1154) );
NAND3_X1 U828 ( .A1(n1046), .A2(n1156), .A3(n1157), .ZN(n1151) );
INV_X1 U829 ( .A(n1084), .ZN(n1150) );
NAND4_X1 U830 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1084) );
NAND3_X1 U831 ( .A1(n1162), .A2(n1038), .A3(n1163), .ZN(n1158) );
XNOR2_X1 U832 ( .A(n1018), .B(KEYINPUT59), .ZN(n1163) );
AND4_X1 U833 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1108) );
NOR4_X1 U834 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR2_X1 U835 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U836 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
INV_X1 U837 ( .A(KEYINPUT57), .ZN(n1175) );
NOR3_X1 U838 ( .A1(n1006), .A2(n1004), .A3(n1005), .ZN(n1169) );
NOR4_X1 U839 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1048), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1018), .A2(n1179), .ZN(n1177) );
NOR4_X1 U841 ( .A1(KEYINPUT57), .A2(n1180), .A3(n1181), .A4(n1004), .ZN(n1179) );
INV_X1 U842 ( .A(n1182), .ZN(n1004) );
NOR2_X1 U843 ( .A1(n1183), .A2(n1172), .ZN(n1176) );
NOR2_X1 U844 ( .A1(n1184), .A2(n1122), .ZN(n1166) );
AND3_X1 U845 ( .A1(n1185), .A2(n1182), .A3(n1038), .ZN(n1122) );
XOR2_X1 U846 ( .A(n1087), .B(KEYINPUT41), .Z(n1149) );
NAND2_X1 U847 ( .A1(n1046), .A2(n1186), .ZN(n1087) );
XOR2_X1 U848 ( .A(KEYINPUT52), .B(n1187), .Z(n1186) );
NOR2_X1 U849 ( .A1(n1044), .A2(G952), .ZN(n1109) );
XNOR2_X1 U850 ( .A(G146), .B(n1188), .ZN(G48) );
NAND3_X1 U851 ( .A1(n1038), .A2(n1018), .A3(n1162), .ZN(n1188) );
XOR2_X1 U852 ( .A(n1159), .B(n1189), .Z(G45) );
NAND2_X1 U853 ( .A1(KEYINPUT4), .A2(G143), .ZN(n1189) );
OR4_X1 U854 ( .A1(n1190), .A2(n1172), .A3(n1181), .A4(n1180), .ZN(n1159) );
XNOR2_X1 U855 ( .A(G140), .B(n1160), .ZN(G42) );
NAND3_X1 U856 ( .A1(n1046), .A2(n1033), .A3(n1191), .ZN(n1160) );
XNOR2_X1 U857 ( .A(G137), .B(n1161), .ZN(G39) );
NAND3_X1 U858 ( .A1(n1046), .A2(n1192), .A3(n1162), .ZN(n1161) );
XOR2_X1 U859 ( .A(G134), .B(n1193), .Z(G36) );
NOR4_X1 U860 ( .A1(KEYINPUT31), .A2(n1006), .A3(n1023), .A4(n1190), .ZN(n1193) );
XNOR2_X1 U861 ( .A(G131), .B(n1194), .ZN(G33) );
NAND2_X1 U862 ( .A1(n1187), .A2(n1046), .ZN(n1194) );
INV_X1 U863 ( .A(n1023), .ZN(n1046) );
NAND2_X1 U864 ( .A1(n1195), .A2(n1060), .ZN(n1023) );
INV_X1 U865 ( .A(n1021), .ZN(n1060) );
AND2_X1 U866 ( .A1(n1157), .A2(n1038), .ZN(n1187) );
INV_X1 U867 ( .A(n1190), .ZN(n1157) );
NAND3_X1 U868 ( .A1(n1033), .A2(n1196), .A3(n1197), .ZN(n1190) );
NAND2_X1 U869 ( .A1(n1198), .A2(n1199), .ZN(G30) );
NAND2_X1 U870 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U871 ( .A(n1202), .B(n1203), .Z(n1198) );
NOR2_X1 U872 ( .A1(n1200), .A2(n1201), .ZN(n1203) );
INV_X1 U873 ( .A(KEYINPUT47), .ZN(n1201) );
NAND2_X1 U874 ( .A1(n1155), .A2(n1018), .ZN(n1202) );
AND2_X1 U875 ( .A1(n1162), .A2(n1156), .ZN(n1155) );
INV_X1 U876 ( .A(n1006), .ZN(n1156) );
AND4_X1 U877 ( .A1(n1033), .A2(n1204), .A3(n1196), .A4(n1052), .ZN(n1162) );
XOR2_X1 U878 ( .A(n1205), .B(n1184), .Z(G3) );
NOR3_X1 U879 ( .A1(n1032), .A2(n1005), .A3(n1049), .ZN(n1184) );
INV_X1 U880 ( .A(n1197), .ZN(n1049) );
NAND2_X1 U881 ( .A1(KEYINPUT20), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U882 ( .A(G125), .B(n1152), .ZN(G27) );
NAND3_X1 U883 ( .A1(n1039), .A2(n1018), .A3(n1191), .ZN(n1152) );
AND4_X1 U884 ( .A1(n1051), .A2(n1038), .A3(n1196), .A4(n1052), .ZN(n1191) );
NAND2_X1 U885 ( .A1(n1026), .A2(n1207), .ZN(n1196) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1209), .ZN(n1207) );
INV_X1 U887 ( .A(G900), .ZN(n1209) );
INV_X1 U888 ( .A(n1172), .ZN(n1018) );
XNOR2_X1 U889 ( .A(G122), .B(n1174), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1039), .A2(n1182), .A3(n1210), .A4(n1211), .ZN(n1174) );
NOR2_X1 U891 ( .A1(n1180), .A2(n1181), .ZN(n1210) );
NOR2_X1 U892 ( .A1(n1052), .A2(n1204), .ZN(n1182) );
XOR2_X1 U893 ( .A(n1212), .B(n1213), .Z(G21) );
AND4_X1 U894 ( .A1(n1214), .A2(n1211), .A3(n1039), .A4(n1183), .ZN(n1213) );
NOR3_X1 U895 ( .A1(n1051), .A2(n1061), .A3(n1032), .ZN(n1183) );
INV_X1 U896 ( .A(n1052), .ZN(n1061) );
INV_X1 U897 ( .A(KEYINPUT56), .ZN(n1214) );
XNOR2_X1 U898 ( .A(G119), .B(KEYINPUT22), .ZN(n1212) );
XNOR2_X1 U899 ( .A(G116), .B(n1164), .ZN(G18) );
NAND3_X1 U900 ( .A1(n1197), .A2(n1211), .A3(n1030), .ZN(n1164) );
NOR2_X1 U901 ( .A1(n1048), .A2(n1006), .ZN(n1030) );
NAND2_X1 U902 ( .A1(n1181), .A2(n1215), .ZN(n1006) );
XNOR2_X1 U903 ( .A(n1216), .B(n1217), .ZN(G15) );
NOR3_X1 U904 ( .A1(n1218), .A2(KEYINPUT55), .A3(n1172), .ZN(n1217) );
XNOR2_X1 U905 ( .A(KEYINPUT1), .B(n1173), .ZN(n1218) );
NAND4_X1 U906 ( .A1(n1039), .A2(n1038), .A3(n1197), .A4(n1219), .ZN(n1173) );
NOR2_X1 U907 ( .A1(n1052), .A2(n1051), .ZN(n1197) );
NOR2_X1 U908 ( .A1(n1215), .A2(n1181), .ZN(n1038) );
INV_X1 U909 ( .A(n1048), .ZN(n1039) );
NAND2_X1 U910 ( .A1(n1220), .A2(n1036), .ZN(n1048) );
XNOR2_X1 U911 ( .A(n1037), .B(KEYINPUT29), .ZN(n1220) );
XOR2_X1 U912 ( .A(n1165), .B(n1221), .Z(G12) );
NAND2_X1 U913 ( .A1(KEYINPUT62), .A2(G110), .ZN(n1221) );
NAND4_X1 U914 ( .A1(n1192), .A2(n1185), .A3(n1051), .A4(n1052), .ZN(n1165) );
NAND3_X1 U915 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1052) );
NAND2_X1 U916 ( .A1(n1225), .A2(n1111), .ZN(n1224) );
OR3_X1 U917 ( .A1(n1111), .A2(n1225), .A3(G902), .ZN(n1223) );
NOR2_X1 U918 ( .A1(n1113), .A2(G234), .ZN(n1225) );
INV_X1 U919 ( .A(G217), .ZN(n1113) );
XOR2_X1 U920 ( .A(n1226), .B(n1227), .Z(n1111) );
XOR2_X1 U921 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U922 ( .A(G146), .B(KEYINPUT25), .ZN(n1229) );
NAND2_X1 U923 ( .A1(n1230), .A2(n1231), .ZN(n1228) );
NAND2_X1 U924 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U925 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U926 ( .A1(KEYINPUT14), .A2(n1236), .ZN(n1235) );
INV_X1 U927 ( .A(KEYINPUT44), .ZN(n1234) );
NAND2_X1 U928 ( .A1(n1135), .A2(n1237), .ZN(n1230) );
NAND2_X1 U929 ( .A1(KEYINPUT14), .A2(n1238), .ZN(n1237) );
OR2_X1 U930 ( .A1(n1232), .A2(KEYINPUT44), .ZN(n1238) );
XNOR2_X1 U931 ( .A(G119), .B(n1200), .ZN(n1232) );
INV_X1 U932 ( .A(G128), .ZN(n1200) );
INV_X1 U933 ( .A(n1236), .ZN(n1135) );
XOR2_X1 U934 ( .A(n1239), .B(n1091), .Z(n1226) );
XNOR2_X1 U935 ( .A(n1148), .B(G140), .ZN(n1091) );
NAND2_X1 U936 ( .A1(KEYINPUT40), .A2(n1240), .ZN(n1239) );
XNOR2_X1 U937 ( .A(G137), .B(n1241), .ZN(n1240) );
NAND2_X1 U938 ( .A1(G221), .A2(n1242), .ZN(n1241) );
NAND2_X1 U939 ( .A1(G902), .A2(G217), .ZN(n1222) );
INV_X1 U940 ( .A(n1204), .ZN(n1051) );
XNOR2_X1 U941 ( .A(n1062), .B(n1243), .ZN(n1204) );
NOR2_X1 U942 ( .A1(KEYINPUT43), .A2(n1063), .ZN(n1243) );
INV_X1 U943 ( .A(G472), .ZN(n1063) );
NAND2_X1 U944 ( .A1(n1244), .A2(n1245), .ZN(n1062) );
XNOR2_X1 U945 ( .A(n1125), .B(n1246), .ZN(n1244) );
XNOR2_X1 U946 ( .A(n1128), .B(KEYINPUT26), .ZN(n1246) );
XNOR2_X1 U947 ( .A(n1247), .B(n1248), .ZN(n1125) );
XOR2_X1 U948 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U949 ( .A(n1251), .B(n1206), .ZN(n1250) );
INV_X1 U950 ( .A(G101), .ZN(n1206) );
NAND2_X1 U951 ( .A1(KEYINPUT46), .A2(n1216), .ZN(n1251) );
NAND2_X1 U952 ( .A1(G210), .A2(n1252), .ZN(n1249) );
XNOR2_X1 U953 ( .A(n1253), .B(n1090), .ZN(n1247) );
INV_X1 U954 ( .A(n1005), .ZN(n1185) );
NAND2_X1 U955 ( .A1(n1033), .A2(n1211), .ZN(n1005) );
NOR2_X1 U956 ( .A1(n1172), .A2(n1178), .ZN(n1211) );
INV_X1 U957 ( .A(n1219), .ZN(n1178) );
NAND2_X1 U958 ( .A1(n1026), .A2(n1254), .ZN(n1219) );
NAND4_X1 U959 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1100), .ZN(n1254) );
INV_X1 U960 ( .A(G898), .ZN(n1100) );
NAND3_X1 U961 ( .A1(n1208), .A2(n1044), .A3(G952), .ZN(n1026) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1208) );
NAND2_X1 U963 ( .A1(n1195), .A2(n1255), .ZN(n1172) );
XNOR2_X1 U964 ( .A(KEYINPUT0), .B(n1021), .ZN(n1255) );
NAND3_X1 U965 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1021) );
OR2_X1 U966 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND3_X1 U967 ( .A1(n1260), .A2(n1259), .A3(n1245), .ZN(n1257) );
NAND2_X1 U968 ( .A1(G237), .A2(G210), .ZN(n1259) );
XNOR2_X1 U969 ( .A(n1144), .B(n1261), .ZN(n1260) );
XNOR2_X1 U970 ( .A(n1148), .B(n1262), .ZN(n1261) );
NOR2_X1 U971 ( .A1(KEYINPUT36), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U972 ( .A(n1128), .B(KEYINPUT15), .ZN(n1263) );
XOR2_X1 U973 ( .A(n1264), .B(n1265), .Z(n1128) );
XOR2_X1 U974 ( .A(G143), .B(n1266), .Z(n1265) );
NOR2_X1 U975 ( .A1(G146), .A2(KEYINPUT30), .ZN(n1266) );
XOR2_X1 U976 ( .A(n1267), .B(n1103), .Z(n1144) );
XOR2_X1 U977 ( .A(G122), .B(n1236), .Z(n1103) );
XOR2_X1 U978 ( .A(n1268), .B(n1269), .Z(n1267) );
AND2_X1 U979 ( .A1(n1044), .A2(G224), .ZN(n1269) );
NAND3_X1 U980 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1268) );
NAND2_X1 U981 ( .A1(n1105), .A2(n1273), .ZN(n1272) );
NAND2_X1 U982 ( .A1(n1274), .A2(KEYINPUT11), .ZN(n1273) );
XOR2_X1 U983 ( .A(n1102), .B(KEYINPUT39), .Z(n1274) );
NAND3_X1 U984 ( .A1(KEYINPUT11), .A2(n1275), .A3(n1102), .ZN(n1271) );
INV_X1 U985 ( .A(n1105), .ZN(n1275) );
XOR2_X1 U986 ( .A(n1276), .B(n1216), .Z(n1105) );
NAND2_X1 U987 ( .A1(KEYINPUT12), .A2(n1277), .ZN(n1276) );
XOR2_X1 U988 ( .A(KEYINPUT32), .B(n1253), .Z(n1277) );
XNOR2_X1 U989 ( .A(G116), .B(n1278), .ZN(n1253) );
INV_X1 U990 ( .A(G119), .ZN(n1278) );
OR2_X1 U991 ( .A1(n1102), .A2(KEYINPUT11), .ZN(n1270) );
XOR2_X1 U992 ( .A(n1279), .B(n1280), .Z(n1102) );
NOR2_X1 U993 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1280) );
NAND2_X1 U994 ( .A1(G902), .A2(G210), .ZN(n1256) );
XNOR2_X1 U995 ( .A(KEYINPUT38), .B(n1058), .ZN(n1195) );
INV_X1 U996 ( .A(n1022), .ZN(n1058) );
NAND2_X1 U997 ( .A1(G214), .A2(n1281), .ZN(n1022) );
OR2_X1 U998 ( .A1(G237), .A2(G902), .ZN(n1281) );
NOR2_X1 U999 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
AND2_X1 U1000 ( .A1(G221), .A2(n1282), .ZN(n1037) );
NAND2_X1 U1001 ( .A1(G234), .A2(n1245), .ZN(n1282) );
XOR2_X1 U1002 ( .A(n1067), .B(n1283), .Z(n1036) );
XOR2_X1 U1003 ( .A(KEYINPUT9), .B(G469), .Z(n1283) );
NAND3_X1 U1004 ( .A1(n1284), .A2(n1285), .A3(n1245), .ZN(n1067) );
NAND2_X1 U1005 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
INV_X1 U1006 ( .A(KEYINPUT6), .ZN(n1287) );
XOR2_X1 U1007 ( .A(n1288), .B(n1289), .Z(n1286) );
NAND3_X1 U1008 ( .A1(n1289), .A2(n1288), .A3(KEYINPUT6), .ZN(n1284) );
XOR2_X1 U1009 ( .A(n1134), .B(n1290), .Z(n1288) );
XNOR2_X1 U1010 ( .A(G104), .B(n1093), .ZN(n1290) );
INV_X1 U1011 ( .A(n1140), .ZN(n1093) );
XOR2_X1 U1012 ( .A(n1291), .B(n1264), .Z(n1140) );
XOR2_X1 U1013 ( .A(G128), .B(KEYINPUT45), .Z(n1264) );
XOR2_X1 U1014 ( .A(n1279), .B(n1090), .Z(n1134) );
XNOR2_X1 U1015 ( .A(n1292), .B(n1293), .ZN(n1090) );
XNOR2_X1 U1016 ( .A(G131), .B(G137), .ZN(n1292) );
XNOR2_X1 U1017 ( .A(G101), .B(n1294), .ZN(n1279) );
XOR2_X1 U1018 ( .A(KEYINPUT5), .B(G107), .Z(n1294) );
AND3_X1 U1019 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1289) );
NAND2_X1 U1020 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1021 ( .A1(n1300), .A2(KEYINPUT24), .ZN(n1299) );
XOR2_X1 U1022 ( .A(n1138), .B(KEYINPUT63), .Z(n1300) );
XNOR2_X1 U1023 ( .A(n1301), .B(n1236), .ZN(n1298) );
OR2_X1 U1024 ( .A1(n1138), .A2(KEYINPUT24), .ZN(n1296) );
NAND3_X1 U1025 ( .A1(n1302), .A2(n1138), .A3(KEYINPUT24), .ZN(n1295) );
NAND2_X1 U1026 ( .A1(G227), .A2(n1044), .ZN(n1138) );
XNOR2_X1 U1027 ( .A(G140), .B(n1236), .ZN(n1302) );
XOR2_X1 U1028 ( .A(G110), .B(KEYINPUT10), .Z(n1236) );
INV_X1 U1029 ( .A(n1032), .ZN(n1192) );
NAND2_X1 U1030 ( .A1(n1180), .A2(n1181), .ZN(n1032) );
XOR2_X1 U1031 ( .A(n1303), .B(G475), .Z(n1181) );
OR2_X1 U1032 ( .A1(n1121), .A2(G902), .ZN(n1303) );
XNOR2_X1 U1033 ( .A(n1304), .B(n1305), .ZN(n1121) );
XOR2_X1 U1034 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U1035 ( .A(n1308), .B(n1216), .ZN(n1307) );
INV_X1 U1036 ( .A(G113), .ZN(n1216) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1252), .ZN(n1308) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1252) );
XNOR2_X1 U1039 ( .A(G131), .B(G122), .ZN(n1306) );
XOR2_X1 U1040 ( .A(n1309), .B(n1132), .Z(n1304) );
XNOR2_X1 U1041 ( .A(G104), .B(n1301), .ZN(n1132) );
INV_X1 U1042 ( .A(G140), .ZN(n1301) );
XOR2_X1 U1043 ( .A(n1310), .B(n1291), .Z(n1309) );
XNOR2_X1 U1044 ( .A(G143), .B(n1311), .ZN(n1291) );
INV_X1 U1045 ( .A(G146), .ZN(n1311) );
NAND2_X1 U1046 ( .A1(KEYINPUT23), .A2(n1148), .ZN(n1310) );
INV_X1 U1047 ( .A(G125), .ZN(n1148) );
INV_X1 U1048 ( .A(n1215), .ZN(n1180) );
XNOR2_X1 U1049 ( .A(n1312), .B(G478), .ZN(n1215) );
NAND2_X1 U1050 ( .A1(n1117), .A2(n1245), .ZN(n1312) );
INV_X1 U1051 ( .A(G902), .ZN(n1245) );
XNOR2_X1 U1052 ( .A(n1313), .B(n1314), .ZN(n1117) );
XOR2_X1 U1053 ( .A(G107), .B(n1315), .Z(n1314) );
XNOR2_X1 U1054 ( .A(n1316), .B(G116), .ZN(n1315) );
INV_X1 U1055 ( .A(G122), .ZN(n1316) );
XOR2_X1 U1056 ( .A(n1317), .B(n1318), .Z(n1313) );
NOR2_X1 U1057 ( .A1(KEYINPUT28), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1058 ( .A(n1320), .B(n1293), .Z(n1319) );
XOR2_X1 U1059 ( .A(G134), .B(KEYINPUT37), .Z(n1293) );
XNOR2_X1 U1060 ( .A(G128), .B(G143), .ZN(n1320) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1242), .ZN(n1317) );
AND2_X1 U1062 ( .A1(G234), .A2(n1044), .ZN(n1242) );
INV_X1 U1063 ( .A(G953), .ZN(n1044) );
endmodule


