//Key = 0100001010010000011001101001000101101011001101000010010100111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;

XNOR2_X1 U773 ( .A(G107), .B(n1072), .ZN(G9) );
NOR2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(G75) );
NOR4_X1 U775 ( .A1(n1075), .A2(n1076), .A3(G953), .A4(n1077), .ZN(n1074) );
NOR3_X1 U776 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1076) );
NOR2_X1 U777 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
INV_X1 U778 ( .A(n1083), .ZN(n1078) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1075) );
NAND3_X1 U780 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NAND3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NAND2_X1 U784 ( .A1(KEYINPUT40), .A2(n1096), .ZN(n1094) );
NAND4_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1091) );
INV_X1 U786 ( .A(n1095), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1101), .ZN(n1099) );
INV_X1 U788 ( .A(KEYINPUT40), .ZN(n1101) );
NAND3_X1 U789 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1098) );
XNOR2_X1 U790 ( .A(n1105), .B(KEYINPUT62), .ZN(n1104) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1097) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U793 ( .A1(n1083), .A2(n1110), .ZN(n1089) );
NAND2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR3_X1 U796 ( .A1(n1115), .A2(n1116), .A3(n1095), .ZN(n1083) );
NOR3_X1 U797 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1073) );
AND4_X1 U798 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1077) );
NOR4_X1 U799 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U801 ( .A1(n1113), .A2(n1103), .ZN(n1119) );
XOR2_X1 U802 ( .A(n1127), .B(n1128), .Z(n1118) );
XOR2_X1 U803 ( .A(KEYINPUT44), .B(G469), .Z(n1128) );
NOR2_X1 U804 ( .A1(n1129), .A2(KEYINPUT14), .ZN(n1127) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(G72) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR3_X1 U807 ( .A1(n1134), .A2(G953), .A3(n1135), .ZN(n1133) );
XNOR2_X1 U808 ( .A(KEYINPUT42), .B(KEYINPUT30), .ZN(n1134) );
NAND2_X1 U809 ( .A1(n1136), .A2(n1137), .ZN(n1132) );
NAND2_X1 U810 ( .A1(G953), .A2(n1138), .ZN(n1137) );
XOR2_X1 U811 ( .A(n1139), .B(n1140), .Z(n1136) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NOR2_X1 U814 ( .A1(KEYINPUT47), .A2(n1145), .ZN(n1144) );
AND2_X1 U815 ( .A1(KEYINPUT51), .A2(n1145), .ZN(n1143) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(n1145) );
XNOR2_X1 U817 ( .A(n1148), .B(G134), .ZN(n1147) );
NAND2_X1 U818 ( .A1(G953), .A2(n1149), .ZN(n1130) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1149) );
NAND2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1160), .A2(G953), .ZN(n1150) );
XOR2_X1 U826 ( .A(n1161), .B(n1158), .Z(n1160) );
XOR2_X1 U827 ( .A(n1156), .B(KEYINPUT50), .Z(n1158) );
NAND3_X1 U828 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1156) );
NAND2_X1 U829 ( .A1(G953), .A2(n1165), .ZN(n1164) );
NAND2_X1 U830 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
INV_X1 U831 ( .A(KEYINPUT60), .ZN(n1167) );
NAND2_X1 U832 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NAND2_X1 U833 ( .A1(KEYINPUT60), .A2(n1170), .ZN(n1162) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1161) );
NOR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(G66) );
XOR2_X1 U836 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND3_X1 U837 ( .A1(G217), .A2(n1175), .A3(G902), .ZN(n1173) );
XNOR2_X1 U838 ( .A(KEYINPUT45), .B(n1176), .ZN(n1175) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1177), .ZN(G63) );
XOR2_X1 U840 ( .A(n1178), .B(n1179), .Z(n1177) );
NAND2_X1 U841 ( .A1(n1180), .A2(G478), .ZN(n1178) );
NOR2_X1 U842 ( .A1(n1171), .A2(n1181), .ZN(G60) );
XOR2_X1 U843 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U844 ( .A1(n1180), .A2(G475), .ZN(n1182) );
XOR2_X1 U845 ( .A(G104), .B(n1184), .Z(G6) );
NOR2_X1 U846 ( .A1(n1185), .A2(n1186), .ZN(G57) );
XOR2_X1 U847 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U848 ( .A(n1189), .B(G101), .ZN(n1188) );
NAND3_X1 U849 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1187) );
NAND2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
OR4_X1 U851 ( .A1(n1193), .A2(KEYINPUT19), .A3(n1194), .A4(n1195), .ZN(n1191) );
INV_X1 U852 ( .A(KEYINPUT6), .ZN(n1194) );
NAND2_X1 U853 ( .A1(n1180), .A2(G472), .ZN(n1193) );
NAND2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1190) );
NAND3_X1 U855 ( .A1(G472), .A2(n1197), .A3(n1180), .ZN(n1196) );
INV_X1 U856 ( .A(KEYINPUT19), .ZN(n1197) );
XOR2_X1 U857 ( .A(n1198), .B(n1199), .Z(n1195) );
XNOR2_X1 U858 ( .A(n1200), .B(n1201), .ZN(n1199) );
NOR2_X1 U859 ( .A1(KEYINPUT2), .A2(n1202), .ZN(n1201) );
NAND2_X1 U860 ( .A1(KEYINPUT33), .A2(n1203), .ZN(n1200) );
NOR2_X1 U861 ( .A1(G952), .A2(n1204), .ZN(n1185) );
XNOR2_X1 U862 ( .A(KEYINPUT21), .B(n1153), .ZN(n1204) );
NOR2_X1 U863 ( .A1(n1171), .A2(n1205), .ZN(G54) );
XNOR2_X1 U864 ( .A(n1206), .B(n1207), .ZN(n1205) );
XOR2_X1 U865 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR4_X1 U866 ( .A1(KEYINPUT3), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1209) );
INV_X1 U867 ( .A(n1213), .ZN(n1211) );
NAND2_X1 U868 ( .A1(n1180), .A2(G469), .ZN(n1208) );
NOR2_X1 U869 ( .A1(n1171), .A2(n1214), .ZN(G51) );
NOR2_X1 U870 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NOR2_X1 U871 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U872 ( .A(KEYINPUT20), .B(n1219), .Z(n1218) );
NOR2_X1 U873 ( .A1(n1125), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U874 ( .A(KEYINPUT48), .B(n1221), .ZN(n1217) );
NOR3_X1 U875 ( .A1(n1221), .A2(n1125), .A3(n1220), .ZN(n1215) );
INV_X1 U876 ( .A(n1180), .ZN(n1220) );
NOR2_X1 U877 ( .A1(n1222), .A2(n1084), .ZN(n1180) );
INV_X1 U878 ( .A(n1176), .ZN(n1084) );
NAND2_X1 U879 ( .A1(n1135), .A2(n1159), .ZN(n1176) );
INV_X1 U880 ( .A(n1157), .ZN(n1159) );
NAND4_X1 U881 ( .A1(n1223), .A2(n1072), .A3(n1224), .A4(n1225), .ZN(n1157) );
NOR3_X1 U882 ( .A1(n1184), .A2(n1226), .A3(n1227), .ZN(n1225) );
AND4_X1 U883 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1184) );
NAND2_X1 U884 ( .A1(n1231), .A2(n1232), .ZN(n1224) );
NAND2_X1 U885 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND3_X1 U886 ( .A1(n1106), .A2(n1228), .A3(n1235), .ZN(n1234) );
XNOR2_X1 U887 ( .A(KEYINPUT24), .B(n1236), .ZN(n1233) );
NAND4_X1 U888 ( .A1(n1237), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1072) );
INV_X1 U889 ( .A(n1238), .ZN(n1230) );
NAND3_X1 U890 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1223) );
NAND2_X1 U891 ( .A1(n1242), .A2(n1243), .ZN(n1239) );
NAND4_X1 U892 ( .A1(n1244), .A2(n1088), .A3(n1245), .A4(n1086), .ZN(n1243) );
NOR2_X1 U893 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U894 ( .A(n1106), .B(KEYINPUT61), .ZN(n1244) );
NAND3_X1 U895 ( .A1(n1106), .A2(n1248), .A3(n1105), .ZN(n1242) );
AND2_X1 U896 ( .A1(n1249), .A2(n1250), .ZN(n1135) );
AND4_X1 U897 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
NOR4_X1 U898 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1249) );
NOR3_X1 U899 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
NOR2_X1 U900 ( .A1(KEYINPUT1), .A2(n1262), .ZN(n1261) );
NOR2_X1 U901 ( .A1(n1263), .A2(n1229), .ZN(n1262) );
INV_X1 U902 ( .A(n1264), .ZN(n1263) );
NOR2_X1 U903 ( .A1(n1265), .A2(n1266), .ZN(n1260) );
INV_X1 U904 ( .A(KEYINPUT1), .ZN(n1266) );
INV_X1 U905 ( .A(n1267), .ZN(n1257) );
XOR2_X1 U906 ( .A(n1170), .B(n1268), .Z(n1221) );
NOR3_X1 U907 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1268) );
NOR2_X1 U908 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
AND2_X1 U909 ( .A1(n1274), .A2(KEYINPUT27), .ZN(n1272) );
AND4_X1 U910 ( .A1(n1273), .A2(KEYINPUT43), .A3(n1274), .A4(KEYINPUT27), .ZN(n1270) );
NOR2_X1 U911 ( .A1(KEYINPUT43), .A2(n1274), .ZN(n1269) );
XNOR2_X1 U912 ( .A(n1275), .B(KEYINPUT15), .ZN(n1274) );
NOR2_X1 U913 ( .A1(n1153), .A2(G952), .ZN(n1171) );
XNOR2_X1 U914 ( .A(G146), .B(n1251), .ZN(G48) );
NAND4_X1 U915 ( .A1(n1228), .A2(n1265), .A3(n1241), .A4(n1248), .ZN(n1251) );
XOR2_X1 U916 ( .A(G143), .B(n1276), .Z(G45) );
NOR2_X1 U917 ( .A1(KEYINPUT13), .A2(n1267), .ZN(n1276) );
NAND3_X1 U918 ( .A1(n1082), .A2(n1265), .A3(n1277), .ZN(n1267) );
NOR3_X1 U919 ( .A1(n1111), .A2(n1246), .A3(n1247), .ZN(n1277) );
XOR2_X1 U920 ( .A(G140), .B(n1256), .Z(G42) );
AND2_X1 U921 ( .A1(n1278), .A2(n1279), .ZN(n1256) );
XOR2_X1 U922 ( .A(n1280), .B(n1281), .Z(G39) );
NAND2_X1 U923 ( .A1(KEYINPUT58), .A2(n1148), .ZN(n1281) );
INV_X1 U924 ( .A(G137), .ZN(n1148) );
NAND2_X1 U925 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND4_X1 U926 ( .A1(n1229), .A2(n1248), .A3(n1093), .A4(n1284), .ZN(n1283) );
NOR3_X1 U927 ( .A1(n1264), .A2(n1115), .A3(n1285), .ZN(n1284) );
NAND2_X1 U928 ( .A1(n1255), .A2(n1285), .ZN(n1282) );
INV_X1 U929 ( .A(KEYINPUT7), .ZN(n1285) );
AND3_X1 U930 ( .A1(n1278), .A2(n1248), .A3(n1105), .ZN(n1255) );
XOR2_X1 U931 ( .A(n1286), .B(n1287), .Z(G36) );
XOR2_X1 U932 ( .A(KEYINPUT39), .B(G134), .Z(n1287) );
NAND2_X1 U933 ( .A1(n1288), .A2(n1265), .ZN(n1286) );
INV_X1 U934 ( .A(n1259), .ZN(n1288) );
NAND3_X1 U935 ( .A1(n1093), .A2(n1237), .A3(n1082), .ZN(n1259) );
XNOR2_X1 U936 ( .A(G131), .B(n1254), .ZN(G33) );
NAND3_X1 U937 ( .A1(n1278), .A2(n1228), .A3(n1082), .ZN(n1254) );
AND2_X1 U938 ( .A1(n1093), .A2(n1265), .ZN(n1278) );
INV_X1 U939 ( .A(n1080), .ZN(n1093) );
NAND2_X1 U940 ( .A1(n1114), .A2(n1289), .ZN(n1080) );
XNOR2_X1 U941 ( .A(G128), .B(n1253), .ZN(G30) );
NAND4_X1 U942 ( .A1(n1265), .A2(n1237), .A3(n1241), .A4(n1248), .ZN(n1253) );
INV_X1 U943 ( .A(n1109), .ZN(n1237) );
AND2_X1 U944 ( .A1(n1229), .A2(n1264), .ZN(n1265) );
XOR2_X1 U945 ( .A(G101), .B(n1290), .Z(G3) );
NOR2_X1 U946 ( .A1(n1291), .A2(n1236), .ZN(n1290) );
NAND2_X1 U947 ( .A1(n1235), .A2(n1096), .ZN(n1236) );
INV_X1 U948 ( .A(n1292), .ZN(n1235) );
XNOR2_X1 U949 ( .A(G125), .B(n1252), .ZN(G27) );
NAND4_X1 U950 ( .A1(n1106), .A2(n1279), .A3(n1241), .A4(n1264), .ZN(n1252) );
NAND2_X1 U951 ( .A1(n1095), .A2(n1293), .ZN(n1264) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1138), .ZN(n1293) );
INV_X1 U953 ( .A(G900), .ZN(n1138) );
AND2_X1 U954 ( .A1(n1228), .A2(n1081), .ZN(n1279) );
XNOR2_X1 U955 ( .A(G122), .B(n1295), .ZN(G24) );
NAND3_X1 U956 ( .A1(n1296), .A2(n1106), .A3(n1297), .ZN(n1295) );
NOR3_X1 U957 ( .A1(n1238), .A2(n1246), .A3(n1247), .ZN(n1297) );
NAND3_X1 U958 ( .A1(n1086), .A2(n1240), .A3(n1088), .ZN(n1238) );
XNOR2_X1 U959 ( .A(n1122), .B(KEYINPUT56), .ZN(n1086) );
XNOR2_X1 U960 ( .A(n1241), .B(KEYINPUT17), .ZN(n1296) );
XOR2_X1 U961 ( .A(n1298), .B(n1299), .Z(G21) );
XNOR2_X1 U962 ( .A(G119), .B(KEYINPUT12), .ZN(n1299) );
NAND4_X1 U963 ( .A1(n1300), .A2(n1240), .A3(n1241), .A4(n1301), .ZN(n1298) );
NOR2_X1 U964 ( .A1(n1116), .A2(n1115), .ZN(n1301) );
XOR2_X1 U965 ( .A(n1248), .B(KEYINPUT16), .Z(n1300) );
NAND2_X1 U966 ( .A1(n1302), .A2(n1303), .ZN(n1248) );
NAND3_X1 U967 ( .A1(n1122), .A2(n1121), .A3(n1304), .ZN(n1303) );
INV_X1 U968 ( .A(KEYINPUT25), .ZN(n1304) );
NAND2_X1 U969 ( .A1(KEYINPUT25), .A2(n1081), .ZN(n1302) );
XOR2_X1 U970 ( .A(n1227), .B(n1305), .Z(G18) );
NOR2_X1 U971 ( .A1(KEYINPUT10), .A2(n1306), .ZN(n1305) );
NOR4_X1 U972 ( .A1(n1292), .A2(n1116), .A3(n1109), .A4(n1111), .ZN(n1227) );
INV_X1 U973 ( .A(n1241), .ZN(n1111) );
NAND2_X1 U974 ( .A1(n1247), .A2(n1123), .ZN(n1109) );
XOR2_X1 U975 ( .A(n1307), .B(n1308), .Z(G15) );
NOR2_X1 U976 ( .A1(KEYINPUT41), .A2(n1309), .ZN(n1308) );
NOR4_X1 U977 ( .A1(n1291), .A2(n1310), .A3(n1108), .A4(n1292), .ZN(n1307) );
NAND2_X1 U978 ( .A1(n1082), .A2(n1240), .ZN(n1292) );
AND2_X1 U979 ( .A1(n1088), .A2(n1122), .ZN(n1082) );
INV_X1 U980 ( .A(n1228), .ZN(n1108) );
NOR2_X1 U981 ( .A1(n1123), .A2(n1247), .ZN(n1228) );
XNOR2_X1 U982 ( .A(n1106), .B(KEYINPUT54), .ZN(n1310) );
INV_X1 U983 ( .A(n1116), .ZN(n1106) );
NAND2_X1 U984 ( .A1(n1102), .A2(n1311), .ZN(n1116) );
INV_X1 U985 ( .A(n1231), .ZN(n1291) );
XOR2_X1 U986 ( .A(G110), .B(n1226), .Z(G12) );
AND4_X1 U987 ( .A1(n1096), .A2(n1081), .A3(n1231), .A4(n1240), .ZN(n1226) );
NAND2_X1 U988 ( .A1(n1095), .A2(n1312), .ZN(n1240) );
NAND4_X1 U989 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1165), .ZN(n1312) );
INV_X1 U990 ( .A(G898), .ZN(n1165) );
NAND3_X1 U991 ( .A1(n1294), .A2(n1153), .A3(G952), .ZN(n1095) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1294) );
XOR2_X1 U993 ( .A(n1241), .B(KEYINPUT35), .Z(n1231) );
NOR2_X1 U994 ( .A1(n1114), .A2(n1113), .ZN(n1241) );
INV_X1 U995 ( .A(n1289), .ZN(n1113) );
NAND2_X1 U996 ( .A1(n1313), .A2(G214), .ZN(n1289) );
XOR2_X1 U997 ( .A(n1314), .B(KEYINPUT4), .Z(n1313) );
XOR2_X1 U998 ( .A(n1315), .B(n1126), .Z(n1114) );
NAND3_X1 U999 ( .A1(n1316), .A2(n1222), .A3(n1317), .ZN(n1126) );
XOR2_X1 U1000 ( .A(KEYINPUT55), .B(n1318), .Z(n1317) );
NOR2_X1 U1001 ( .A1(n1170), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1002 ( .A1(n1170), .A2(n1319), .ZN(n1316) );
XOR2_X1 U1003 ( .A(n1320), .B(n1273), .Z(n1319) );
XNOR2_X1 U1004 ( .A(n1198), .B(n1321), .ZN(n1273) );
XOR2_X1 U1005 ( .A(n1275), .B(KEYINPUT38), .Z(n1320) );
NAND2_X1 U1006 ( .A1(G224), .A2(n1153), .ZN(n1275) );
XNOR2_X1 U1007 ( .A(n1169), .B(n1168), .ZN(n1170) );
XOR2_X1 U1008 ( .A(G122), .B(n1322), .Z(n1168) );
XOR2_X1 U1009 ( .A(n1323), .B(n1324), .Z(n1169) );
NOR2_X1 U1010 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NOR3_X1 U1011 ( .A1(n1327), .A2(G119), .A3(n1306), .ZN(n1326) );
INV_X1 U1012 ( .A(KEYINPUT23), .ZN(n1327) );
NOR2_X1 U1013 ( .A1(KEYINPUT23), .A2(n1328), .ZN(n1325) );
XNOR2_X1 U1014 ( .A(n1329), .B(n1309), .ZN(n1323) );
NAND2_X1 U1015 ( .A1(n1330), .A2(KEYINPUT8), .ZN(n1315) );
XOR2_X1 U1016 ( .A(n1125), .B(KEYINPUT57), .Z(n1330) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1314), .ZN(n1125) );
NAND2_X1 U1018 ( .A1(n1222), .A2(n1331), .ZN(n1314) );
INV_X1 U1019 ( .A(G237), .ZN(n1331) );
NOR2_X1 U1020 ( .A1(n1122), .A2(n1088), .ZN(n1081) );
INV_X1 U1021 ( .A(n1121), .ZN(n1088) );
NAND3_X1 U1022 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1121) );
OR2_X1 U1023 ( .A1(n1335), .A2(n1174), .ZN(n1334) );
NAND3_X1 U1024 ( .A1(n1174), .A2(n1335), .A3(n1222), .ZN(n1333) );
NAND2_X1 U1025 ( .A1(G217), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1026 ( .A(n1337), .B(n1338), .Z(n1174) );
XOR2_X1 U1027 ( .A(n1339), .B(n1340), .Z(n1338) );
XNOR2_X1 U1028 ( .A(n1341), .B(G137), .ZN(n1340) );
INV_X1 U1029 ( .A(G146), .ZN(n1341) );
NOR2_X1 U1030 ( .A1(KEYINPUT46), .A2(n1342), .ZN(n1339) );
XNOR2_X1 U1031 ( .A(n1343), .B(G119), .ZN(n1342) );
XOR2_X1 U1032 ( .A(n1344), .B(n1141), .Z(n1337) );
XOR2_X1 U1033 ( .A(n1345), .B(n1346), .Z(n1344) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1347), .ZN(n1345) );
NAND2_X1 U1035 ( .A1(G902), .A2(G217), .ZN(n1332) );
XNOR2_X1 U1036 ( .A(n1348), .B(G472), .ZN(n1122) );
NAND2_X1 U1037 ( .A1(n1349), .A2(n1222), .ZN(n1348) );
XOR2_X1 U1038 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1039 ( .A(n1352), .B(KEYINPUT11), .Z(n1351) );
NAND2_X1 U1040 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1041 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1042 ( .A1(KEYINPUT31), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1043 ( .A1(n1203), .A2(n1358), .ZN(n1357) );
INV_X1 U1044 ( .A(n1359), .ZN(n1355) );
NAND2_X1 U1045 ( .A1(n1360), .A2(n1361), .ZN(n1353) );
NAND2_X1 U1046 ( .A1(n1358), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1047 ( .A1(KEYINPUT31), .A2(n1359), .ZN(n1362) );
XNOR2_X1 U1048 ( .A(n1202), .B(n1198), .ZN(n1359) );
XNOR2_X1 U1049 ( .A(G128), .B(n1363), .ZN(n1198) );
INV_X1 U1050 ( .A(KEYINPUT9), .ZN(n1358) );
INV_X1 U1051 ( .A(n1203), .ZN(n1360) );
XOR2_X1 U1052 ( .A(G113), .B(n1328), .Z(n1203) );
XNOR2_X1 U1053 ( .A(n1306), .B(G119), .ZN(n1328) );
NAND3_X1 U1054 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1350) );
NAND2_X1 U1055 ( .A1(n1189), .A2(G101), .ZN(n1366) );
NAND2_X1 U1056 ( .A1(n1367), .A2(n1368), .ZN(n1365) );
INV_X1 U1057 ( .A(KEYINPUT36), .ZN(n1368) );
NAND2_X1 U1058 ( .A1(n1369), .A2(n1370), .ZN(n1367) );
XNOR2_X1 U1059 ( .A(KEYINPUT37), .B(G101), .ZN(n1369) );
NAND2_X1 U1060 ( .A1(KEYINPUT36), .A2(n1371), .ZN(n1364) );
NAND2_X1 U1061 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
OR3_X1 U1062 ( .A1(n1189), .A2(G101), .A3(KEYINPUT37), .ZN(n1373) );
INV_X1 U1063 ( .A(n1370), .ZN(n1189) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1374), .ZN(n1370) );
NAND2_X1 U1065 ( .A1(KEYINPUT37), .A2(G101), .ZN(n1372) );
AND2_X1 U1066 ( .A1(n1105), .A2(n1229), .ZN(n1096) );
NOR2_X1 U1067 ( .A1(n1102), .A2(n1103), .ZN(n1229) );
INV_X1 U1068 ( .A(n1311), .ZN(n1103) );
NAND2_X1 U1069 ( .A1(G221), .A2(n1375), .ZN(n1311) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1222), .ZN(n1375) );
XNOR2_X1 U1071 ( .A(n1129), .B(G469), .ZN(n1102) );
AND2_X1 U1072 ( .A1(n1376), .A2(n1222), .ZN(n1129) );
XOR2_X1 U1073 ( .A(n1377), .B(n1378), .Z(n1376) );
XNOR2_X1 U1074 ( .A(n1379), .B(n1380), .ZN(n1378) );
INV_X1 U1075 ( .A(n1206), .ZN(n1380) );
XOR2_X1 U1076 ( .A(n1142), .B(n1381), .Z(n1206) );
XOR2_X1 U1077 ( .A(n1202), .B(n1329), .Z(n1381) );
XNOR2_X1 U1078 ( .A(G101), .B(n1382), .ZN(n1329) );
XNOR2_X1 U1079 ( .A(n1383), .B(G104), .ZN(n1382) );
NAND2_X1 U1080 ( .A1(n1384), .A2(n1385), .ZN(n1202) );
OR2_X1 U1081 ( .A1(n1386), .A2(n1146), .ZN(n1385) );
XOR2_X1 U1082 ( .A(n1387), .B(KEYINPUT28), .Z(n1384) );
NAND2_X1 U1083 ( .A1(n1386), .A2(n1146), .ZN(n1387) );
INV_X1 U1084 ( .A(G131), .ZN(n1146) );
XOR2_X1 U1085 ( .A(G137), .B(n1388), .Z(n1386) );
NOR2_X1 U1086 ( .A1(G134), .A2(KEYINPUT29), .ZN(n1388) );
XOR2_X1 U1087 ( .A(G128), .B(n1389), .Z(n1142) );
NOR2_X1 U1088 ( .A1(KEYINPUT49), .A2(n1363), .ZN(n1389) );
NAND4_X1 U1089 ( .A1(n1213), .A2(n1390), .A3(n1391), .A4(n1392), .ZN(n1379) );
NAND2_X1 U1090 ( .A1(n1212), .A2(n1393), .ZN(n1392) );
AND2_X1 U1091 ( .A1(n1394), .A2(n1346), .ZN(n1212) );
OR2_X1 U1092 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
XOR2_X1 U1093 ( .A(n1395), .B(n1396), .Z(n1394) );
INV_X1 U1094 ( .A(KEYINPUT0), .ZN(n1393) );
INV_X1 U1095 ( .A(n1210), .ZN(n1390) );
NOR3_X1 U1096 ( .A1(n1346), .A2(n1396), .A3(n1395), .ZN(n1210) );
INV_X1 U1097 ( .A(n1322), .ZN(n1346) );
NAND3_X1 U1098 ( .A1(n1322), .A2(n1395), .A3(n1396), .ZN(n1213) );
XNOR2_X1 U1099 ( .A(G140), .B(KEYINPUT26), .ZN(n1396) );
NAND2_X1 U1100 ( .A1(G227), .A2(n1153), .ZN(n1395) );
INV_X1 U1101 ( .A(G953), .ZN(n1153) );
XNOR2_X1 U1102 ( .A(G110), .B(KEYINPUT53), .ZN(n1322) );
XNOR2_X1 U1103 ( .A(KEYINPUT32), .B(KEYINPUT18), .ZN(n1377) );
INV_X1 U1104 ( .A(n1115), .ZN(n1105) );
NAND2_X1 U1105 ( .A1(n1246), .A2(n1247), .ZN(n1115) );
XOR2_X1 U1106 ( .A(n1117), .B(KEYINPUT63), .Z(n1247) );
XOR2_X1 U1107 ( .A(n1397), .B(G475), .Z(n1117) );
NAND2_X1 U1108 ( .A1(n1183), .A2(n1222), .ZN(n1397) );
XNOR2_X1 U1109 ( .A(n1398), .B(n1399), .ZN(n1183) );
XNOR2_X1 U1110 ( .A(n1363), .B(n1141), .ZN(n1399) );
XOR2_X1 U1111 ( .A(G140), .B(n1321), .Z(n1141) );
XOR2_X1 U1112 ( .A(G125), .B(KEYINPUT22), .Z(n1321) );
XNOR2_X1 U1113 ( .A(G143), .B(G146), .ZN(n1363) );
XOR2_X1 U1114 ( .A(n1400), .B(n1401), .Z(n1398) );
XNOR2_X1 U1115 ( .A(G131), .B(n1402), .ZN(n1401) );
NAND2_X1 U1116 ( .A1(n1403), .A2(KEYINPUT59), .ZN(n1402) );
XNOR2_X1 U1117 ( .A(G104), .B(n1404), .ZN(n1403) );
XNOR2_X1 U1118 ( .A(G122), .B(n1309), .ZN(n1404) );
INV_X1 U1119 ( .A(G113), .ZN(n1309) );
NAND2_X1 U1120 ( .A1(G214), .A2(n1374), .ZN(n1400) );
NOR2_X1 U1121 ( .A1(G953), .A2(G237), .ZN(n1374) );
INV_X1 U1122 ( .A(n1123), .ZN(n1246) );
XNOR2_X1 U1123 ( .A(n1405), .B(G478), .ZN(n1123) );
NAND2_X1 U1124 ( .A1(n1179), .A2(n1222), .ZN(n1405) );
INV_X1 U1125 ( .A(G902), .ZN(n1222) );
XNOR2_X1 U1126 ( .A(n1406), .B(n1407), .ZN(n1179) );
XNOR2_X1 U1127 ( .A(n1343), .B(n1408), .ZN(n1407) );
XOR2_X1 U1128 ( .A(G143), .B(G134), .Z(n1408) );
INV_X1 U1129 ( .A(G128), .ZN(n1343) );
XOR2_X1 U1130 ( .A(n1409), .B(n1410), .Z(n1406) );
AND2_X1 U1131 ( .A1(n1347), .A2(G217), .ZN(n1410) );
NOR2_X1 U1132 ( .A1(n1336), .A2(G953), .ZN(n1347) );
INV_X1 U1133 ( .A(G234), .ZN(n1336) );
NAND3_X1 U1134 ( .A1(n1411), .A2(n1412), .A3(KEYINPUT34), .ZN(n1409) );
NAND2_X1 U1135 ( .A1(n1413), .A2(n1383), .ZN(n1412) );
INV_X1 U1136 ( .A(G107), .ZN(n1383) );
NAND2_X1 U1137 ( .A1(n1414), .A2(n1415), .ZN(n1413) );
NAND2_X1 U1138 ( .A1(KEYINPUT52), .A2(n1416), .ZN(n1415) );
NAND3_X1 U1139 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1411) );
INV_X1 U1140 ( .A(KEYINPUT52), .ZN(n1419) );
NAND2_X1 U1141 ( .A1(n1414), .A2(n1420), .ZN(n1418) );
NAND2_X1 U1142 ( .A1(G107), .A2(n1416), .ZN(n1420) );
INV_X1 U1143 ( .A(KEYINPUT5), .ZN(n1416) );
OR2_X1 U1144 ( .A1(n1414), .A2(KEYINPUT5), .ZN(n1417) );
XNOR2_X1 U1145 ( .A(n1306), .B(G122), .ZN(n1414) );
INV_X1 U1146 ( .A(G116), .ZN(n1306) );
endmodule


