//Key = 0110001100101000100110100101001111000000111100111100011001111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XOR2_X1 U741 ( .A(n1022), .B(n1023), .Z(G9) );
NOR2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U743 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND3_X1 U744 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1026) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND4_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NOR3_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U750 ( .A1(KEYINPUT56), .A2(n1045), .ZN(n1043) );
NOR2_X1 U751 ( .A1(KEYINPUT56), .A2(n1046), .ZN(n1040) );
NAND3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1047) );
NAND3_X1 U754 ( .A1(n1037), .A2(n1052), .A3(n1036), .ZN(n1051) );
NAND2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1055), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1036), .A2(n1058), .ZN(n1057) );
OR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1037), .A2(n1061), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U763 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1024) );
INV_X1 U764 ( .A(n1029), .ZN(n1066) );
NAND4_X1 U765 ( .A1(n1067), .A2(n1049), .A3(n1068), .A4(n1069), .ZN(n1029) );
NOR3_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
XNOR2_X1 U767 ( .A(n1073), .B(n1074), .ZN(n1072) );
NAND2_X1 U768 ( .A1(KEYINPUT40), .A2(n1075), .ZN(n1073) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND3_X1 U770 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1070) );
NOR3_X1 U771 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1068) );
NOR3_X1 U772 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
AND2_X1 U773 ( .A1(n1084), .A2(n1086), .ZN(n1082) );
INV_X1 U774 ( .A(KEYINPUT1), .ZN(n1084) );
XOR2_X1 U775 ( .A(G478), .B(n1087), .Z(n1081) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U778 ( .A1(G953), .A2(n1092), .ZN(n1091) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1092) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U781 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1093) );
XNOR2_X1 U783 ( .A(n1098), .B(n1099), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1096) );
XOR2_X1 U785 ( .A(n1102), .B(G140), .Z(n1101) );
NAND2_X1 U786 ( .A1(KEYINPUT58), .A2(G131), .ZN(n1102) );
NAND2_X1 U787 ( .A1(KEYINPUT42), .A2(n1103), .ZN(n1100) );
AND2_X1 U788 ( .A1(n1028), .A2(n1030), .ZN(n1088) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND3_X1 U790 ( .A1(n1106), .A2(n1107), .A3(G953), .ZN(n1105) );
XOR2_X1 U791 ( .A(n1108), .B(KEYINPUT38), .Z(n1104) );
NAND2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U793 ( .A1(G953), .A2(n1111), .ZN(n1110) );
OR2_X1 U794 ( .A1(n1107), .A2(n1106), .ZN(n1111) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1106) );
XNOR2_X1 U796 ( .A(n1027), .B(n1107), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U798 ( .A1(n1114), .A2(G953), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1112) );
XOR2_X1 U800 ( .A(n1117), .B(G122), .Z(n1116) );
NAND3_X1 U801 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
OR3_X1 U803 ( .A1(n1122), .A2(n1121), .A3(n1123), .ZN(n1119) );
INV_X1 U804 ( .A(KEYINPUT32), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(n1118) );
NAND2_X1 U806 ( .A1(n1125), .A2(KEYINPUT32), .ZN(n1124) );
XOR2_X1 U807 ( .A(n1121), .B(KEYINPUT53), .Z(n1125) );
XOR2_X1 U808 ( .A(n1126), .B(KEYINPUT16), .Z(n1121) );
XNOR2_X1 U809 ( .A(n1127), .B(G104), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR3_X1 U812 ( .A1(n1132), .A2(KEYINPUT13), .A3(n1086), .ZN(n1131) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1133), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1087), .A2(n1134), .A3(n1135), .ZN(n1133) );
NOR3_X1 U815 ( .A1(n1136), .A2(n1137), .A3(n1132), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1137), .ZN(n1138) );
INV_X1 U818 ( .A(G478), .ZN(n1137) );
NOR2_X1 U819 ( .A1(n1027), .A2(n1028), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1128), .A2(n1141), .ZN(G60) );
XOR2_X1 U821 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U822 ( .A1(n1077), .A2(n1132), .ZN(n1143) );
NAND2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(G6) );
NAND4_X1 U824 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
INV_X1 U825 ( .A(KEYINPUT44), .ZN(n1149) );
XOR2_X1 U826 ( .A(KEYINPUT12), .B(G104), .Z(n1148) );
NAND2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1151) );
NAND2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NAND2_X1 U830 ( .A1(KEYINPUT44), .A2(KEYINPUT12), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1128), .A2(n1154), .ZN(G57) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U833 ( .A(n1126), .B(n1157), .Z(n1156) );
XOR2_X1 U834 ( .A(n1158), .B(n1159), .Z(n1155) );
XOR2_X1 U835 ( .A(n1160), .B(n1161), .Z(n1158) );
NOR2_X1 U836 ( .A1(n1162), .A2(n1132), .ZN(n1161) );
INV_X1 U837 ( .A(G472), .ZN(n1162) );
NAND2_X1 U838 ( .A1(KEYINPUT63), .A2(n1163), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1128), .A2(n1164), .ZN(G54) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U841 ( .A(n1167), .B(n1168), .ZN(n1166) );
XOR2_X1 U842 ( .A(n1169), .B(n1170), .Z(n1165) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1132), .ZN(n1170) );
INV_X1 U844 ( .A(G469), .ZN(n1171) );
XOR2_X1 U845 ( .A(n1172), .B(KEYINPUT60), .Z(n1169) );
NOR2_X1 U846 ( .A1(n1128), .A2(n1173), .ZN(G51) );
XOR2_X1 U847 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U848 ( .A1(n1074), .A2(n1132), .ZN(n1175) );
NAND2_X1 U849 ( .A1(G902), .A2(n1176), .ZN(n1132) );
OR2_X1 U850 ( .A1(n1028), .A2(n1027), .ZN(n1176) );
NAND4_X1 U851 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1023), .ZN(n1027) );
NAND3_X1 U852 ( .A1(n1180), .A2(n1147), .A3(n1181), .ZN(n1023) );
NAND3_X1 U853 ( .A1(n1147), .A2(n1182), .A3(n1183), .ZN(n1178) );
XOR2_X1 U854 ( .A(n1053), .B(KEYINPUT10), .Z(n1183) );
XOR2_X1 U855 ( .A(KEYINPUT17), .B(n1180), .Z(n1182) );
AND2_X1 U856 ( .A1(n1184), .A2(n1037), .ZN(n1147) );
NAND2_X1 U857 ( .A1(n1180), .A2(n1185), .ZN(n1177) );
NAND4_X1 U858 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
AND2_X1 U859 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NAND3_X1 U860 ( .A1(n1059), .A2(n1192), .A3(n1193), .ZN(n1186) );
NAND4_X1 U861 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1028) );
NOR4_X1 U862 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
INV_X1 U863 ( .A(n1202), .ZN(n1201) );
NAND2_X1 U864 ( .A1(n1146), .A2(n1203), .ZN(n1196) );
NAND2_X1 U865 ( .A1(n1059), .A2(n1204), .ZN(n1194) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND4_X1 U867 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
INV_X1 U868 ( .A(KEYINPUT33), .ZN(n1210) );
INV_X1 U869 ( .A(n1211), .ZN(n1207) );
NAND2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1205) );
NAND2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U872 ( .A1(n1181), .A2(n1216), .ZN(n1215) );
XOR2_X1 U873 ( .A(KEYINPUT4), .B(n1036), .Z(n1216) );
NAND2_X1 U874 ( .A1(KEYINPUT33), .A2(n1208), .ZN(n1214) );
NOR2_X1 U875 ( .A1(n1217), .A2(n1218), .ZN(n1174) );
XOR2_X1 U876 ( .A(KEYINPUT28), .B(n1219), .Z(n1218) );
NOR2_X1 U877 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
AND2_X1 U878 ( .A1(n1221), .A2(n1220), .ZN(n1217) );
XNOR2_X1 U879 ( .A(n1222), .B(n1159), .ZN(n1221) );
XOR2_X1 U880 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U881 ( .A1(G125), .A2(KEYINPUT8), .ZN(n1224) );
NOR2_X1 U882 ( .A1(n1030), .A2(G952), .ZN(n1128) );
XOR2_X1 U883 ( .A(n1225), .B(n1226), .Z(G48) );
NOR2_X1 U884 ( .A1(KEYINPUT51), .A2(n1227), .ZN(n1226) );
NOR3_X1 U885 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1225) );
XOR2_X1 U886 ( .A(n1062), .B(KEYINPUT29), .Z(n1230) );
XOR2_X1 U887 ( .A(n1053), .B(KEYINPUT37), .Z(n1229) );
XOR2_X1 U888 ( .A(n1231), .B(n1195), .Z(G45) );
NAND4_X1 U889 ( .A1(n1232), .A2(n1212), .A3(n1233), .A4(n1234), .ZN(n1195) );
XOR2_X1 U890 ( .A(n1235), .B(n1200), .Z(G42) );
AND3_X1 U891 ( .A1(n1060), .A2(n1212), .A3(n1208), .ZN(n1200) );
AND2_X1 U892 ( .A1(n1192), .A2(n1036), .ZN(n1208) );
NAND2_X1 U893 ( .A1(KEYINPUT22), .A2(n1236), .ZN(n1235) );
INV_X1 U894 ( .A(G140), .ZN(n1236) );
XOR2_X1 U895 ( .A(n1199), .B(n1237), .Z(G39) );
NOR2_X1 U896 ( .A1(KEYINPUT21), .A2(n1238), .ZN(n1237) );
INV_X1 U897 ( .A(G137), .ZN(n1238) );
AND3_X1 U898 ( .A1(n1036), .A2(n1203), .A3(n1038), .ZN(n1199) );
INV_X1 U899 ( .A(n1228), .ZN(n1203) );
XOR2_X1 U900 ( .A(G134), .B(n1239), .Z(G36) );
NOR2_X1 U901 ( .A1(n1054), .A2(n1240), .ZN(n1239) );
XOR2_X1 U902 ( .A(G131), .B(n1241), .Z(G33) );
NOR2_X1 U903 ( .A1(n1053), .A2(n1240), .ZN(n1241) );
NAND3_X1 U904 ( .A1(n1036), .A2(n1212), .A3(n1059), .ZN(n1240) );
AND2_X1 U905 ( .A1(n1065), .A2(n1242), .ZN(n1036) );
XOR2_X1 U906 ( .A(G128), .B(n1198), .Z(G30) );
NOR3_X1 U907 ( .A1(n1054), .A2(n1062), .A3(n1228), .ZN(n1198) );
NAND3_X1 U908 ( .A1(n1243), .A2(n1244), .A3(n1212), .ZN(n1228) );
AND2_X1 U909 ( .A1(n1209), .A2(n1211), .ZN(n1212) );
INV_X1 U910 ( .A(n1181), .ZN(n1054) );
XNOR2_X1 U911 ( .A(G101), .B(n1179), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1038), .A2(n1184), .A3(n1232), .ZN(n1179) );
XOR2_X1 U913 ( .A(n1103), .B(n1202), .Z(G27) );
NAND4_X1 U914 ( .A1(n1146), .A2(n1060), .A3(n1049), .A4(n1211), .ZN(n1202) );
NAND2_X1 U915 ( .A1(n1245), .A2(n1246), .ZN(n1211) );
NAND2_X1 U916 ( .A1(n1247), .A2(n1095), .ZN(n1246) );
INV_X1 U917 ( .A(G900), .ZN(n1095) );
NOR2_X1 U918 ( .A1(n1053), .A2(n1062), .ZN(n1146) );
XOR2_X1 U919 ( .A(G122), .B(n1248), .Z(G24) );
NOR3_X1 U920 ( .A1(n1190), .A2(KEYINPUT55), .A3(n1249), .ZN(n1248) );
XOR2_X1 U921 ( .A(n1062), .B(KEYINPUT3), .Z(n1249) );
NAND4_X1 U922 ( .A1(n1193), .A2(n1037), .A3(n1233), .A4(n1234), .ZN(n1190) );
NOR2_X1 U923 ( .A1(n1244), .A2(n1243), .ZN(n1037) );
XNOR2_X1 U924 ( .A(G119), .B(n1250), .ZN(G21) );
NAND2_X1 U925 ( .A1(n1251), .A2(n1180), .ZN(n1250) );
XOR2_X1 U926 ( .A(n1187), .B(KEYINPUT61), .Z(n1251) );
NAND4_X1 U927 ( .A1(n1193), .A2(n1038), .A3(n1243), .A4(n1244), .ZN(n1187) );
INV_X1 U928 ( .A(n1067), .ZN(n1243) );
XOR2_X1 U929 ( .A(G116), .B(n1252), .Z(G18) );
NOR2_X1 U930 ( .A1(n1253), .A2(n1062), .ZN(n1252) );
XOR2_X1 U931 ( .A(n1189), .B(KEYINPUT50), .Z(n1253) );
NAND3_X1 U932 ( .A1(n1059), .A2(n1181), .A3(n1193), .ZN(n1189) );
NOR2_X1 U933 ( .A1(n1234), .A2(n1254), .ZN(n1181) );
XOR2_X1 U934 ( .A(n1255), .B(n1256), .Z(G15) );
NAND4_X1 U935 ( .A1(KEYINPUT25), .A2(n1193), .A3(n1232), .A4(n1192), .ZN(n1256) );
INV_X1 U936 ( .A(n1053), .ZN(n1192) );
NAND2_X1 U937 ( .A1(n1254), .A2(n1234), .ZN(n1053) );
INV_X1 U938 ( .A(n1233), .ZN(n1254) );
AND2_X1 U939 ( .A1(n1059), .A2(n1180), .ZN(n1232) );
NOR2_X1 U940 ( .A1(n1244), .A2(n1067), .ZN(n1059) );
AND2_X1 U941 ( .A1(n1049), .A2(n1257), .ZN(n1193) );
INV_X1 U942 ( .A(n1046), .ZN(n1049) );
NAND2_X1 U943 ( .A1(n1258), .A2(n1044), .ZN(n1046) );
INV_X1 U944 ( .A(n1045), .ZN(n1258) );
XOR2_X1 U945 ( .A(n1259), .B(n1260), .Z(G12) );
NAND3_X1 U946 ( .A1(KEYINPUT6), .A2(n1180), .A3(n1261), .ZN(n1260) );
XOR2_X1 U947 ( .A(n1191), .B(KEYINPUT19), .Z(n1261) );
NAND3_X1 U948 ( .A1(n1038), .A2(n1184), .A3(n1060), .ZN(n1191) );
AND2_X1 U949 ( .A1(n1067), .A2(n1244), .ZN(n1060) );
NAND2_X1 U950 ( .A1(n1078), .A2(n1262), .ZN(n1244) );
OR2_X1 U951 ( .A1(n1086), .A2(n1085), .ZN(n1262) );
NAND2_X1 U952 ( .A1(n1085), .A2(n1086), .ZN(n1078) );
NAND2_X1 U953 ( .A1(G217), .A2(n1263), .ZN(n1086) );
NOR2_X1 U954 ( .A1(n1130), .A2(G902), .ZN(n1085) );
XOR2_X1 U955 ( .A(n1264), .B(n1265), .Z(n1130) );
XOR2_X1 U956 ( .A(n1266), .B(n1267), .Z(n1265) );
NAND3_X1 U957 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
OR2_X1 U958 ( .A1(n1259), .A2(KEYINPUT7), .ZN(n1270) );
NAND3_X1 U959 ( .A1(KEYINPUT7), .A2(n1271), .A3(n1272), .ZN(n1269) );
OR2_X1 U960 ( .A1(n1272), .A2(n1271), .ZN(n1268) );
NOR2_X1 U961 ( .A1(G110), .A2(KEYINPUT5), .ZN(n1271) );
XOR2_X1 U962 ( .A(G119), .B(G128), .Z(n1272) );
NAND2_X1 U963 ( .A1(n1273), .A2(KEYINPUT2), .ZN(n1266) );
XOR2_X1 U964 ( .A(n1274), .B(G137), .Z(n1273) );
NAND2_X1 U965 ( .A1(G221), .A2(n1275), .ZN(n1274) );
XOR2_X1 U966 ( .A(n1276), .B(G472), .Z(n1067) );
NAND2_X1 U967 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U968 ( .A(n1279), .B(n1280), .Z(n1277) );
XNOR2_X1 U969 ( .A(n1281), .B(n1282), .ZN(n1280) );
NOR2_X1 U970 ( .A1(KEYINPUT11), .A2(n1126), .ZN(n1282) );
NAND2_X1 U971 ( .A1(KEYINPUT47), .A2(n1283), .ZN(n1281) );
XOR2_X1 U972 ( .A(n1157), .B(n1163), .Z(n1279) );
XOR2_X1 U973 ( .A(n1284), .B(G101), .Z(n1157) );
NAND2_X1 U974 ( .A1(G210), .A2(n1285), .ZN(n1284) );
AND2_X1 U975 ( .A1(n1209), .A2(n1257), .ZN(n1184) );
NAND2_X1 U976 ( .A1(n1245), .A2(n1286), .ZN(n1257) );
NAND2_X1 U977 ( .A1(n1247), .A2(n1114), .ZN(n1286) );
XNOR2_X1 U978 ( .A(G898), .B(KEYINPUT24), .ZN(n1114) );
NOR3_X1 U979 ( .A1(n1278), .A2(n1041), .A3(n1030), .ZN(n1247) );
INV_X1 U980 ( .A(n1048), .ZN(n1041) );
NAND3_X1 U981 ( .A1(n1048), .A2(n1030), .A3(n1287), .ZN(n1245) );
XOR2_X1 U982 ( .A(n1032), .B(KEYINPUT39), .Z(n1287) );
XNOR2_X1 U983 ( .A(G952), .B(KEYINPUT46), .ZN(n1032) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1048) );
AND2_X1 U985 ( .A1(n1045), .A2(n1044), .ZN(n1209) );
NAND2_X1 U986 ( .A1(G221), .A2(n1263), .ZN(n1044) );
NAND2_X1 U987 ( .A1(G234), .A2(n1278), .ZN(n1263) );
XNOR2_X1 U988 ( .A(n1288), .B(G469), .ZN(n1045) );
NAND2_X1 U989 ( .A1(n1289), .A2(n1278), .ZN(n1288) );
XOR2_X1 U990 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U991 ( .A(n1292), .B(n1167), .Z(n1291) );
XOR2_X1 U992 ( .A(n1293), .B(n1163), .Z(n1167) );
XNOR2_X1 U993 ( .A(n1294), .B(n1098), .ZN(n1163) );
XOR2_X1 U994 ( .A(G134), .B(G137), .Z(n1098) );
XNOR2_X1 U995 ( .A(G131), .B(KEYINPUT23), .ZN(n1294) );
XOR2_X1 U996 ( .A(n1259), .B(G140), .Z(n1293) );
NAND2_X1 U997 ( .A1(KEYINPUT41), .A2(n1168), .ZN(n1292) );
XOR2_X1 U998 ( .A(n1099), .B(n1295), .Z(n1168) );
XOR2_X1 U999 ( .A(G101), .B(n1296), .Z(n1295) );
NOR2_X1 U1000 ( .A1(KEYINPUT52), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1001 ( .A(n1153), .B(n1298), .Z(n1297) );
NOR2_X1 U1002 ( .A1(KEYINPUT18), .A2(n1022), .ZN(n1298) );
INV_X1 U1003 ( .A(G107), .ZN(n1022) );
XOR2_X1 U1004 ( .A(n1299), .B(n1300), .Z(n1099) );
XNOR2_X1 U1005 ( .A(n1301), .B(KEYINPUT30), .ZN(n1300) );
NAND2_X1 U1006 ( .A1(KEYINPUT27), .A2(n1231), .ZN(n1301) );
XOR2_X1 U1007 ( .A(n1172), .B(n1302), .Z(n1290) );
XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(KEYINPUT35), .ZN(n1302) );
NAND2_X1 U1009 ( .A1(G227), .A2(n1030), .ZN(n1172) );
NOR2_X1 U1010 ( .A1(n1234), .A2(n1233), .ZN(n1038) );
XNOR2_X1 U1011 ( .A(n1087), .B(n1303), .ZN(n1233) );
NOR2_X1 U1012 ( .A1(G478), .A2(KEYINPUT0), .ZN(n1303) );
NOR2_X1 U1013 ( .A1(n1139), .A2(G902), .ZN(n1087) );
INV_X1 U1014 ( .A(n1136), .ZN(n1139) );
XOR2_X1 U1015 ( .A(n1304), .B(n1305), .Z(n1136) );
XOR2_X1 U1016 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1017 ( .A(G128), .B(G122), .Z(n1307) );
XOR2_X1 U1018 ( .A(KEYINPUT14), .B(G143), .Z(n1306) );
XOR2_X1 U1019 ( .A(n1308), .B(n1309), .Z(n1304) );
XOR2_X1 U1020 ( .A(G116), .B(G107), .Z(n1309) );
XOR2_X1 U1021 ( .A(n1310), .B(n1311), .Z(n1308) );
NOR2_X1 U1022 ( .A1(KEYINPUT15), .A2(G134), .ZN(n1311) );
NAND2_X1 U1023 ( .A1(G217), .A2(n1275), .ZN(n1310) );
AND2_X1 U1024 ( .A1(G234), .A2(n1030), .ZN(n1275) );
NAND3_X1 U1025 ( .A1(n1312), .A2(n1313), .A3(n1079), .ZN(n1234) );
NAND2_X1 U1026 ( .A1(n1076), .A2(n1077), .ZN(n1079) );
NAND2_X1 U1027 ( .A1(KEYINPUT45), .A2(n1077), .ZN(n1313) );
OR3_X1 U1028 ( .A1(n1076), .A2(KEYINPUT45), .A3(n1077), .ZN(n1312) );
INV_X1 U1029 ( .A(G475), .ZN(n1077) );
NOR2_X1 U1030 ( .A1(n1142), .A2(G902), .ZN(n1076) );
XOR2_X1 U1031 ( .A(n1314), .B(n1315), .Z(n1142) );
XOR2_X1 U1032 ( .A(G113), .B(n1316), .Z(n1315) );
NOR2_X1 U1033 ( .A1(KEYINPUT26), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1034 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1035 ( .A(KEYINPUT36), .B(G143), .Z(n1319) );
XOR2_X1 U1036 ( .A(n1320), .B(G131), .Z(n1318) );
NAND3_X1 U1037 ( .A1(G214), .A2(n1285), .A3(KEYINPUT31), .ZN(n1320) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1285) );
XOR2_X1 U1039 ( .A(n1264), .B(n1321), .Z(n1314) );
XOR2_X1 U1040 ( .A(n1103), .B(n1322), .Z(n1264) );
XOR2_X1 U1041 ( .A(G146), .B(G140), .Z(n1322) );
INV_X1 U1042 ( .A(G125), .ZN(n1103) );
INV_X1 U1043 ( .A(n1062), .ZN(n1180) );
NAND2_X1 U1044 ( .A1(n1323), .A2(n1242), .ZN(n1062) );
XOR2_X1 U1045 ( .A(n1064), .B(KEYINPUT57), .Z(n1242) );
INV_X1 U1046 ( .A(n1080), .ZN(n1064) );
NAND2_X1 U1047 ( .A1(G214), .A2(n1324), .ZN(n1080) );
XOR2_X1 U1048 ( .A(KEYINPUT20), .B(n1065), .Z(n1323) );
XOR2_X1 U1049 ( .A(n1325), .B(n1075), .Z(n1065) );
NAND3_X1 U1050 ( .A1(n1326), .A2(n1278), .A3(n1327), .ZN(n1075) );
NAND2_X1 U1051 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1052 ( .A(n1283), .B(G125), .Z(n1328) );
INV_X1 U1053 ( .A(n1159), .ZN(n1283) );
NAND2_X1 U1054 ( .A1(n1330), .A2(n1331), .ZN(n1326) );
XOR2_X1 U1055 ( .A(KEYINPUT59), .B(n1329), .Z(n1331) );
XOR2_X1 U1056 ( .A(n1220), .B(n1223), .Z(n1329) );
NAND2_X1 U1057 ( .A1(G224), .A2(n1030), .ZN(n1223) );
INV_X1 U1058 ( .A(G953), .ZN(n1030) );
XOR2_X1 U1059 ( .A(n1332), .B(n1333), .Z(n1220) );
XNOR2_X1 U1060 ( .A(n1127), .B(n1321), .ZN(n1333) );
XNOR2_X1 U1061 ( .A(n1153), .B(G122), .ZN(n1321) );
INV_X1 U1062 ( .A(G104), .ZN(n1153) );
XOR2_X1 U1063 ( .A(n1334), .B(n1335), .Z(n1127) );
XOR2_X1 U1064 ( .A(G107), .B(G101), .Z(n1335) );
XNOR2_X1 U1065 ( .A(KEYINPUT9), .B(KEYINPUT34), .ZN(n1334) );
XNOR2_X1 U1066 ( .A(n1126), .B(n1117), .ZN(n1332) );
NAND2_X1 U1067 ( .A1(KEYINPUT48), .A2(n1259), .ZN(n1117) );
XOR2_X1 U1068 ( .A(n1255), .B(n1336), .Z(n1126) );
XOR2_X1 U1069 ( .A(G119), .B(G116), .Z(n1336) );
INV_X1 U1070 ( .A(G113), .ZN(n1255) );
XOR2_X1 U1071 ( .A(G125), .B(n1159), .Z(n1330) );
XNOR2_X1 U1072 ( .A(n1231), .B(n1337), .ZN(n1159) );
INV_X1 U1073 ( .A(n1299), .ZN(n1337) );
XOR2_X1 U1074 ( .A(n1227), .B(G128), .Z(n1299) );
INV_X1 U1075 ( .A(G146), .ZN(n1227) );
INV_X1 U1076 ( .A(G143), .ZN(n1231) );
NAND2_X1 U1077 ( .A1(KEYINPUT54), .A2(n1074), .ZN(n1325) );
NAND2_X1 U1078 ( .A1(G210), .A2(n1324), .ZN(n1074) );
NAND2_X1 U1079 ( .A1(n1338), .A2(n1278), .ZN(n1324) );
INV_X1 U1080 ( .A(G902), .ZN(n1278) );
XOR2_X1 U1081 ( .A(n1339), .B(G237), .Z(n1338) );
XNOR2_X1 U1082 ( .A(KEYINPUT62), .B(KEYINPUT43), .ZN(n1339) );
INV_X1 U1083 ( .A(G110), .ZN(n1259) );
endmodule


