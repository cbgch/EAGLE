//Key = 1100001010000110000001110100001001110101101011000111001111100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312;

XOR2_X1 U713 ( .A(n986), .B(n987), .Z(G9) );
NOR2_X1 U714 ( .A1(KEYINPUT28), .A2(n988), .ZN(n987) );
NOR2_X1 U715 ( .A1(n989), .A2(n990), .ZN(G75) );
NOR4_X1 U716 ( .A1(G953), .A2(n991), .A3(n992), .A4(n993), .ZN(n990) );
NOR2_X1 U717 ( .A1(n994), .A2(n995), .ZN(n992) );
INV_X1 U718 ( .A(n996), .ZN(n995) );
NOR2_X1 U719 ( .A1(n997), .A2(n998), .ZN(n994) );
NOR3_X1 U720 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NOR4_X1 U721 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
NOR2_X1 U722 ( .A1(KEYINPUT24), .A2(n1006), .ZN(n1005) );
NOR2_X1 U723 ( .A1(n1007), .A2(n1008), .ZN(n1003) );
NOR2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U725 ( .A1(n1011), .A2(n1012), .ZN(n1000) );
AND2_X1 U726 ( .A1(n1013), .A2(KEYINPUT24), .ZN(n1012) );
NOR4_X1 U727 ( .A1(n1014), .A2(n1015), .A3(n1008), .A4(n1016), .ZN(n997) );
NOR3_X1 U728 ( .A1(n1002), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR2_X1 U729 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1021), .ZN(n1014) );
NOR2_X1 U731 ( .A1(n1022), .A2(n999), .ZN(n1021) );
INV_X1 U732 ( .A(n1023), .ZN(n999) );
NOR2_X1 U733 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U734 ( .A1(n991), .A2(G953), .A3(G952), .ZN(n989) );
AND4_X1 U735 ( .A1(n1026), .A2(n1025), .A3(n1027), .A4(n1028), .ZN(n991) );
NOR3_X1 U736 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
XNOR2_X1 U737 ( .A(n1032), .B(n1033), .ZN(n1031) );
XNOR2_X1 U738 ( .A(G475), .B(n1034), .ZN(n1030) );
NAND3_X1 U739 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1029) );
XOR2_X1 U740 ( .A(KEYINPUT0), .B(n1038), .Z(n1036) );
NOR2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
XNOR2_X1 U742 ( .A(KEYINPUT38), .B(n1041), .ZN(n1040) );
NOR3_X1 U743 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1027) );
INV_X1 U744 ( .A(n1045), .ZN(n1044) );
XOR2_X1 U745 ( .A(KEYINPUT14), .B(n1046), .Z(n1026) );
NOR2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND4_X1 U747 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(G72) );
OR2_X1 U748 ( .A1(n1053), .A2(KEYINPUT22), .ZN(n1052) );
NAND3_X1 U749 ( .A1(n1054), .A2(n1053), .A3(KEYINPUT22), .ZN(n1051) );
NAND2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U751 ( .A1(G953), .A2(n1057), .ZN(n1056) );
NAND3_X1 U752 ( .A1(G227), .A2(n1058), .A3(G900), .ZN(n1050) );
NAND2_X1 U753 ( .A1(KEYINPUT22), .A2(n1059), .ZN(n1058) );
OR2_X1 U754 ( .A1(n1053), .A2(n1060), .ZN(n1059) );
NAND2_X1 U755 ( .A1(n1061), .A2(n1060), .ZN(n1049) );
NAND2_X1 U756 ( .A1(n1062), .A2(KEYINPUT22), .ZN(n1061) );
XOR2_X1 U757 ( .A(n1053), .B(n1063), .Z(n1062) );
NOR2_X1 U758 ( .A1(n1064), .A2(KEYINPUT16), .ZN(n1063) );
NOR2_X1 U759 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U760 ( .A1(n1067), .A2(n1055), .ZN(n1053) );
INV_X1 U761 ( .A(n1068), .ZN(n1055) );
XOR2_X1 U762 ( .A(n1069), .B(n1070), .Z(n1067) );
XOR2_X1 U763 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U764 ( .A1(KEYINPUT33), .A2(n1073), .ZN(n1071) );
NAND2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(G69) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1060), .ZN(n1075) );
XOR2_X1 U767 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U768 ( .A1(n1079), .A2(G953), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1082), .ZN(n1081) );
NAND2_X1 U771 ( .A1(G224), .A2(n1083), .ZN(n1080) );
NAND2_X1 U772 ( .A1(G898), .A2(n1077), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1077) );
NAND2_X1 U774 ( .A1(G953), .A2(n1086), .ZN(n1085) );
XOR2_X1 U775 ( .A(n1087), .B(n1088), .Z(n1084) );
XNOR2_X1 U776 ( .A(n1089), .B(KEYINPUT13), .ZN(n1088) );
NAND2_X1 U777 ( .A1(KEYINPUT6), .A2(n1090), .ZN(n1089) );
NOR2_X1 U778 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U780 ( .A(n1095), .B(KEYINPUT12), .Z(n1093) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1047), .ZN(n1095) );
NOR2_X1 U782 ( .A1(n1091), .A2(n1097), .ZN(G63) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U784 ( .A1(n1096), .A2(G478), .A3(KEYINPUT25), .ZN(n1098) );
NOR2_X1 U785 ( .A1(n1091), .A2(n1100), .ZN(G60) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U787 ( .A(KEYINPUT2), .B(n1103), .Z(n1102) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
AND2_X1 U789 ( .A1(n1105), .A2(n1104), .ZN(n1101) );
XNOR2_X1 U790 ( .A(n1106), .B(KEYINPUT1), .ZN(n1104) );
NAND2_X1 U791 ( .A1(n1096), .A2(G475), .ZN(n1105) );
XNOR2_X1 U792 ( .A(n1107), .B(n1108), .ZN(G6) );
NAND2_X1 U793 ( .A1(KEYINPUT57), .A2(G104), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1091), .A2(n1109), .ZN(G57) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(n1109) );
XNOR2_X1 U796 ( .A(n1112), .B(n1113), .ZN(n1111) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR3_X1 U798 ( .A1(n1116), .A2(KEYINPUT29), .A3(n1117), .ZN(n1114) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1110) );
NOR2_X1 U800 ( .A1(KEYINPUT48), .A2(n1120), .ZN(n1119) );
XOR2_X1 U801 ( .A(n1121), .B(KEYINPUT19), .Z(n1118) );
NOR2_X1 U802 ( .A1(n1091), .A2(n1122), .ZN(G54) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U804 ( .A(n1125), .B(n1072), .Z(n1124) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1123) );
NAND2_X1 U806 ( .A1(n1096), .A2(G469), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1091), .A2(n1128), .ZN(G51) );
XOR2_X1 U808 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U809 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND2_X1 U810 ( .A1(n1096), .A2(n1032), .ZN(n1131) );
INV_X1 U811 ( .A(n1116), .ZN(n1096) );
NAND2_X1 U812 ( .A1(G902), .A2(n993), .ZN(n1116) );
NAND3_X1 U813 ( .A1(n1133), .A2(n1134), .A3(n1078), .ZN(n993) );
AND2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1078) );
NOR4_X1 U815 ( .A1(n1137), .A2(n1107), .A3(n986), .A4(n1138), .ZN(n1136) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
AND3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1010), .ZN(n986) );
AND3_X1 U818 ( .A1(n1141), .A2(n1142), .A3(n1009), .ZN(n1107) );
NOR4_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1135) );
XOR2_X1 U820 ( .A(KEYINPUT39), .B(n1065), .Z(n1134) );
INV_X1 U821 ( .A(n1066), .ZN(n1133) );
NAND4_X1 U822 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1066) );
AND3_X1 U823 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NAND2_X1 U824 ( .A1(n1023), .A2(n1154), .ZN(n1149) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U826 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U827 ( .A(KEYINPUT11), .B(n1016), .ZN(n1158) );
XOR2_X1 U828 ( .A(KEYINPUT56), .B(n1159), .Z(n1155) );
NOR2_X1 U829 ( .A1(n1060), .A2(G952), .ZN(n1091) );
XNOR2_X1 U830 ( .A(G146), .B(n1147), .ZN(G48) );
NAND3_X1 U831 ( .A1(n1009), .A2(n1017), .A3(n1157), .ZN(n1147) );
XOR2_X1 U832 ( .A(G143), .B(n1065), .Z(G45) );
AND3_X1 U833 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1065) );
NAND2_X1 U834 ( .A1(n1163), .A2(n1164), .ZN(G42) );
NAND2_X1 U835 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1163) );
NOR2_X1 U837 ( .A1(n1165), .A2(n1166), .ZN(n1168) );
INV_X1 U838 ( .A(KEYINPUT62), .ZN(n1166) );
INV_X1 U839 ( .A(G140), .ZN(n1165) );
NAND2_X1 U840 ( .A1(n1159), .A2(n1023), .ZN(n1167) );
NOR3_X1 U841 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1159) );
INV_X1 U842 ( .A(n1162), .ZN(n1171) );
XNOR2_X1 U843 ( .A(G137), .B(n1172), .ZN(G39) );
NAND3_X1 U844 ( .A1(n1157), .A2(n1173), .A3(n1023), .ZN(n1172) );
XNOR2_X1 U845 ( .A(G134), .B(n1148), .ZN(G36) );
NAND2_X1 U846 ( .A1(n1174), .A2(n1010), .ZN(n1148) );
XNOR2_X1 U847 ( .A(G131), .B(n1151), .ZN(G33) );
NAND2_X1 U848 ( .A1(n1174), .A2(n1009), .ZN(n1151) );
AND3_X1 U849 ( .A1(n1162), .A2(n1160), .A3(n1023), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1019), .A2(n1042), .ZN(n1023) );
INV_X1 U851 ( .A(n1020), .ZN(n1042) );
XNOR2_X1 U852 ( .A(G128), .B(n1153), .ZN(G30) );
NAND3_X1 U853 ( .A1(n1010), .A2(n1017), .A3(n1157), .ZN(n1153) );
AND3_X1 U854 ( .A1(n1175), .A2(n1176), .A3(n1162), .ZN(n1157) );
NOR2_X1 U855 ( .A1(n1177), .A2(n1178), .ZN(n1162) );
INV_X1 U856 ( .A(n1179), .ZN(n1178) );
XOR2_X1 U857 ( .A(G101), .B(n1145), .Z(G3) );
AND2_X1 U858 ( .A1(n1004), .A2(n1141), .ZN(n1145) );
AND2_X1 U859 ( .A1(n1160), .A2(n1173), .ZN(n1004) );
XNOR2_X1 U860 ( .A(G125), .B(n1152), .ZN(G27) );
NAND4_X1 U861 ( .A1(n1017), .A2(n1179), .A3(n1011), .A4(n1180), .ZN(n1152) );
NOR2_X1 U862 ( .A1(n1170), .A2(n1169), .ZN(n1180) );
NAND2_X1 U863 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NAND3_X1 U864 ( .A1(G902), .A2(n996), .A3(n1068), .ZN(n1182) );
NOR2_X1 U865 ( .A1(n1060), .A2(G900), .ZN(n1068) );
XOR2_X1 U866 ( .A(G122), .B(n1137), .Z(G24) );
AND4_X1 U867 ( .A1(n1161), .A2(n1011), .A3(n1142), .A4(n1183), .ZN(n1137) );
INV_X1 U868 ( .A(n1008), .ZN(n1142) );
NAND2_X1 U869 ( .A1(n1184), .A2(n1185), .ZN(n1008) );
AND3_X1 U870 ( .A1(n1017), .A2(n1186), .A3(n1187), .ZN(n1161) );
XOR2_X1 U871 ( .A(n1188), .B(KEYINPUT36), .Z(n1187) );
XNOR2_X1 U872 ( .A(G119), .B(n1189), .ZN(G21) );
NAND2_X1 U873 ( .A1(n1190), .A2(n1017), .ZN(n1189) );
XOR2_X1 U874 ( .A(n1140), .B(KEYINPUT21), .Z(n1190) );
NAND4_X1 U875 ( .A1(n1175), .A2(n1173), .A3(n1191), .A4(n1011), .ZN(n1140) );
NOR2_X1 U876 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U877 ( .A(n1194), .B(n1144), .ZN(G18) );
AND2_X1 U878 ( .A1(n1195), .A2(n1010), .ZN(n1144) );
AND2_X1 U879 ( .A1(n1196), .A2(n1186), .ZN(n1010) );
XNOR2_X1 U880 ( .A(KEYINPUT61), .B(n1188), .ZN(n1196) );
XOR2_X1 U881 ( .A(n1197), .B(n1143), .Z(G15) );
AND2_X1 U882 ( .A1(n1195), .A2(n1009), .ZN(n1143) );
INV_X1 U883 ( .A(n1170), .ZN(n1009) );
NAND2_X1 U884 ( .A1(n1037), .A2(n1188), .ZN(n1170) );
INV_X1 U885 ( .A(n1186), .ZN(n1037) );
AND4_X1 U886 ( .A1(n1160), .A2(n1011), .A3(n1017), .A4(n1183), .ZN(n1195) );
INV_X1 U887 ( .A(n1139), .ZN(n1017) );
INV_X1 U888 ( .A(n1002), .ZN(n1011) );
NAND2_X1 U889 ( .A1(n1024), .A2(n1025), .ZN(n1002) );
INV_X1 U890 ( .A(n1198), .ZN(n1024) );
AND2_X1 U891 ( .A1(n1184), .A2(n1176), .ZN(n1160) );
XNOR2_X1 U892 ( .A(G113), .B(KEYINPUT40), .ZN(n1197) );
XOR2_X1 U893 ( .A(n1199), .B(G110), .Z(G12) );
NAND2_X1 U894 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND4_X1 U895 ( .A1(n1183), .A2(n1139), .A3(n1202), .A4(n1203), .ZN(n1201) );
INV_X1 U896 ( .A(KEYINPUT44), .ZN(n1203) );
NOR2_X1 U897 ( .A1(n1177), .A2(n1006), .ZN(n1202) );
INV_X1 U898 ( .A(n1013), .ZN(n1006) );
NAND2_X1 U899 ( .A1(n1146), .A2(KEYINPUT44), .ZN(n1200) );
AND2_X1 U900 ( .A1(n1013), .A2(n1141), .ZN(n1146) );
NOR3_X1 U901 ( .A1(n1139), .A2(n1192), .A3(n1177), .ZN(n1141) );
NAND2_X1 U902 ( .A1(n1025), .A2(n1198), .ZN(n1177) );
NAND2_X1 U903 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NAND2_X1 U904 ( .A1(n1206), .A2(n1041), .ZN(n1205) );
XNOR2_X1 U905 ( .A(n1043), .B(KEYINPUT9), .ZN(n1204) );
NOR2_X1 U906 ( .A1(n1041), .A2(n1206), .ZN(n1043) );
INV_X1 U907 ( .A(n1039), .ZN(n1206) );
NAND2_X1 U908 ( .A1(n1207), .A2(n1208), .ZN(n1039) );
XOR2_X1 U909 ( .A(n1209), .B(n1210), .Z(n1207) );
XNOR2_X1 U910 ( .A(n1125), .B(n1211), .ZN(n1210) );
NOR2_X1 U911 ( .A1(KEYINPUT7), .A2(n1212), .ZN(n1211) );
XOR2_X1 U912 ( .A(n1213), .B(n1072), .Z(n1212) );
XNOR2_X1 U913 ( .A(n1214), .B(G143), .ZN(n1072) );
NAND2_X1 U914 ( .A1(KEYINPUT30), .A2(G128), .ZN(n1214) );
XNOR2_X1 U915 ( .A(n1215), .B(n1216), .ZN(n1125) );
XOR2_X1 U916 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U917 ( .A1(G953), .A2(n1057), .ZN(n1217) );
INV_X1 U918 ( .A(G227), .ZN(n1057) );
XOR2_X1 U919 ( .A(n1219), .B(G104), .Z(n1215) );
XNOR2_X1 U920 ( .A(G140), .B(KEYINPUT34), .ZN(n1209) );
INV_X1 U921 ( .A(G469), .ZN(n1041) );
NAND2_X1 U922 ( .A1(G221), .A2(n1220), .ZN(n1025) );
INV_X1 U923 ( .A(n1183), .ZN(n1192) );
NAND2_X1 U924 ( .A1(n1181), .A2(n1221), .ZN(n1183) );
NAND4_X1 U925 ( .A1(G953), .A2(G902), .A3(n996), .A4(n1086), .ZN(n1221) );
INV_X1 U926 ( .A(G898), .ZN(n1086) );
NAND3_X1 U927 ( .A1(n996), .A2(n1060), .A3(n1222), .ZN(n1181) );
XOR2_X1 U928 ( .A(KEYINPUT5), .B(G952), .Z(n1222) );
NAND2_X1 U929 ( .A1(G237), .A2(G234), .ZN(n996) );
NAND2_X1 U930 ( .A1(n1019), .A2(n1020), .ZN(n1139) );
NAND2_X1 U931 ( .A1(G214), .A2(n1223), .ZN(n1020) );
XOR2_X1 U932 ( .A(n1033), .B(n1224), .Z(n1019) );
NOR2_X1 U933 ( .A1(n1032), .A2(KEYINPUT60), .ZN(n1224) );
AND2_X1 U934 ( .A1(G210), .A2(n1223), .ZN(n1032) );
NAND2_X1 U935 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
INV_X1 U936 ( .A(G237), .ZN(n1225) );
NAND2_X1 U937 ( .A1(n1227), .A2(n1208), .ZN(n1033) );
XOR2_X1 U938 ( .A(n1129), .B(n1228), .Z(n1227) );
NOR2_X1 U939 ( .A1(KEYINPUT18), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U940 ( .A(n1132), .B(KEYINPUT46), .ZN(n1229) );
NOR2_X1 U941 ( .A1(n1082), .A2(G953), .ZN(n1132) );
INV_X1 U942 ( .A(G224), .ZN(n1082) );
XOR2_X1 U943 ( .A(n1230), .B(n1231), .Z(n1129) );
XNOR2_X1 U944 ( .A(G125), .B(n1090), .ZN(n1231) );
NAND3_X1 U945 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1090) );
OR2_X1 U946 ( .A1(G113), .A2(KEYINPUT55), .ZN(n1234) );
NAND3_X1 U947 ( .A1(KEYINPUT55), .A2(G113), .A3(n1235), .ZN(n1233) );
INV_X1 U948 ( .A(n1236), .ZN(n1235) );
NAND2_X1 U949 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
NAND2_X1 U950 ( .A1(KEYINPUT55), .A2(n1238), .ZN(n1237) );
XOR2_X1 U951 ( .A(KEYINPUT59), .B(G113), .Z(n1238) );
XOR2_X1 U952 ( .A(n1087), .B(n1239), .Z(n1230) );
XOR2_X1 U953 ( .A(n1240), .B(n1241), .Z(n1087) );
XNOR2_X1 U954 ( .A(n1218), .B(KEYINPUT3), .ZN(n1240) );
XOR2_X1 U955 ( .A(n1242), .B(n1243), .Z(n1218) );
XNOR2_X1 U956 ( .A(G107), .B(G110), .ZN(n1242) );
NOR2_X1 U957 ( .A1(n1169), .A2(n1016), .ZN(n1013) );
INV_X1 U958 ( .A(n1173), .ZN(n1016) );
NOR2_X1 U959 ( .A1(n1186), .A2(n1188), .ZN(n1173) );
NAND3_X1 U960 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1188) );
OR2_X1 U961 ( .A1(n1247), .A2(n1034), .ZN(n1246) );
NAND3_X1 U962 ( .A1(n1034), .A2(n1247), .A3(G475), .ZN(n1245) );
NAND2_X1 U963 ( .A1(n1248), .A2(n1249), .ZN(n1244) );
INV_X1 U964 ( .A(G475), .ZN(n1249) );
NAND2_X1 U965 ( .A1(n1250), .A2(n1247), .ZN(n1248) );
INV_X1 U966 ( .A(KEYINPUT4), .ZN(n1247) );
XOR2_X1 U967 ( .A(n1034), .B(KEYINPUT63), .Z(n1250) );
NAND2_X1 U968 ( .A1(n1251), .A2(n1208), .ZN(n1034) );
XOR2_X1 U969 ( .A(n1106), .B(KEYINPUT27), .Z(n1251) );
XOR2_X1 U970 ( .A(n1252), .B(n1253), .Z(n1106) );
XOR2_X1 U971 ( .A(n1069), .B(n1254), .Z(n1253) );
XOR2_X1 U972 ( .A(n1255), .B(n1241), .Z(n1254) );
XOR2_X1 U973 ( .A(G104), .B(G122), .Z(n1241) );
NAND2_X1 U974 ( .A1(G214), .A2(n1256), .ZN(n1255) );
XOR2_X1 U975 ( .A(n1257), .B(G131), .Z(n1069) );
XOR2_X1 U976 ( .A(n1258), .B(n1259), .Z(n1252) );
XOR2_X1 U977 ( .A(G143), .B(G113), .Z(n1259) );
XNOR2_X1 U978 ( .A(KEYINPUT49), .B(KEYINPUT42), .ZN(n1258) );
XNOR2_X1 U979 ( .A(n1260), .B(G478), .ZN(n1186) );
NAND2_X1 U980 ( .A1(n1261), .A2(n1099), .ZN(n1260) );
XNOR2_X1 U981 ( .A(n1262), .B(n1263), .ZN(n1099) );
XNOR2_X1 U982 ( .A(n1264), .B(n1265), .ZN(n1263) );
XNOR2_X1 U983 ( .A(G143), .B(n1266), .ZN(n1265) );
INV_X1 U984 ( .A(G134), .ZN(n1266) );
XOR2_X1 U985 ( .A(n1267), .B(n1268), .Z(n1262) );
AND2_X1 U986 ( .A1(n1269), .A2(G217), .ZN(n1268) );
XNOR2_X1 U987 ( .A(n1270), .B(n988), .ZN(n1267) );
INV_X1 U988 ( .A(G107), .ZN(n988) );
NAND2_X1 U989 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U990 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U991 ( .A1(KEYINPUT23), .A2(n1275), .ZN(n1274) );
NAND2_X1 U992 ( .A1(n1194), .A2(n1276), .ZN(n1275) );
INV_X1 U993 ( .A(n1277), .ZN(n1273) );
NAND2_X1 U994 ( .A1(G116), .A2(n1278), .ZN(n1271) );
NAND2_X1 U995 ( .A1(n1276), .A2(n1279), .ZN(n1278) );
NAND2_X1 U996 ( .A1(KEYINPUT23), .A2(n1277), .ZN(n1279) );
XOR2_X1 U997 ( .A(G122), .B(KEYINPUT26), .Z(n1277) );
INV_X1 U998 ( .A(KEYINPUT20), .ZN(n1276) );
XOR2_X1 U999 ( .A(KEYINPUT47), .B(n1208), .Z(n1261) );
NAND2_X1 U1000 ( .A1(n1175), .A2(n1185), .ZN(n1169) );
XNOR2_X1 U1001 ( .A(n1193), .B(KEYINPUT35), .ZN(n1185) );
INV_X1 U1002 ( .A(n1176), .ZN(n1193) );
XNOR2_X1 U1003 ( .A(n1035), .B(KEYINPUT53), .ZN(n1176) );
XNOR2_X1 U1004 ( .A(n1280), .B(n1117), .ZN(n1035) );
INV_X1 U1005 ( .A(G472), .ZN(n1117) );
NAND2_X1 U1006 ( .A1(n1281), .A2(n1208), .ZN(n1280) );
XNOR2_X1 U1007 ( .A(n1120), .B(n1282), .ZN(n1281) );
XOR2_X1 U1008 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U1009 ( .A1(KEYINPUT58), .A2(n1115), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(G113), .B(n1236), .ZN(n1115) );
XOR2_X1 U1011 ( .A(G119), .B(n1194), .Z(n1236) );
INV_X1 U1012 ( .A(G116), .ZN(n1194) );
NAND3_X1 U1013 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1283) );
NAND2_X1 U1014 ( .A1(KEYINPUT41), .A2(n1121), .ZN(n1287) );
NAND3_X1 U1015 ( .A1(n1288), .A2(n1289), .A3(n1243), .ZN(n1286) );
INV_X1 U1016 ( .A(KEYINPUT41), .ZN(n1289) );
OR2_X1 U1017 ( .A1(n1243), .A2(n1288), .ZN(n1285) );
NOR2_X1 U1018 ( .A1(KEYINPUT52), .A2(n1121), .ZN(n1288) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1256), .ZN(n1121) );
NOR2_X1 U1020 ( .A1(G953), .A2(G237), .ZN(n1256) );
INV_X1 U1021 ( .A(n1112), .ZN(n1243) );
XOR2_X1 U1022 ( .A(G101), .B(KEYINPUT15), .Z(n1112) );
XNOR2_X1 U1023 ( .A(n1219), .B(n1239), .ZN(n1120) );
XNOR2_X1 U1024 ( .A(n1290), .B(n1291), .ZN(n1239) );
XNOR2_X1 U1025 ( .A(G143), .B(n1264), .ZN(n1291) );
NAND2_X1 U1026 ( .A1(KEYINPUT37), .A2(n1213), .ZN(n1290) );
NAND3_X1 U1027 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1219) );
NAND2_X1 U1028 ( .A1(KEYINPUT43), .A2(n1295), .ZN(n1294) );
INV_X1 U1029 ( .A(n1073), .ZN(n1295) );
OR3_X1 U1030 ( .A1(n1296), .A2(KEYINPUT43), .A3(G131), .ZN(n1293) );
NAND2_X1 U1031 ( .A1(G131), .A2(n1296), .ZN(n1292) );
NAND2_X1 U1032 ( .A1(KEYINPUT45), .A2(n1073), .ZN(n1296) );
XOR2_X1 U1033 ( .A(n1297), .B(n1298), .Z(n1073) );
INV_X1 U1034 ( .A(n1299), .ZN(n1298) );
XNOR2_X1 U1035 ( .A(G134), .B(KEYINPUT10), .ZN(n1297) );
XNOR2_X1 U1036 ( .A(n1184), .B(KEYINPUT32), .ZN(n1175) );
NAND2_X1 U1037 ( .A1(n1300), .A2(n1301), .ZN(n1184) );
NAND2_X1 U1038 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
INV_X1 U1039 ( .A(KEYINPUT51), .ZN(n1303) );
NAND2_X1 U1040 ( .A1(n1045), .A2(n1304), .ZN(n1302) );
OR2_X1 U1041 ( .A1(n1048), .A2(n1047), .ZN(n1304) );
NAND2_X1 U1042 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U1043 ( .A1(KEYINPUT51), .A2(n1305), .ZN(n1300) );
XOR2_X1 U1044 ( .A(n1048), .B(n1047), .Z(n1305) );
AND2_X1 U1045 ( .A1(G217), .A2(n1220), .ZN(n1047) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1226), .ZN(n1220) );
NAND2_X1 U1047 ( .A1(n1094), .A2(n1208), .ZN(n1048) );
XNOR2_X1 U1048 ( .A(n1226), .B(KEYINPUT8), .ZN(n1208) );
INV_X1 U1049 ( .A(G902), .ZN(n1226) );
XNOR2_X1 U1050 ( .A(n1306), .B(n1307), .ZN(n1094) );
XOR2_X1 U1051 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1052 ( .A(n1310), .B(G110), .Z(n1309) );
NAND2_X1 U1053 ( .A1(KEYINPUT50), .A2(n1264), .ZN(n1310) );
INV_X1 U1054 ( .A(G128), .ZN(n1264) );
XNOR2_X1 U1055 ( .A(G119), .B(KEYINPUT17), .ZN(n1308) );
XOR2_X1 U1056 ( .A(n1257), .B(n1311), .Z(n1306) );
XNOR2_X1 U1057 ( .A(n1312), .B(n1299), .ZN(n1311) );
XOR2_X1 U1058 ( .A(G137), .B(KEYINPUT31), .Z(n1299) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1269), .ZN(n1312) );
AND2_X1 U1060 ( .A1(G234), .A2(n1060), .ZN(n1269) );
INV_X1 U1061 ( .A(G953), .ZN(n1060) );
XNOR2_X1 U1062 ( .A(n1127), .B(G125), .ZN(n1257) );
XOR2_X1 U1063 ( .A(G140), .B(n1213), .Z(n1127) );
XOR2_X1 U1064 ( .A(G146), .B(KEYINPUT54), .Z(n1213) );
endmodule


