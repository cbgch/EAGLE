//Key = 1100101100111010101000100111101101001011111011101010010100111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;

NAND2_X1 U724 ( .A1(n1002), .A2(n1003), .ZN(G9) );
NAND2_X1 U725 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U726 ( .A1(G107), .A2(n1006), .ZN(n1002) );
NAND2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
OR2_X1 U729 ( .A1(n1010), .A2(n1004), .ZN(n1007) );
NOR2_X1 U730 ( .A1(KEYINPUT19), .A2(n1011), .ZN(n1004) );
INV_X1 U731 ( .A(n1009), .ZN(n1011) );
INV_X1 U732 ( .A(KEYINPUT11), .ZN(n1010) );
NOR2_X1 U733 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U734 ( .A1(n1014), .A2(n1015), .A3(G953), .A4(n1016), .ZN(n1013) );
NOR4_X1 U735 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1015) );
NAND2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1018) );
NAND2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U738 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND3_X1 U739 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NAND3_X1 U741 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND2_X1 U742 ( .A1(KEYINPUT63), .A2(n1035), .ZN(n1034) );
NAND4_X1 U743 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND4_X1 U744 ( .A1(n1038), .A2(n1021), .A3(n1040), .A4(n1041), .ZN(n1033) );
NAND2_X1 U745 ( .A1(n1042), .A2(n1020), .ZN(n1041) );
OR2_X1 U746 ( .A1(n1043), .A2(KEYINPUT53), .ZN(n1042) );
NAND3_X1 U747 ( .A1(n1044), .A2(n1045), .A3(n1036), .ZN(n1040) );
NAND2_X1 U748 ( .A1(KEYINPUT53), .A2(n1046), .ZN(n1044) );
NAND3_X1 U749 ( .A1(n1039), .A2(n1047), .A3(n1036), .ZN(n1032) );
INV_X1 U750 ( .A(n1020), .ZN(n1036) );
NAND2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1021), .A2(n1050), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U755 ( .A1(n1038), .A2(n1055), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
OR2_X1 U757 ( .A1(n1058), .A2(KEYINPUT63), .ZN(n1057) );
NOR3_X1 U758 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n1012) );
AND4_X1 U759 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1016) );
NOR4_X1 U760 ( .A1(n1025), .A2(n1063), .A3(n1053), .A4(n1064), .ZN(n1062) );
INV_X1 U761 ( .A(n1065), .ZN(n1064) );
NOR3_X1 U762 ( .A1(n1017), .A2(n1066), .A3(n1067), .ZN(n1061) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XNOR2_X1 U764 ( .A(KEYINPUT15), .B(n1070), .ZN(n1068) );
NOR2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
XNOR2_X1 U766 ( .A(KEYINPUT14), .B(n1070), .ZN(n1072) );
XNOR2_X1 U767 ( .A(n1073), .B(n1074), .ZN(n1060) );
NOR2_X1 U768 ( .A1(G469), .A2(KEYINPUT21), .ZN(n1074) );
XNOR2_X1 U769 ( .A(KEYINPUT62), .B(n1075), .ZN(n1059) );
XOR2_X1 U770 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1082), .B(n1083), .Z(n1081) );
XNOR2_X1 U774 ( .A(n1084), .B(n1085), .ZN(n1083) );
NOR2_X1 U775 ( .A1(KEYINPUT8), .A2(n1086), .ZN(n1085) );
XNOR2_X1 U776 ( .A(n1087), .B(KEYINPUT0), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1088), .A2(KEYINPUT46), .ZN(n1084) );
XNOR2_X1 U778 ( .A(G125), .B(G140), .ZN(n1088) );
NOR2_X1 U779 ( .A1(G953), .A2(n1027), .ZN(n1078) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1076) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(G69) );
NAND2_X1 U783 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
OR2_X1 U784 ( .A1(n1090), .A2(G224), .ZN(n1094) );
NAND3_X1 U785 ( .A1(G953), .A2(n1095), .A3(n1096), .ZN(n1091) );
XNOR2_X1 U786 ( .A(n1093), .B(KEYINPUT23), .ZN(n1096) );
XNOR2_X1 U787 ( .A(n1097), .B(n1098), .ZN(n1093) );
NOR2_X1 U788 ( .A1(n1029), .A2(G953), .ZN(n1098) );
NAND2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U790 ( .A1(G953), .A2(n1101), .ZN(n1100) );
XNOR2_X1 U791 ( .A(n1102), .B(n1103), .ZN(n1099) );
XNOR2_X1 U792 ( .A(n1104), .B(KEYINPUT61), .ZN(n1103) );
NAND2_X1 U793 ( .A1(KEYINPUT60), .A2(n1105), .ZN(n1104) );
XOR2_X1 U794 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1095) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U797 ( .A(KEYINPUT37), .B(n1110), .Z(n1109) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(n1108) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1115), .ZN(G63) );
XNOR2_X1 U801 ( .A(n1116), .B(n1117), .ZN(n1115) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1114), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1110), .A2(n1119), .ZN(G60) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1114), .ZN(n1120) );
XNOR2_X1 U806 ( .A(G104), .B(n1123), .ZN(G6) );
NAND4_X1 U807 ( .A1(n1124), .A2(n1046), .A3(n1125), .A4(n1021), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U809 ( .A(n1051), .B(KEYINPUT6), .Z(n1124) );
NOR2_X1 U810 ( .A1(n1110), .A2(n1128), .ZN(G57) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U812 ( .A(KEYINPUT47), .B(n1131), .Z(n1130) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
AND2_X1 U814 ( .A1(n1133), .A2(n1132), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(n1132) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1114), .ZN(n1135) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U819 ( .A(KEYINPUT4), .B(n1141), .Z(n1137) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1139), .ZN(n1141) );
XNOR2_X1 U821 ( .A(n1142), .B(n1143), .ZN(n1139) );
NOR2_X1 U822 ( .A1(n1110), .A2(n1144), .ZN(G54) );
XOR2_X1 U823 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U824 ( .A(n1147), .B(n1143), .ZN(n1146) );
NOR2_X1 U825 ( .A1(n1148), .A2(n1114), .ZN(n1147) );
XNOR2_X1 U826 ( .A(n1149), .B(n1150), .ZN(n1145) );
NOR2_X1 U827 ( .A1(n1110), .A2(n1151), .ZN(G51) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U829 ( .A(n1154), .B(n1155), .ZN(n1153) );
XOR2_X1 U830 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U831 ( .A1(n1070), .A2(n1114), .ZN(n1157) );
NAND2_X1 U832 ( .A1(G902), .A2(n1158), .ZN(n1114) );
NAND2_X1 U833 ( .A1(n1029), .A2(n1027), .ZN(n1158) );
AND4_X1 U834 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1027) );
NOR4_X1 U835 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1046), .A2(n1038), .A3(n1167), .ZN(n1161) );
NAND3_X1 U837 ( .A1(n1168), .A2(n1169), .A3(n1030), .ZN(n1159) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
AND4_X1 U839 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1029) );
NOR4_X1 U840 ( .A1(n1176), .A2(n1177), .A3(n1009), .A4(n1178), .ZN(n1175) );
NOR3_X1 U841 ( .A1(n1043), .A2(n1179), .A3(n1180), .ZN(n1178) );
NOR3_X1 U842 ( .A1(n1045), .A2(n1179), .A3(n1180), .ZN(n1009) );
INV_X1 U843 ( .A(n1021), .ZN(n1179) );
NOR4_X1 U844 ( .A1(n1126), .A2(n1017), .A3(n1181), .A4(n1182), .ZN(n1177) );
XNOR2_X1 U845 ( .A(KEYINPUT39), .B(n1019), .ZN(n1182) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1184), .ZN(n1174) );
NAND2_X1 U847 ( .A1(KEYINPUT42), .A2(n1185), .ZN(n1156) );
NOR2_X1 U848 ( .A1(n1090), .A2(G952), .ZN(n1110) );
XNOR2_X1 U849 ( .A(n1160), .B(n1186), .ZN(G48) );
NOR2_X1 U850 ( .A1(KEYINPUT20), .A2(n1187), .ZN(n1186) );
INV_X1 U851 ( .A(G146), .ZN(n1187) );
NAND3_X1 U852 ( .A1(n1188), .A2(n1046), .A3(n1168), .ZN(n1160) );
XOR2_X1 U853 ( .A(G143), .B(n1166), .Z(G45) );
AND4_X1 U854 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1166) );
NOR2_X1 U855 ( .A1(n1058), .A2(n1193), .ZN(n1192) );
XNOR2_X1 U856 ( .A(n1194), .B(n1165), .ZN(G42) );
NOR4_X1 U857 ( .A1(n1195), .A2(n1193), .A3(n1043), .A4(n1056), .ZN(n1165) );
XOR2_X1 U858 ( .A(G137), .B(n1196), .Z(G39) );
NOR3_X1 U859 ( .A1(n1171), .A2(n1197), .A3(n1193), .ZN(n1196) );
XNOR2_X1 U860 ( .A(n1030), .B(KEYINPUT5), .ZN(n1197) );
NAND3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1039), .ZN(n1171) );
XOR2_X1 U862 ( .A(G134), .B(n1164), .Z(G36) );
NOR4_X1 U863 ( .A1(n1195), .A2(n1193), .A3(n1058), .A4(n1045), .ZN(n1164) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(G33) );
NAND2_X1 U865 ( .A1(G131), .A2(n1202), .ZN(n1201) );
XOR2_X1 U866 ( .A(n1203), .B(KEYINPUT56), .Z(n1200) );
OR2_X1 U867 ( .A1(n1202), .A2(G131), .ZN(n1203) );
NAND4_X1 U868 ( .A1(n1204), .A2(n1168), .A3(n1046), .A4(n1037), .ZN(n1202) );
XNOR2_X1 U869 ( .A(n1030), .B(KEYINPUT30), .ZN(n1204) );
INV_X1 U870 ( .A(n1195), .ZN(n1030) );
NAND2_X1 U871 ( .A1(n1026), .A2(n1205), .ZN(n1195) );
XNOR2_X1 U872 ( .A(n1206), .B(n1163), .ZN(G30) );
NOR3_X1 U873 ( .A1(n1181), .A2(n1045), .A3(n1193), .ZN(n1163) );
INV_X1 U874 ( .A(n1168), .ZN(n1193) );
NOR2_X1 U875 ( .A1(n1051), .A2(n1207), .ZN(n1168) );
INV_X1 U876 ( .A(n1208), .ZN(n1045) );
XOR2_X1 U877 ( .A(G101), .B(n1176), .Z(G3) );
NOR3_X1 U878 ( .A1(n1017), .A2(n1180), .A3(n1058), .ZN(n1176) );
INV_X1 U879 ( .A(n1037), .ZN(n1058) );
XOR2_X1 U880 ( .A(n1209), .B(n1210), .Z(G27) );
NOR2_X1 U881 ( .A1(KEYINPUT24), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U882 ( .A(KEYINPUT35), .B(n1212), .ZN(n1211) );
NAND3_X1 U883 ( .A1(n1167), .A2(n1046), .A3(n1213), .ZN(n1209) );
XNOR2_X1 U884 ( .A(n1038), .B(KEYINPUT45), .ZN(n1213) );
NOR3_X1 U885 ( .A1(n1023), .A2(n1207), .A3(n1056), .ZN(n1167) );
AND2_X1 U886 ( .A1(n1020), .A2(n1214), .ZN(n1207) );
NAND3_X1 U887 ( .A1(G902), .A2(n1215), .A3(n1080), .ZN(n1214) );
NOR2_X1 U888 ( .A1(n1090), .A2(G900), .ZN(n1080) );
XNOR2_X1 U889 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1216), .A2(n1021), .A3(n1189), .A4(n1190), .ZN(n1172) );
NOR2_X1 U891 ( .A1(n1199), .A2(n1198), .ZN(n1021) );
XNOR2_X1 U892 ( .A(G119), .B(n1217), .ZN(G21) );
NAND4_X1 U893 ( .A1(KEYINPUT33), .A2(n1188), .A3(n1218), .A4(n1038), .ZN(n1217) );
INV_X1 U894 ( .A(n1019), .ZN(n1038) );
NOR2_X1 U895 ( .A1(n1126), .A2(n1017), .ZN(n1218) );
INV_X1 U896 ( .A(n1181), .ZN(n1188) );
NAND3_X1 U897 ( .A1(n1198), .A2(n1199), .A3(n1191), .ZN(n1181) );
XNOR2_X1 U898 ( .A(G116), .B(n1219), .ZN(G18) );
NAND2_X1 U899 ( .A1(KEYINPUT27), .A2(n1220), .ZN(n1219) );
INV_X1 U900 ( .A(n1173), .ZN(n1220) );
NAND3_X1 U901 ( .A1(n1037), .A2(n1208), .A3(n1216), .ZN(n1173) );
NOR3_X1 U902 ( .A1(n1023), .A2(n1126), .A3(n1019), .ZN(n1216) );
INV_X1 U903 ( .A(n1191), .ZN(n1023) );
NOR2_X1 U904 ( .A1(n1190), .A2(n1221), .ZN(n1208) );
XOR2_X1 U905 ( .A(n1222), .B(n1184), .Z(G15) );
NOR4_X1 U906 ( .A1(n1127), .A2(n1126), .A3(n1019), .A4(n1170), .ZN(n1184) );
NAND2_X1 U907 ( .A1(n1037), .A2(n1046), .ZN(n1170) );
INV_X1 U908 ( .A(n1043), .ZN(n1046) );
NAND2_X1 U909 ( .A1(n1221), .A2(n1190), .ZN(n1043) );
INV_X1 U910 ( .A(n1189), .ZN(n1221) );
NOR2_X1 U911 ( .A1(n1199), .A2(n1075), .ZN(n1037) );
NAND2_X1 U912 ( .A1(n1054), .A2(n1223), .ZN(n1019) );
NAND2_X1 U913 ( .A1(KEYINPUT16), .A2(n1224), .ZN(n1222) );
XOR2_X1 U914 ( .A(G110), .B(n1183), .Z(G12) );
NOR3_X1 U915 ( .A1(n1017), .A2(n1180), .A3(n1056), .ZN(n1183) );
NAND2_X1 U916 ( .A1(n1075), .A2(n1199), .ZN(n1056) );
NAND3_X1 U917 ( .A1(n1225), .A2(n1226), .A3(n1065), .ZN(n1199) );
NAND2_X1 U918 ( .A1(n1227), .A2(n1113), .ZN(n1065) );
NAND2_X1 U919 ( .A1(n1063), .A2(n1228), .ZN(n1226) );
INV_X1 U920 ( .A(KEYINPUT43), .ZN(n1228) );
NOR2_X1 U921 ( .A1(n1113), .A2(n1227), .ZN(n1063) );
NOR2_X1 U922 ( .A1(n1229), .A2(n1112), .ZN(n1227) );
XNOR2_X1 U923 ( .A(n1230), .B(n1231), .ZN(n1112) );
XOR2_X1 U924 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U925 ( .A(G137), .B(G140), .ZN(n1233) );
NAND2_X1 U926 ( .A1(KEYINPUT55), .A2(n1234), .ZN(n1232) );
XOR2_X1 U927 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U928 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U929 ( .A1(KEYINPUT57), .A2(G119), .ZN(n1238) );
NOR2_X1 U930 ( .A1(KEYINPUT18), .A2(n1239), .ZN(n1237) );
XNOR2_X1 U931 ( .A(G128), .B(n1240), .ZN(n1235) );
XNOR2_X1 U932 ( .A(n1241), .B(n1242), .ZN(n1230) );
XOR2_X1 U933 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR2_X1 U934 ( .A1(G125), .A2(KEYINPUT3), .ZN(n1244) );
NOR2_X1 U935 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
INV_X1 U936 ( .A(G221), .ZN(n1245) );
XNOR2_X1 U937 ( .A(n1247), .B(KEYINPUT2), .ZN(n1229) );
NAND2_X1 U938 ( .A1(KEYINPUT43), .A2(n1113), .ZN(n1225) );
NAND2_X1 U939 ( .A1(G217), .A2(n1248), .ZN(n1113) );
INV_X1 U940 ( .A(n1198), .ZN(n1075) );
XOR2_X1 U941 ( .A(n1249), .B(n1136), .Z(n1198) );
INV_X1 U942 ( .A(G472), .ZN(n1136) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1247), .ZN(n1249) );
XOR2_X1 U944 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U945 ( .A(n1133), .B(n1143), .ZN(n1252) );
XNOR2_X1 U946 ( .A(n1253), .B(G101), .ZN(n1133) );
NAND3_X1 U947 ( .A1(n1254), .A2(n1255), .A3(G210), .ZN(n1253) );
XNOR2_X1 U948 ( .A(n1140), .B(n1256), .ZN(n1251) );
NOR2_X1 U949 ( .A1(KEYINPUT17), .A2(n1142), .ZN(n1256) );
XNOR2_X1 U950 ( .A(n1257), .B(n1258), .ZN(n1142) );
XOR2_X1 U951 ( .A(n1106), .B(n1259), .Z(n1140) );
XNOR2_X1 U952 ( .A(n1260), .B(KEYINPUT28), .ZN(n1259) );
NAND2_X1 U953 ( .A1(n1261), .A2(KEYINPUT48), .ZN(n1260) );
XNOR2_X1 U954 ( .A(n1107), .B(KEYINPUT29), .ZN(n1261) );
OR3_X1 U955 ( .A1(n1127), .A2(n1126), .A3(n1051), .ZN(n1180) );
OR2_X1 U956 ( .A1(n1054), .A2(n1053), .ZN(n1051) );
INV_X1 U957 ( .A(n1223), .ZN(n1053) );
NAND2_X1 U958 ( .A1(G221), .A2(n1248), .ZN(n1223) );
NAND2_X1 U959 ( .A1(n1262), .A2(n1247), .ZN(n1248) );
XOR2_X1 U960 ( .A(n1073), .B(n1263), .Z(n1054) );
NOR2_X1 U961 ( .A1(KEYINPUT9), .A2(n1148), .ZN(n1263) );
INV_X1 U962 ( .A(G469), .ZN(n1148) );
NAND2_X1 U963 ( .A1(n1264), .A2(n1247), .ZN(n1073) );
XNOR2_X1 U964 ( .A(n1150), .B(n1265), .ZN(n1264) );
XOR2_X1 U965 ( .A(n1266), .B(KEYINPUT26), .Z(n1265) );
NAND2_X1 U966 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U967 ( .A1(n1087), .A2(n1269), .ZN(n1268) );
NAND2_X1 U968 ( .A1(n1149), .A2(n1270), .ZN(n1269) );
NAND2_X1 U969 ( .A1(KEYINPUT52), .A2(n1271), .ZN(n1270) );
NAND3_X1 U970 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1267) );
INV_X1 U971 ( .A(KEYINPUT52), .ZN(n1274) );
NAND2_X1 U972 ( .A1(n1149), .A2(n1275), .ZN(n1273) );
NAND2_X1 U973 ( .A1(n1143), .A2(n1271), .ZN(n1275) );
INV_X1 U974 ( .A(n1087), .ZN(n1143) );
XOR2_X1 U975 ( .A(G131), .B(n1276), .Z(n1087) );
XOR2_X1 U976 ( .A(G137), .B(G134), .Z(n1276) );
NAND2_X1 U977 ( .A1(n1277), .A2(n1271), .ZN(n1272) );
INV_X1 U978 ( .A(KEYINPUT34), .ZN(n1271) );
INV_X1 U979 ( .A(n1149), .ZN(n1277) );
XNOR2_X1 U980 ( .A(n1278), .B(n1082), .ZN(n1149) );
XNOR2_X1 U981 ( .A(n1257), .B(G128), .ZN(n1082) );
XOR2_X1 U982 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U983 ( .A1(KEYINPUT59), .A2(n1281), .ZN(n1279) );
INV_X1 U984 ( .A(G104), .ZN(n1281) );
XNOR2_X1 U985 ( .A(n1282), .B(n1240), .ZN(n1150) );
XNOR2_X1 U986 ( .A(n1283), .B(n1194), .ZN(n1282) );
NAND2_X1 U987 ( .A1(G227), .A2(n1255), .ZN(n1283) );
AND2_X1 U988 ( .A1(n1020), .A2(n1284), .ZN(n1126) );
NAND4_X1 U989 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1101), .ZN(n1284) );
INV_X1 U990 ( .A(G898), .ZN(n1101) );
NAND3_X1 U991 ( .A1(n1215), .A2(n1090), .A3(G952), .ZN(n1020) );
INV_X1 U992 ( .A(G953), .ZN(n1090) );
NAND2_X1 U993 ( .A1(n1262), .A2(n1285), .ZN(n1215) );
XNOR2_X1 U994 ( .A(KEYINPUT32), .B(n1286), .ZN(n1285) );
XNOR2_X1 U995 ( .A(G234), .B(KEYINPUT38), .ZN(n1262) );
XOR2_X1 U996 ( .A(n1191), .B(KEYINPUT25), .Z(n1127) );
NOR2_X1 U997 ( .A1(n1026), .A2(n1025), .ZN(n1191) );
INV_X1 U998 ( .A(n1205), .ZN(n1025) );
NAND2_X1 U999 ( .A1(G214), .A2(n1287), .ZN(n1205) );
XOR2_X1 U1000 ( .A(n1071), .B(n1070), .Z(n1026) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1287), .ZN(n1070) );
NAND2_X1 U1002 ( .A1(n1247), .A2(n1286), .ZN(n1287) );
INV_X1 U1003 ( .A(n1069), .ZN(n1071) );
NAND2_X1 U1004 ( .A1(n1288), .A2(n1247), .ZN(n1069) );
XOR2_X1 U1005 ( .A(n1154), .B(n1289), .Z(n1288) );
XOR2_X1 U1006 ( .A(n1290), .B(n1185), .Z(n1289) );
AND2_X1 U1007 ( .A1(n1291), .A2(G224), .ZN(n1185) );
XNOR2_X1 U1008 ( .A(n1255), .B(KEYINPUT40), .ZN(n1291) );
NAND2_X1 U1009 ( .A1(KEYINPUT41), .A2(n1155), .ZN(n1290) );
XOR2_X1 U1010 ( .A(n1292), .B(n1258), .Z(n1155) );
XNOR2_X1 U1011 ( .A(n1293), .B(KEYINPUT13), .ZN(n1258) );
NAND2_X1 U1012 ( .A1(KEYINPUT31), .A2(n1206), .ZN(n1293) );
INV_X1 U1013 ( .A(G128), .ZN(n1206) );
XNOR2_X1 U1014 ( .A(n1294), .B(n1295), .ZN(n1154) );
INV_X1 U1015 ( .A(n1102), .ZN(n1295) );
XNOR2_X1 U1016 ( .A(n1296), .B(n1297), .ZN(n1102) );
XOR2_X1 U1017 ( .A(n1298), .B(n1280), .Z(n1297) );
XNOR2_X1 U1018 ( .A(G101), .B(n1005), .ZN(n1280) );
XOR2_X1 U1019 ( .A(n1299), .B(n1240), .Z(n1296) );
XOR2_X1 U1020 ( .A(G110), .B(KEYINPUT1), .Z(n1240) );
XNOR2_X1 U1021 ( .A(G104), .B(KEYINPUT10), .ZN(n1299) );
NAND2_X1 U1022 ( .A1(n1300), .A2(KEYINPUT12), .ZN(n1294) );
XNOR2_X1 U1023 ( .A(n1107), .B(n1106), .ZN(n1300) );
XNOR2_X1 U1024 ( .A(G113), .B(n1239), .ZN(n1106) );
INV_X1 U1025 ( .A(G119), .ZN(n1239) );
XOR2_X1 U1026 ( .A(G116), .B(KEYINPUT58), .Z(n1107) );
INV_X1 U1027 ( .A(n1039), .ZN(n1017) );
NOR2_X1 U1028 ( .A1(n1189), .A2(n1190), .ZN(n1039) );
XOR2_X1 U1029 ( .A(n1301), .B(n1122), .Z(n1190) );
INV_X1 U1030 ( .A(G475), .ZN(n1122) );
OR2_X1 U1031 ( .A1(n1121), .A2(G902), .ZN(n1301) );
XOR2_X1 U1032 ( .A(n1302), .B(n1224), .Z(n1121) );
INV_X1 U1033 ( .A(G113), .ZN(n1224) );
XOR2_X1 U1034 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1035 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1036 ( .A(n1194), .B(G131), .ZN(n1306) );
INV_X1 U1037 ( .A(G140), .ZN(n1194) );
XOR2_X1 U1038 ( .A(KEYINPUT36), .B(KEYINPUT22), .Z(n1305) );
XOR2_X1 U1039 ( .A(n1307), .B(n1308), .Z(n1303) );
XNOR2_X1 U1040 ( .A(G104), .B(n1309), .ZN(n1308) );
NAND3_X1 U1041 ( .A1(n1254), .A2(n1255), .A3(G214), .ZN(n1309) );
XNOR2_X1 U1042 ( .A(n1286), .B(KEYINPUT44), .ZN(n1254) );
INV_X1 U1043 ( .A(G237), .ZN(n1286) );
XOR2_X1 U1044 ( .A(n1292), .B(n1310), .Z(n1307) );
NOR2_X1 U1045 ( .A1(KEYINPUT49), .A2(n1298), .ZN(n1310) );
XNOR2_X1 U1046 ( .A(n1257), .B(n1212), .ZN(n1292) );
INV_X1 U1047 ( .A(G125), .ZN(n1212) );
XNOR2_X1 U1048 ( .A(G143), .B(n1241), .ZN(n1257) );
XOR2_X1 U1049 ( .A(G146), .B(KEYINPUT51), .Z(n1241) );
XOR2_X1 U1050 ( .A(n1311), .B(n1118), .Z(n1189) );
INV_X1 U1051 ( .A(G478), .ZN(n1118) );
NAND2_X1 U1052 ( .A1(n1116), .A2(n1247), .ZN(n1311) );
INV_X1 U1053 ( .A(G902), .ZN(n1247) );
XNOR2_X1 U1054 ( .A(n1312), .B(n1313), .ZN(n1116) );
XOR2_X1 U1055 ( .A(n1298), .B(n1314), .Z(n1313) );
XNOR2_X1 U1056 ( .A(n1005), .B(n1315), .ZN(n1314) );
NOR2_X1 U1057 ( .A1(n1246), .A2(n1316), .ZN(n1315) );
INV_X1 U1058 ( .A(G217), .ZN(n1316) );
NAND2_X1 U1059 ( .A1(n1317), .A2(n1255), .ZN(n1246) );
XOR2_X1 U1060 ( .A(G953), .B(KEYINPUT50), .Z(n1255) );
XNOR2_X1 U1061 ( .A(G234), .B(KEYINPUT7), .ZN(n1317) );
INV_X1 U1062 ( .A(G107), .ZN(n1005) );
XOR2_X1 U1063 ( .A(G122), .B(KEYINPUT54), .Z(n1298) );
XOR2_X1 U1064 ( .A(n1318), .B(n1319), .Z(n1312) );
XOR2_X1 U1065 ( .A(G143), .B(G134), .Z(n1319) );
XNOR2_X1 U1066 ( .A(G116), .B(G128), .ZN(n1318) );
endmodule


