//Key = 1001101100010100101100111101111011000000111111111010000100010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;

NAND2_X1 U739 ( .A1(n1014), .A2(n1015), .ZN(G9) );
NAND2_X1 U740 ( .A1(G107), .A2(n1016), .ZN(n1015) );
XOR2_X1 U741 ( .A(n1017), .B(KEYINPUT15), .Z(n1014) );
OR2_X1 U742 ( .A1(n1016), .A2(G107), .ZN(n1017) );
NOR2_X1 U743 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
NOR2_X1 U745 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XNOR2_X1 U746 ( .A(KEYINPUT62), .B(n1026), .ZN(n1025) );
NOR3_X1 U747 ( .A1(n1027), .A2(n1026), .A3(n1028), .ZN(n1022) );
NAND4_X1 U748 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1026) );
NOR2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND3_X1 U750 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1020) );
NAND3_X1 U751 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
INV_X1 U752 ( .A(n1034), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND3_X1 U754 ( .A1(n1031), .A2(n1043), .A3(n1044), .ZN(n1042) );
OR2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NAND3_X1 U756 ( .A1(n1030), .A2(n1047), .A3(n1029), .ZN(n1041) );
NAND3_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1044), .A2(n1051), .ZN(n1050) );
NAND2_X1 U759 ( .A1(n1031), .A2(n1052), .ZN(n1048) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U762 ( .A(n1057), .ZN(n1038) );
NOR3_X1 U763 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1018) );
INV_X1 U764 ( .A(n1035), .ZN(n1058) );
NAND4_X1 U765 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1035) );
NOR4_X1 U766 ( .A1(n1055), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1062) );
XOR2_X1 U767 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U768 ( .A1(G472), .A2(KEYINPUT2), .ZN(n1067) );
XNOR2_X1 U769 ( .A(n1068), .B(n1069), .ZN(n1064) );
NAND2_X1 U770 ( .A1(KEYINPUT48), .A2(n1070), .ZN(n1068) );
INV_X1 U771 ( .A(n1027), .ZN(n1063) );
NOR2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1061) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1072) );
NOR2_X1 U774 ( .A1(KEYINPUT61), .A2(n1075), .ZN(n1074) );
XOR2_X1 U775 ( .A(n1076), .B(n1077), .Z(n1060) );
XOR2_X1 U776 ( .A(n1078), .B(KEYINPUT10), .Z(n1076) );
XOR2_X1 U777 ( .A(n1056), .B(KEYINPUT35), .Z(n1059) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U779 ( .A1(n1081), .A2(n1036), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1036), .ZN(n1085) );
XOR2_X1 U783 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
INV_X1 U785 ( .A(n1091), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1092), .B(KEYINPUT33), .Z(n1089) );
NAND3_X1 U787 ( .A1(G900), .A2(n1088), .A3(G953), .ZN(n1084) );
XNOR2_X1 U788 ( .A(n1093), .B(n1094), .ZN(n1088) );
NOR2_X1 U789 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U790 ( .A(KEYINPUT54), .B(n1097), .Z(n1096) );
NOR2_X1 U791 ( .A1(G140), .A2(n1098), .ZN(n1097) );
XOR2_X1 U792 ( .A(n1099), .B(KEYINPUT51), .Z(n1098) );
NAND2_X1 U793 ( .A1(KEYINPUT45), .A2(n1100), .ZN(n1093) );
XOR2_X1 U794 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U795 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U796 ( .A1(KEYINPUT26), .A2(n1105), .ZN(n1104) );
XOR2_X1 U797 ( .A(n1106), .B(KEYINPUT21), .Z(n1101) );
XOR2_X1 U798 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U799 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1036), .ZN(n1110) );
NOR2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1109) );
NAND2_X1 U803 ( .A1(G953), .A2(n1113), .ZN(n1115) );
XOR2_X1 U804 ( .A(n1116), .B(n1117), .Z(n1114) );
NOR2_X1 U805 ( .A1(KEYINPUT39), .A2(n1118), .ZN(n1117) );
NAND2_X1 U806 ( .A1(n1036), .A2(n1119), .ZN(n1107) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(G66) );
NOR3_X1 U808 ( .A1(n1073), .A2(n1122), .A3(n1123), .ZN(n1121) );
AND3_X1 U809 ( .A1(n1124), .A2(G217), .A3(n1125), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1124), .ZN(n1122) );
AND2_X1 U811 ( .A1(n1021), .A2(G217), .ZN(n1126) );
INV_X1 U812 ( .A(n1127), .ZN(n1021) );
NOR2_X1 U813 ( .A1(n1120), .A2(n1128), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1077), .A2(n1129), .A3(n1130), .ZN(n1128) );
AND3_X1 U815 ( .A1(n1131), .A2(G478), .A3(n1125), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1131), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1127), .A2(n1078), .ZN(n1132) );
NOR3_X1 U818 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1136), .A2(G953), .A3(G952), .ZN(n1135) );
AND2_X1 U820 ( .A1(n1136), .A2(n1120), .ZN(n1134) );
INV_X1 U821 ( .A(KEYINPUT1), .ZN(n1136) );
XNOR2_X1 U822 ( .A(n1137), .B(n1138), .ZN(n1133) );
AND2_X1 U823 ( .A1(G475), .A2(n1125), .ZN(n1138) );
XNOR2_X1 U824 ( .A(G104), .B(n1139), .ZN(G6) );
NAND2_X1 U825 ( .A1(KEYINPUT16), .A2(n1140), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1120), .A2(n1141), .ZN(G57) );
XOR2_X1 U827 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U828 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U829 ( .A(n1146), .B(n1147), .Z(n1142) );
AND2_X1 U830 ( .A1(G472), .A2(n1125), .ZN(n1147) );
NAND2_X1 U831 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NOR2_X1 U832 ( .A1(n1120), .A2(n1150), .ZN(G54) );
XOR2_X1 U833 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U834 ( .A1(G469), .A2(n1125), .ZN(n1152) );
NOR3_X1 U835 ( .A1(n1153), .A2(KEYINPUT52), .A3(n1154), .ZN(n1151) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U837 ( .A(KEYINPUT8), .B(n1157), .Z(n1153) );
AND2_X1 U838 ( .A1(n1156), .A2(n1155), .ZN(n1157) );
NAND2_X1 U839 ( .A1(n1158), .A2(n1159), .ZN(n1155) );
NAND2_X1 U840 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U841 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1106), .ZN(n1163) );
INV_X1 U843 ( .A(n1165), .ZN(n1160) );
NAND2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(n1158) );
NAND2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1106), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1170), .B(n1171), .ZN(n1156) );
NAND2_X1 U848 ( .A1(KEYINPUT41), .A2(n1172), .ZN(n1170) );
NOR2_X1 U849 ( .A1(n1120), .A2(n1173), .ZN(G51) );
XNOR2_X1 U850 ( .A(n1174), .B(n1175), .ZN(n1173) );
XOR2_X1 U851 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND3_X1 U852 ( .A1(n1125), .A2(n1178), .A3(KEYINPUT24), .ZN(n1177) );
NOR2_X1 U853 ( .A1(n1179), .A2(n1127), .ZN(n1125) );
NOR3_X1 U854 ( .A1(n1119), .A2(n1091), .A3(n1092), .ZN(n1127) );
NAND4_X1 U855 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1092) );
NAND3_X1 U856 ( .A1(n1184), .A2(n1185), .A3(n1045), .ZN(n1180) );
NAND4_X1 U857 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1091) );
NAND4_X1 U858 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1187) );
XNOR2_X1 U859 ( .A(n1045), .B(KEYINPUT19), .ZN(n1190) );
NAND3_X1 U860 ( .A1(n1194), .A2(n1051), .A3(n1195), .ZN(n1186) );
NAND4_X1 U861 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1119) );
NOR4_X1 U862 ( .A1(n1200), .A2(n1201), .A3(n1140), .A4(n1202), .ZN(n1199) );
INV_X1 U863 ( .A(n1016), .ZN(n1202) );
NAND3_X1 U864 ( .A1(n1051), .A2(n1203), .A3(n1204), .ZN(n1016) );
AND3_X1 U865 ( .A1(n1204), .A2(n1203), .A3(n1184), .ZN(n1140) );
NOR2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(n1198) );
NOR3_X1 U867 ( .A1(n1207), .A2(n1208), .A3(n1024), .ZN(n1206) );
XOR2_X1 U868 ( .A(n1209), .B(KEYINPUT59), .Z(n1208) );
NAND3_X1 U869 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1176) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
INV_X1 U871 ( .A(KEYINPUT11), .ZN(n1214) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1099), .ZN(n1213) );
XOR2_X1 U873 ( .A(KEYINPUT38), .B(n1216), .Z(n1215) );
NAND2_X1 U874 ( .A1(KEYINPUT11), .A2(n1217), .ZN(n1210) );
NAND2_X1 U875 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
OR3_X1 U876 ( .A1(n1220), .A2(G125), .A3(KEYINPUT38), .ZN(n1219) );
NAND2_X1 U877 ( .A1(KEYINPUT38), .A2(n1220), .ZN(n1218) );
NOR2_X1 U878 ( .A1(n1036), .A2(G952), .ZN(n1120) );
XOR2_X1 U879 ( .A(n1221), .B(n1181), .Z(G48) );
NAND3_X1 U880 ( .A1(n1195), .A2(n1194), .A3(n1184), .ZN(n1181) );
XNOR2_X1 U881 ( .A(G143), .B(n1182), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1195), .A2(n1046), .A3(n1222), .A4(n1071), .ZN(n1182) );
NAND2_X1 U883 ( .A1(n1223), .A2(n1224), .ZN(G42) );
NAND2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U885 ( .A(KEYINPUT30), .B(n1227), .Z(n1223) );
NOR2_X1 U886 ( .A1(n1225), .A2(n1226), .ZN(n1227) );
NAND3_X1 U887 ( .A1(n1228), .A2(n1045), .A3(n1229), .ZN(n1226) );
NOR3_X1 U888 ( .A1(n1230), .A2(n1231), .A3(n1053), .ZN(n1229) );
XOR2_X1 U889 ( .A(n1057), .B(KEYINPUT3), .Z(n1228) );
XNOR2_X1 U890 ( .A(KEYINPUT0), .B(G140), .ZN(n1225) );
XNOR2_X1 U891 ( .A(G137), .B(n1183), .ZN(G39) );
NAND3_X1 U892 ( .A1(n1194), .A2(n1185), .A3(n1031), .ZN(n1183) );
XNOR2_X1 U893 ( .A(G134), .B(n1188), .ZN(G36) );
NAND3_X1 U894 ( .A1(n1185), .A2(n1051), .A3(n1046), .ZN(n1188) );
XNOR2_X1 U895 ( .A(G131), .B(n1189), .ZN(G33) );
NAND3_X1 U896 ( .A1(n1046), .A2(n1185), .A3(n1184), .ZN(n1189) );
NOR3_X1 U897 ( .A1(n1053), .A2(n1231), .A3(n1057), .ZN(n1185) );
NAND2_X1 U898 ( .A1(n1232), .A2(n1027), .ZN(n1057) );
XOR2_X1 U899 ( .A(n1233), .B(n1234), .Z(G30) );
NAND4_X1 U900 ( .A1(KEYINPUT6), .A2(n1195), .A3(n1051), .A4(n1235), .ZN(n1234) );
XOR2_X1 U901 ( .A(KEYINPUT5), .B(n1194), .Z(n1235) );
NOR3_X1 U902 ( .A1(n1024), .A2(n1231), .A3(n1053), .ZN(n1195) );
INV_X1 U903 ( .A(n1193), .ZN(n1231) );
XNOR2_X1 U904 ( .A(n1205), .B(n1236), .ZN(G3) );
NAND2_X1 U905 ( .A1(KEYINPUT7), .A2(G101), .ZN(n1236) );
AND4_X1 U906 ( .A1(n1046), .A2(n1031), .A3(n1204), .A4(n1237), .ZN(n1205) );
XOR2_X1 U907 ( .A(n1099), .B(n1238), .Z(G27) );
NAND4_X1 U908 ( .A1(n1191), .A2(n1045), .A3(n1192), .A4(n1193), .ZN(n1238) );
NAND2_X1 U909 ( .A1(n1034), .A2(n1239), .ZN(n1193) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1240), .A4(n1083), .ZN(n1239) );
INV_X1 U911 ( .A(G900), .ZN(n1083) );
XOR2_X1 U912 ( .A(n1241), .B(n1196), .Z(G24) );
NAND4_X1 U913 ( .A1(n1044), .A2(n1203), .A3(n1222), .A4(n1071), .ZN(n1196) );
NOR3_X1 U914 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1203) );
XOR2_X1 U915 ( .A(n1245), .B(n1197), .Z(G21) );
NAND4_X1 U916 ( .A1(n1044), .A2(n1031), .A3(n1194), .A4(n1237), .ZN(n1197) );
NOR2_X1 U917 ( .A1(n1030), .A2(n1029), .ZN(n1194) );
XNOR2_X1 U918 ( .A(G116), .B(n1246), .ZN(G18) );
NOR2_X1 U919 ( .A1(KEYINPUT60), .A2(n1247), .ZN(n1246) );
NOR2_X1 U920 ( .A1(n1244), .A2(n1207), .ZN(n1247) );
NAND3_X1 U921 ( .A1(n1046), .A2(n1051), .A3(n1044), .ZN(n1207) );
NOR2_X1 U922 ( .A1(n1071), .A2(n1248), .ZN(n1051) );
NAND2_X1 U923 ( .A1(n1249), .A2(n1250), .ZN(G15) );
NAND2_X1 U924 ( .A1(n1201), .A2(n1251), .ZN(n1250) );
XOR2_X1 U925 ( .A(KEYINPUT28), .B(n1252), .Z(n1249) );
NOR2_X1 U926 ( .A1(n1201), .A2(n1251), .ZN(n1252) );
AND3_X1 U927 ( .A1(n1046), .A2(n1237), .A3(n1191), .ZN(n1201) );
INV_X1 U928 ( .A(n1049), .ZN(n1191) );
NAND2_X1 U929 ( .A1(n1044), .A2(n1184), .ZN(n1049) );
INV_X1 U930 ( .A(n1230), .ZN(n1184) );
NAND2_X1 U931 ( .A1(n1248), .A2(n1071), .ZN(n1230) );
INV_X1 U932 ( .A(n1033), .ZN(n1044) );
NAND2_X1 U933 ( .A1(n1056), .A2(n1253), .ZN(n1033) );
XOR2_X1 U934 ( .A(KEYINPUT27), .B(n1055), .Z(n1253) );
INV_X1 U935 ( .A(n1254), .ZN(n1055) );
NOR2_X1 U936 ( .A1(n1243), .A2(n1029), .ZN(n1046) );
INV_X1 U937 ( .A(n1030), .ZN(n1243) );
XOR2_X1 U938 ( .A(n1200), .B(n1255), .Z(G12) );
NOR2_X1 U939 ( .A1(KEYINPUT20), .A2(n1256), .ZN(n1255) );
AND4_X1 U940 ( .A1(n1045), .A2(n1031), .A3(n1204), .A4(n1237), .ZN(n1200) );
INV_X1 U941 ( .A(n1244), .ZN(n1237) );
NAND2_X1 U942 ( .A1(n1192), .A2(n1209), .ZN(n1244) );
NAND2_X1 U943 ( .A1(n1257), .A2(n1034), .ZN(n1209) );
NAND3_X1 U944 ( .A1(n1240), .A2(n1036), .A3(G952), .ZN(n1034) );
XOR2_X1 U945 ( .A(KEYINPUT13), .B(n1258), .Z(n1257) );
AND4_X1 U946 ( .A1(n1113), .A2(n1240), .A3(G902), .A4(G953), .ZN(n1258) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1240) );
INV_X1 U948 ( .A(G898), .ZN(n1113) );
INV_X1 U949 ( .A(n1024), .ZN(n1192) );
NAND2_X1 U950 ( .A1(n1028), .A2(n1027), .ZN(n1024) );
NAND2_X1 U951 ( .A1(G214), .A2(n1259), .ZN(n1027) );
INV_X1 U952 ( .A(n1232), .ZN(n1028) );
XOR2_X1 U953 ( .A(n1260), .B(n1178), .Z(n1232) );
INV_X1 U954 ( .A(n1070), .ZN(n1178) );
NAND2_X1 U955 ( .A1(G210), .A2(n1259), .ZN(n1070) );
NAND2_X1 U956 ( .A1(n1261), .A2(n1179), .ZN(n1259) );
INV_X1 U957 ( .A(G237), .ZN(n1261) );
XOR2_X1 U958 ( .A(n1069), .B(KEYINPUT56), .Z(n1260) );
NAND4_X1 U959 ( .A1(n1262), .A2(n1179), .A3(n1263), .A4(n1264), .ZN(n1069) );
NAND3_X1 U960 ( .A1(n1174), .A2(n1216), .A3(G125), .ZN(n1264) );
NAND2_X1 U961 ( .A1(n1265), .A2(n1099), .ZN(n1263) );
XOR2_X1 U962 ( .A(n1174), .B(n1216), .Z(n1265) );
OR2_X1 U963 ( .A1(n1212), .A2(n1174), .ZN(n1262) );
XNOR2_X1 U964 ( .A(n1266), .B(n1267), .ZN(n1174) );
INV_X1 U965 ( .A(n1116), .ZN(n1267) );
XOR2_X1 U966 ( .A(n1268), .B(n1269), .Z(n1116) );
XOR2_X1 U967 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND2_X1 U968 ( .A1(KEYINPUT55), .A2(n1272), .ZN(n1271) );
XOR2_X1 U969 ( .A(KEYINPUT32), .B(n1273), .Z(n1272) );
XOR2_X1 U970 ( .A(n1256), .B(G122), .Z(n1268) );
INV_X1 U971 ( .A(G110), .ZN(n1256) );
XNOR2_X1 U972 ( .A(n1118), .B(n1274), .ZN(n1266) );
NOR2_X1 U973 ( .A1(G953), .A2(n1112), .ZN(n1274) );
INV_X1 U974 ( .A(G224), .ZN(n1112) );
XNOR2_X1 U975 ( .A(n1275), .B(G119), .ZN(n1118) );
NAND2_X1 U976 ( .A1(G125), .A2(n1220), .ZN(n1212) );
INV_X1 U977 ( .A(n1053), .ZN(n1204) );
NAND2_X1 U978 ( .A1(n1276), .A2(n1254), .ZN(n1053) );
NAND2_X1 U979 ( .A1(G221), .A2(n1277), .ZN(n1254) );
INV_X1 U980 ( .A(n1056), .ZN(n1276) );
XNOR2_X1 U981 ( .A(G469), .B(n1278), .ZN(n1056) );
NOR2_X1 U982 ( .A1(G902), .A2(n1279), .ZN(n1278) );
XOR2_X1 U983 ( .A(n1280), .B(n1281), .Z(n1279) );
NOR2_X1 U984 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U985 ( .A(n1284), .B(KEYINPUT46), .Z(n1283) );
NAND4_X1 U986 ( .A1(n1285), .A2(n1162), .A3(n1286), .A4(n1287), .ZN(n1284) );
OR2_X1 U987 ( .A1(n1167), .A2(KEYINPUT22), .ZN(n1287) );
NAND3_X1 U988 ( .A1(n1164), .A2(n1106), .A3(KEYINPUT22), .ZN(n1286) );
NAND2_X1 U989 ( .A1(n1288), .A2(n1169), .ZN(n1162) );
NOR3_X1 U990 ( .A1(n1285), .A2(n1289), .A3(n1290), .ZN(n1282) );
NOR2_X1 U991 ( .A1(n1291), .A2(n1167), .ZN(n1290) );
NAND2_X1 U992 ( .A1(n1288), .A2(n1164), .ZN(n1167) );
NOR2_X1 U993 ( .A1(n1288), .A2(n1292), .ZN(n1289) );
NOR2_X1 U994 ( .A1(n1169), .A2(n1291), .ZN(n1292) );
INV_X1 U995 ( .A(KEYINPUT22), .ZN(n1291) );
INV_X1 U996 ( .A(n1164), .ZN(n1169) );
XOR2_X1 U997 ( .A(n1270), .B(n1273), .Z(n1164) );
XOR2_X1 U998 ( .A(G104), .B(G107), .Z(n1273) );
INV_X1 U999 ( .A(n1106), .ZN(n1288) );
NAND2_X1 U1000 ( .A1(n1293), .A2(n1294), .ZN(n1106) );
NAND2_X1 U1001 ( .A1(G128), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n1296), .Z(n1293) );
NOR2_X1 U1003 ( .A1(G128), .A2(n1295), .ZN(n1296) );
XOR2_X1 U1004 ( .A(n1165), .B(KEYINPUT58), .Z(n1285) );
NAND2_X1 U1005 ( .A1(n1297), .A2(KEYINPUT43), .ZN(n1280) );
XOR2_X1 U1006 ( .A(n1172), .B(n1298), .Z(n1297) );
XOR2_X1 U1007 ( .A(KEYINPUT57), .B(n1171), .Z(n1298) );
XOR2_X1 U1008 ( .A(G110), .B(n1299), .Z(n1171) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1082), .ZN(n1299) );
INV_X1 U1010 ( .A(G227), .ZN(n1082) );
XNOR2_X1 U1011 ( .A(G140), .B(KEYINPUT18), .ZN(n1172) );
NOR2_X1 U1012 ( .A1(n1071), .A2(n1222), .ZN(n1031) );
INV_X1 U1013 ( .A(n1248), .ZN(n1222) );
NAND2_X1 U1014 ( .A1(n1300), .A2(n1301), .ZN(n1248) );
NAND2_X1 U1015 ( .A1(n1302), .A2(n1078), .ZN(n1301) );
INV_X1 U1016 ( .A(G478), .ZN(n1078) );
XOR2_X1 U1017 ( .A(KEYINPUT44), .B(n1077), .Z(n1302) );
NAND2_X1 U1018 ( .A1(n1303), .A2(G478), .ZN(n1300) );
XOR2_X1 U1019 ( .A(KEYINPUT14), .B(n1077), .Z(n1303) );
NOR2_X1 U1020 ( .A1(n1131), .A2(G902), .ZN(n1077) );
XOR2_X1 U1021 ( .A(n1304), .B(n1305), .Z(n1131) );
NOR2_X1 U1022 ( .A1(KEYINPUT37), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1023 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1024 ( .A(G128), .B(n1309), .Z(n1308) );
XOR2_X1 U1025 ( .A(G143), .B(G134), .Z(n1309) );
XNOR2_X1 U1026 ( .A(G107), .B(n1310), .ZN(n1307) );
XOR2_X1 U1027 ( .A(G122), .B(G116), .Z(n1310) );
NAND2_X1 U1028 ( .A1(G217), .A2(n1311), .ZN(n1304) );
XNOR2_X1 U1029 ( .A(n1312), .B(G475), .ZN(n1071) );
NAND2_X1 U1030 ( .A1(n1137), .A2(n1179), .ZN(n1312) );
XNOR2_X1 U1031 ( .A(n1313), .B(n1314), .ZN(n1137) );
XOR2_X1 U1032 ( .A(n1295), .B(n1105), .Z(n1314) );
INV_X1 U1033 ( .A(n1315), .ZN(n1105) );
XOR2_X1 U1034 ( .A(n1316), .B(n1317), .Z(n1313) );
XOR2_X1 U1035 ( .A(n1318), .B(n1319), .Z(n1316) );
AND2_X1 U1036 ( .A1(n1320), .A2(G214), .ZN(n1319) );
NAND2_X1 U1037 ( .A1(n1321), .A2(n1322), .ZN(n1318) );
OR2_X1 U1038 ( .A1(n1323), .A2(G104), .ZN(n1322) );
XOR2_X1 U1039 ( .A(n1324), .B(KEYINPUT12), .Z(n1321) );
NAND2_X1 U1040 ( .A1(G104), .A2(n1323), .ZN(n1324) );
XOR2_X1 U1041 ( .A(n1251), .B(n1241), .Z(n1323) );
INV_X1 U1042 ( .A(G122), .ZN(n1241) );
NOR2_X1 U1043 ( .A1(n1242), .A2(n1030), .ZN(n1045) );
XOR2_X1 U1044 ( .A(n1073), .B(n1075), .Z(n1030) );
NAND2_X1 U1045 ( .A1(n1325), .A2(G217), .ZN(n1075) );
XOR2_X1 U1046 ( .A(n1277), .B(KEYINPUT36), .Z(n1325) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1179), .ZN(n1277) );
NOR2_X1 U1048 ( .A1(n1124), .A2(G902), .ZN(n1073) );
XNOR2_X1 U1049 ( .A(n1326), .B(n1327), .ZN(n1124) );
XOR2_X1 U1050 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1051 ( .A(n1330), .B(n1331), .ZN(n1329) );
NAND3_X1 U1052 ( .A1(n1311), .A2(G221), .A3(KEYINPUT40), .ZN(n1331) );
AND2_X1 U1053 ( .A1(G234), .A2(n1036), .ZN(n1311) );
INV_X1 U1054 ( .A(G953), .ZN(n1036) );
NAND2_X1 U1055 ( .A1(KEYINPUT4), .A2(n1221), .ZN(n1330) );
INV_X1 U1056 ( .A(G146), .ZN(n1221) );
XOR2_X1 U1057 ( .A(n1332), .B(n1333), .Z(n1326) );
XOR2_X1 U1058 ( .A(KEYINPUT53), .B(G110), .Z(n1333) );
XOR2_X1 U1059 ( .A(n1334), .B(n1317), .Z(n1332) );
NOR2_X1 U1060 ( .A1(n1095), .A2(n1335), .ZN(n1317) );
NOR2_X1 U1061 ( .A1(n1099), .A2(G140), .ZN(n1335) );
AND2_X1 U1062 ( .A1(G140), .A2(n1099), .ZN(n1095) );
INV_X1 U1063 ( .A(G125), .ZN(n1099) );
NAND3_X1 U1064 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1334) );
OR2_X1 U1065 ( .A1(n1233), .A2(KEYINPUT23), .ZN(n1338) );
NAND3_X1 U1066 ( .A1(KEYINPUT23), .A2(n1233), .A3(G119), .ZN(n1337) );
NAND2_X1 U1067 ( .A1(n1339), .A2(n1245), .ZN(n1336) );
INV_X1 U1068 ( .A(G119), .ZN(n1245) );
NAND2_X1 U1069 ( .A1(KEYINPUT23), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1070 ( .A(KEYINPUT50), .B(G128), .Z(n1340) );
INV_X1 U1071 ( .A(n1029), .ZN(n1242) );
XOR2_X1 U1072 ( .A(n1066), .B(G472), .Z(n1029) );
NAND2_X1 U1073 ( .A1(n1341), .A2(n1179), .ZN(n1066) );
INV_X1 U1074 ( .A(G902), .ZN(n1179) );
XOR2_X1 U1075 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1076 ( .A(n1344), .B(KEYINPUT29), .ZN(n1343) );
NAND2_X1 U1077 ( .A1(KEYINPUT42), .A2(n1144), .ZN(n1344) );
XOR2_X1 U1078 ( .A(n1165), .B(n1220), .Z(n1144) );
INV_X1 U1079 ( .A(n1216), .ZN(n1220) );
XOR2_X1 U1080 ( .A(n1345), .B(n1295), .Z(n1216) );
XOR2_X1 U1081 ( .A(G143), .B(G146), .Z(n1295) );
XOR2_X1 U1082 ( .A(n1233), .B(KEYINPUT63), .Z(n1345) );
INV_X1 U1083 ( .A(G128), .ZN(n1233) );
XOR2_X1 U1084 ( .A(n1315), .B(n1103), .Z(n1165) );
XOR2_X1 U1085 ( .A(G134), .B(n1346), .Z(n1103) );
INV_X1 U1086 ( .A(n1328), .ZN(n1346) );
XNOR2_X1 U1087 ( .A(G137), .B(KEYINPUT17), .ZN(n1328) );
XNOR2_X1 U1088 ( .A(G131), .B(KEYINPUT25), .ZN(n1315) );
XOR2_X1 U1089 ( .A(n1347), .B(n1145), .Z(n1342) );
XNOR2_X1 U1090 ( .A(n1275), .B(n1348), .ZN(n1145) );
NOR2_X1 U1091 ( .A1(G119), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1092 ( .A(KEYINPUT49), .B(KEYINPUT34), .Z(n1349) );
XOR2_X1 U1093 ( .A(n1251), .B(n1350), .Z(n1275) );
XOR2_X1 U1094 ( .A(KEYINPUT9), .B(G116), .Z(n1350) );
INV_X1 U1095 ( .A(G113), .ZN(n1251) );
NAND2_X1 U1096 ( .A1(n1351), .A2(n1149), .ZN(n1347) );
NAND2_X1 U1097 ( .A1(n1270), .A2(n1352), .ZN(n1149) );
NAND2_X1 U1098 ( .A1(G210), .A2(n1320), .ZN(n1352) );
INV_X1 U1099 ( .A(G101), .ZN(n1270) );
XOR2_X1 U1100 ( .A(n1148), .B(KEYINPUT31), .Z(n1351) );
NAND3_X1 U1101 ( .A1(n1320), .A2(G101), .A3(G210), .ZN(n1148) );
NOR2_X1 U1102 ( .A1(G953), .A2(G237), .ZN(n1320) );
endmodule


