//Key = 1110101000110111001010000101000100011111000011001111101111001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376;

XNOR2_X1 U752 ( .A(n1042), .B(n1043), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1050) );
INV_X1 U757 ( .A(n1056), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1052) );
NAND3_X1 U759 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1046) );
NAND2_X1 U760 ( .A1(n1057), .A2(n1062), .ZN(n1061) );
NAND2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U762 ( .A1(n1065), .A2(n1066), .A3(n1058), .ZN(n1064) );
NAND3_X1 U763 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U766 ( .A(KEYINPUT48), .B(n1074), .Z(n1072) );
NAND3_X1 U767 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1068) );
XNOR2_X1 U768 ( .A(KEYINPUT47), .B(n1055), .ZN(n1076) );
NAND3_X1 U769 ( .A1(n1056), .A2(n1051), .A3(n1078), .ZN(n1067) );
INV_X1 U770 ( .A(KEYINPUT34), .ZN(n1051) );
NAND3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1070), .ZN(n1063) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1065), .A2(n1082), .ZN(n1081) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1058), .A2(n1085), .ZN(n1080) );
NAND2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
INV_X1 U778 ( .A(n1090), .ZN(n1086) );
AND3_X1 U779 ( .A1(n1059), .A2(n1060), .A3(n1091), .ZN(n1044) );
NAND4_X1 U780 ( .A1(n1092), .A2(n1070), .A3(n1093), .A4(n1094), .ZN(n1059) );
NOR4_X1 U781 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
AND2_X1 U782 ( .A1(n1099), .A2(KEYINPUT3), .ZN(n1097) );
NOR3_X1 U783 ( .A1(n1053), .A2(n1100), .A3(n1101), .ZN(n1093) );
NOR2_X1 U784 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U785 ( .A1(KEYINPUT3), .A2(n1104), .ZN(n1103) );
XOR2_X1 U786 ( .A(KEYINPUT32), .B(n1099), .Z(n1104) );
NOR3_X1 U787 ( .A1(n1105), .A2(KEYINPUT3), .A3(n1099), .ZN(n1100) );
XOR2_X1 U788 ( .A(n1106), .B(n1107), .Z(G72) );
XOR2_X1 U789 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U790 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U791 ( .A1(G900), .A2(G227), .ZN(n1110) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
OR2_X1 U793 ( .A1(n1060), .A2(n1113), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(n1111) );
XNOR2_X1 U795 ( .A(G125), .B(G140), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1116), .A2(KEYINPUT39), .ZN(n1114) );
XOR2_X1 U797 ( .A(n1117), .B(n1118), .Z(n1116) );
AND2_X1 U798 ( .A1(n1049), .A2(n1060), .ZN(n1106) );
NAND3_X1 U799 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(G69) );
XOR2_X1 U800 ( .A(KEYINPUT25), .B(n1122), .Z(n1121) );
NOR3_X1 U801 ( .A1(n1060), .A2(n1123), .A3(n1124), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1060), .ZN(n1120) );
XOR2_X1 U803 ( .A(n1123), .B(n1047), .Z(n1125) );
NAND3_X1 U804 ( .A1(n1123), .A2(n1124), .A3(G953), .ZN(n1119) );
AND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1124) );
AND2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
XOR2_X1 U807 ( .A(KEYINPUT0), .B(n1128), .Z(n1126) );
NOR2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR3_X1 U809 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
AND2_X1 U810 ( .A1(n1131), .A2(n1134), .ZN(n1129) );
INV_X1 U811 ( .A(KEYINPUT59), .ZN(n1131) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(G66) );
NOR3_X1 U813 ( .A1(n1099), .A2(n1137), .A3(n1138), .ZN(n1136) );
NOR4_X1 U814 ( .A1(n1139), .A2(n1140), .A3(KEYINPUT33), .A4(n1141), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NOR3_X1 U816 ( .A1(n1141), .A2(KEYINPUT33), .A3(n1144), .ZN(n1142) );
NOR2_X1 U817 ( .A1(n1049), .A2(n1047), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1135), .A2(n1145), .ZN(G63) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U820 ( .A(n1148), .B(KEYINPUT63), .Z(n1147) );
NAND2_X1 U821 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U822 ( .A(n1151), .B(KEYINPUT9), .ZN(n1149) );
NOR2_X1 U823 ( .A1(n1150), .A2(n1152), .ZN(n1146) );
INV_X1 U824 ( .A(n1151), .ZN(n1152) );
AND2_X1 U825 ( .A1(n1153), .A2(G478), .ZN(n1150) );
NOR2_X1 U826 ( .A1(n1135), .A2(n1154), .ZN(G60) );
XNOR2_X1 U827 ( .A(n1155), .B(n1156), .ZN(n1154) );
NAND2_X1 U828 ( .A1(n1153), .A2(G475), .ZN(n1156) );
XOR2_X1 U829 ( .A(G104), .B(n1157), .Z(G6) );
NOR4_X1 U830 ( .A1(KEYINPUT16), .A2(n1158), .A3(n1055), .A4(n1083), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1135), .A2(n1159), .ZN(G57) );
XOR2_X1 U832 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U833 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U834 ( .A1(KEYINPUT4), .A2(n1164), .ZN(n1163) );
NAND2_X1 U835 ( .A1(n1153), .A2(G472), .ZN(n1162) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(n1160) );
NAND2_X1 U837 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U838 ( .A(n1169), .B(KEYINPUT21), .Z(n1167) );
NOR2_X1 U839 ( .A1(n1135), .A2(n1170), .ZN(G54) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U841 ( .A(n1173), .B(n1118), .Z(n1172) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U843 ( .A1(n1153), .A2(G469), .ZN(n1174) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1171) );
XNOR2_X1 U845 ( .A(n1178), .B(n1179), .ZN(n1177) );
XNOR2_X1 U846 ( .A(n1180), .B(n1181), .ZN(n1176) );
NAND2_X1 U847 ( .A1(KEYINPUT6), .A2(n1182), .ZN(n1181) );
NAND2_X1 U848 ( .A1(KEYINPUT35), .A2(n1183), .ZN(n1180) );
NOR2_X1 U849 ( .A1(n1135), .A2(n1184), .ZN(G51) );
XOR2_X1 U850 ( .A(n1185), .B(n1134), .Z(n1184) );
XOR2_X1 U851 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U853 ( .A(KEYINPUT17), .B(n1190), .Z(n1189) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
AND2_X1 U855 ( .A1(n1192), .A2(n1191), .ZN(n1188) );
XOR2_X1 U856 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U857 ( .A1(G125), .A2(KEYINPUT19), .ZN(n1194) );
NAND2_X1 U858 ( .A1(n1153), .A2(n1195), .ZN(n1186) );
INV_X1 U859 ( .A(n1140), .ZN(n1153) );
NAND2_X1 U860 ( .A1(G902), .A2(n1196), .ZN(n1140) );
OR2_X1 U861 ( .A1(n1047), .A2(n1049), .ZN(n1196) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1049) );
NOR4_X1 U863 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
INV_X1 U864 ( .A(n1205), .ZN(n1201) );
NOR2_X1 U865 ( .A1(n1206), .A2(n1207), .ZN(n1199) );
INV_X1 U866 ( .A(n1208), .ZN(n1207) );
NAND4_X1 U867 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1047) );
NOR4_X1 U868 ( .A1(n1213), .A2(n1214), .A3(n1043), .A4(n1215), .ZN(n1212) );
INV_X1 U869 ( .A(n1216), .ZN(n1215) );
NOR3_X1 U870 ( .A1(n1055), .A2(n1158), .A3(n1084), .ZN(n1043) );
NOR3_X1 U871 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1211) );
NOR2_X1 U872 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
INV_X1 U873 ( .A(KEYINPUT44), .ZN(n1220) );
NOR4_X1 U874 ( .A1(KEYINPUT44), .A2(n1222), .A3(n1223), .A4(n1055), .ZN(n1218) );
NOR3_X1 U875 ( .A1(n1224), .A2(n1158), .A3(n1083), .ZN(n1217) );
XNOR2_X1 U876 ( .A(KEYINPUT52), .B(n1055), .ZN(n1224) );
INV_X1 U877 ( .A(n1078), .ZN(n1055) );
NOR2_X1 U878 ( .A1(n1060), .A2(G952), .ZN(n1135) );
XNOR2_X1 U879 ( .A(n1204), .B(n1225), .ZN(G48) );
NAND2_X1 U880 ( .A1(KEYINPUT50), .A2(G146), .ZN(n1225) );
AND3_X1 U881 ( .A1(n1226), .A2(n1056), .A3(n1227), .ZN(n1204) );
XOR2_X1 U882 ( .A(n1203), .B(n1228), .Z(G45) );
NOR2_X1 U883 ( .A1(KEYINPUT58), .A2(n1229), .ZN(n1228) );
AND3_X1 U884 ( .A1(n1223), .A2(n1056), .A3(n1230), .ZN(n1203) );
XNOR2_X1 U885 ( .A(n1178), .B(n1202), .ZN(G42) );
AND4_X1 U886 ( .A1(n1231), .A2(n1074), .A3(n1226), .A4(n1070), .ZN(n1202) );
XNOR2_X1 U887 ( .A(G137), .B(n1205), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1058), .A2(n1070), .A3(n1227), .ZN(n1205) );
XNOR2_X1 U889 ( .A(G134), .B(n1197), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1070), .A2(n1232), .A3(n1230), .ZN(n1197) );
XNOR2_X1 U891 ( .A(G131), .B(n1198), .ZN(G33) );
NAND3_X1 U892 ( .A1(n1226), .A2(n1070), .A3(n1230), .ZN(n1198) );
AND2_X1 U893 ( .A1(n1231), .A2(n1233), .ZN(n1230) );
NOR2_X1 U894 ( .A1(n1234), .A2(n1077), .ZN(n1070) );
XNOR2_X1 U895 ( .A(G128), .B(n1208), .ZN(G30) );
NAND3_X1 U896 ( .A1(n1232), .A2(n1056), .A3(n1227), .ZN(n1208) );
AND3_X1 U897 ( .A1(n1235), .A2(n1098), .A3(n1231), .ZN(n1227) );
AND2_X1 U898 ( .A1(n1090), .A2(n1236), .ZN(n1231) );
XNOR2_X1 U899 ( .A(n1214), .B(n1237), .ZN(G3) );
XNOR2_X1 U900 ( .A(KEYINPUT31), .B(n1164), .ZN(n1237) );
AND3_X1 U901 ( .A1(n1233), .A2(n1238), .A3(n1058), .ZN(n1214) );
XOR2_X1 U902 ( .A(n1206), .B(n1239), .Z(G27) );
NOR2_X1 U903 ( .A1(KEYINPUT30), .A2(n1240), .ZN(n1239) );
AND4_X1 U904 ( .A1(n1056), .A2(n1236), .A3(n1065), .A4(n1241), .ZN(n1206) );
AND2_X1 U905 ( .A1(n1226), .A2(n1074), .ZN(n1241) );
NAND2_X1 U906 ( .A1(n1242), .A2(n1243), .ZN(n1236) );
XOR2_X1 U907 ( .A(KEYINPUT27), .B(n1244), .Z(n1242) );
NOR4_X1 U908 ( .A1(n1245), .A2(n1113), .A3(n1060), .A4(n1246), .ZN(n1244) );
XNOR2_X1 U909 ( .A(G900), .B(KEYINPUT62), .ZN(n1113) );
XNOR2_X1 U910 ( .A(G122), .B(n1221), .ZN(G24) );
NAND3_X1 U911 ( .A1(n1247), .A2(n1078), .A3(n1223), .ZN(n1221) );
NOR2_X1 U912 ( .A1(n1092), .A2(n1248), .ZN(n1223) );
NOR2_X1 U913 ( .A1(n1098), .A2(n1235), .ZN(n1078) );
XNOR2_X1 U914 ( .A(G119), .B(n1209), .ZN(G21) );
NAND4_X1 U915 ( .A1(n1058), .A2(n1247), .A3(n1235), .A4(n1098), .ZN(n1209) );
XNOR2_X1 U916 ( .A(G116), .B(n1210), .ZN(G18) );
NAND3_X1 U917 ( .A1(n1233), .A2(n1232), .A3(n1247), .ZN(n1210) );
INV_X1 U918 ( .A(n1222), .ZN(n1247) );
INV_X1 U919 ( .A(n1084), .ZN(n1232) );
NAND2_X1 U920 ( .A1(n1248), .A2(n1249), .ZN(n1084) );
INV_X1 U921 ( .A(n1073), .ZN(n1233) );
NAND2_X1 U922 ( .A1(n1250), .A2(n1251), .ZN(G15) );
OR2_X1 U923 ( .A1(n1252), .A2(G113), .ZN(n1251) );
NAND2_X1 U924 ( .A1(n1253), .A2(G113), .ZN(n1250) );
NAND2_X1 U925 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U926 ( .A1(KEYINPUT40), .A2(n1213), .ZN(n1255) );
NAND2_X1 U927 ( .A1(n1252), .A2(n1256), .ZN(n1254) );
INV_X1 U928 ( .A(KEYINPUT40), .ZN(n1256) );
NAND2_X1 U929 ( .A1(KEYINPUT38), .A2(n1213), .ZN(n1252) );
NOR3_X1 U930 ( .A1(n1222), .A2(n1073), .A3(n1083), .ZN(n1213) );
INV_X1 U931 ( .A(n1226), .ZN(n1083) );
NOR2_X1 U932 ( .A1(n1249), .A2(n1248), .ZN(n1226) );
NAND2_X1 U933 ( .A1(n1257), .A2(n1098), .ZN(n1073) );
NAND2_X1 U934 ( .A1(n1065), .A2(n1258), .ZN(n1222) );
INV_X1 U935 ( .A(n1053), .ZN(n1065) );
NAND2_X1 U936 ( .A1(n1089), .A2(n1259), .ZN(n1053) );
XNOR2_X1 U937 ( .A(G110), .B(n1216), .ZN(G12) );
NAND3_X1 U938 ( .A1(n1058), .A2(n1238), .A3(n1074), .ZN(n1216) );
NOR2_X1 U939 ( .A1(n1098), .A2(n1257), .ZN(n1074) );
INV_X1 U940 ( .A(n1235), .ZN(n1257) );
XOR2_X1 U941 ( .A(n1102), .B(n1099), .Z(n1235) );
NOR2_X1 U942 ( .A1(n1143), .A2(G902), .ZN(n1099) );
INV_X1 U943 ( .A(n1139), .ZN(n1143) );
XNOR2_X1 U944 ( .A(n1260), .B(n1261), .ZN(n1139) );
NOR2_X1 U945 ( .A1(KEYINPUT46), .A2(n1262), .ZN(n1261) );
XOR2_X1 U946 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U947 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U948 ( .A(n1267), .B(n1182), .ZN(n1265) );
NAND2_X1 U949 ( .A1(KEYINPUT55), .A2(n1240), .ZN(n1267) );
XNOR2_X1 U950 ( .A(G119), .B(n1268), .ZN(n1263) );
XNOR2_X1 U951 ( .A(KEYINPUT43), .B(n1269), .ZN(n1268) );
NAND2_X1 U952 ( .A1(n1270), .A2(n1271), .ZN(n1260) );
NAND2_X1 U953 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U954 ( .A(n1274), .B(KEYINPUT28), .Z(n1270) );
OR2_X1 U955 ( .A1(n1272), .A2(n1273), .ZN(n1274) );
INV_X1 U956 ( .A(G137), .ZN(n1273) );
NAND3_X1 U957 ( .A1(G234), .A2(n1060), .A3(G221), .ZN(n1272) );
INV_X1 U958 ( .A(n1105), .ZN(n1102) );
NAND2_X1 U959 ( .A1(G217), .A2(n1275), .ZN(n1105) );
XNOR2_X1 U960 ( .A(n1276), .B(G472), .ZN(n1098) );
NAND2_X1 U961 ( .A1(n1277), .A2(n1246), .ZN(n1276) );
XOR2_X1 U962 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U963 ( .A(n1165), .B(n1280), .ZN(n1279) );
NOR2_X1 U964 ( .A1(G101), .A2(KEYINPUT53), .ZN(n1280) );
NAND2_X1 U965 ( .A1(G210), .A2(n1281), .ZN(n1165) );
NAND2_X1 U966 ( .A1(n1169), .A2(n1168), .ZN(n1278) );
NAND2_X1 U967 ( .A1(n1282), .A2(n1283), .ZN(n1168) );
NAND2_X1 U968 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U969 ( .A(n1193), .B(n1118), .ZN(n1282) );
NAND3_X1 U970 ( .A1(n1286), .A2(n1285), .A3(n1284), .ZN(n1169) );
XOR2_X1 U971 ( .A(n1287), .B(KEYINPUT7), .Z(n1284) );
OR2_X1 U972 ( .A1(n1288), .A2(G113), .ZN(n1287) );
NAND2_X1 U973 ( .A1(G113), .A2(n1288), .ZN(n1285) );
XNOR2_X1 U974 ( .A(n1289), .B(n1118), .ZN(n1286) );
INV_X1 U975 ( .A(n1158), .ZN(n1238) );
NAND2_X1 U976 ( .A1(n1090), .A2(n1258), .ZN(n1158) );
AND2_X1 U977 ( .A1(n1056), .A2(n1290), .ZN(n1258) );
NAND2_X1 U978 ( .A1(n1291), .A2(n1243), .ZN(n1290) );
INV_X1 U979 ( .A(n1057), .ZN(n1243) );
NOR3_X1 U980 ( .A1(n1245), .A2(G953), .A3(n1091), .ZN(n1057) );
INV_X1 U981 ( .A(G952), .ZN(n1091) );
OR3_X1 U982 ( .A1(n1127), .A2(n1245), .A3(n1246), .ZN(n1291) );
NOR2_X1 U983 ( .A1(n1292), .A2(n1293), .ZN(n1245) );
NAND2_X1 U984 ( .A1(G953), .A2(n1294), .ZN(n1127) );
XOR2_X1 U985 ( .A(KEYINPUT37), .B(G898), .Z(n1294) );
NOR2_X1 U986 ( .A1(n1075), .A2(n1077), .ZN(n1056) );
AND2_X1 U987 ( .A1(G214), .A2(n1295), .ZN(n1077) );
INV_X1 U988 ( .A(n1234), .ZN(n1075) );
XNOR2_X1 U989 ( .A(n1296), .B(n1195), .ZN(n1234) );
AND2_X1 U990 ( .A1(G210), .A2(n1295), .ZN(n1195) );
NAND2_X1 U991 ( .A1(n1246), .A2(n1292), .ZN(n1295) );
INV_X1 U992 ( .A(G237), .ZN(n1292) );
NAND2_X1 U993 ( .A1(n1297), .A2(n1246), .ZN(n1296) );
XNOR2_X1 U994 ( .A(n1134), .B(n1298), .ZN(n1297) );
XOR2_X1 U995 ( .A(n1299), .B(KEYINPUT10), .Z(n1298) );
NAND3_X1 U996 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1299) );
OR2_X1 U997 ( .A1(n1191), .A2(KEYINPUT57), .ZN(n1302) );
NAND3_X1 U998 ( .A1(KEYINPUT57), .A2(n1303), .A3(n1304), .ZN(n1301) );
OR2_X1 U999 ( .A1(n1304), .A2(n1303), .ZN(n1300) );
AND2_X1 U1000 ( .A1(KEYINPUT18), .A2(n1191), .ZN(n1303) );
AND2_X1 U1001 ( .A1(G224), .A2(n1060), .ZN(n1191) );
XNOR2_X1 U1002 ( .A(G125), .B(n1289), .ZN(n1304) );
INV_X1 U1003 ( .A(n1193), .ZN(n1289) );
XOR2_X1 U1004 ( .A(G146), .B(n1305), .Z(n1193) );
XOR2_X1 U1005 ( .A(n1132), .B(n1133), .Z(n1134) );
XOR2_X1 U1006 ( .A(n1306), .B(n1307), .Z(n1133) );
XNOR2_X1 U1007 ( .A(G107), .B(n1308), .ZN(n1307) );
NAND2_X1 U1008 ( .A1(KEYINPUT56), .A2(n1164), .ZN(n1308) );
XOR2_X1 U1009 ( .A(n1309), .B(n1310), .Z(n1306) );
NAND2_X1 U1010 ( .A1(KEYINPUT45), .A2(n1288), .ZN(n1309) );
XNOR2_X1 U1011 ( .A(n1311), .B(G119), .ZN(n1288) );
XOR2_X1 U1012 ( .A(n1312), .B(KEYINPUT54), .Z(n1132) );
NAND3_X1 U1013 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
NAND2_X1 U1014 ( .A1(G110), .A2(n1316), .ZN(n1315) );
INV_X1 U1015 ( .A(G122), .ZN(n1316) );
NAND2_X1 U1016 ( .A1(KEYINPUT42), .A2(n1317), .ZN(n1314) );
NAND2_X1 U1017 ( .A1(n1318), .A2(n1182), .ZN(n1317) );
XNOR2_X1 U1018 ( .A(KEYINPUT15), .B(G122), .ZN(n1318) );
NAND2_X1 U1019 ( .A1(n1319), .A2(n1320), .ZN(n1313) );
INV_X1 U1020 ( .A(KEYINPUT42), .ZN(n1320) );
NAND2_X1 U1021 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
OR2_X1 U1022 ( .A1(G122), .A2(KEYINPUT15), .ZN(n1322) );
NAND3_X1 U1023 ( .A1(G122), .A2(n1182), .A3(KEYINPUT15), .ZN(n1321) );
NOR2_X1 U1024 ( .A1(n1089), .A2(n1088), .ZN(n1090) );
INV_X1 U1025 ( .A(n1259), .ZN(n1088) );
NAND2_X1 U1026 ( .A1(G221), .A2(n1275), .ZN(n1259) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1246), .ZN(n1275) );
XOR2_X1 U1028 ( .A(n1323), .B(G469), .Z(n1089) );
NAND2_X1 U1029 ( .A1(n1324), .A2(n1246), .ZN(n1323) );
XOR2_X1 U1030 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1031 ( .A(n1327), .B(n1175), .ZN(n1326) );
XNOR2_X1 U1032 ( .A(n1117), .B(KEYINPUT36), .ZN(n1175) );
NAND2_X1 U1033 ( .A1(n1328), .A2(n1329), .ZN(n1117) );
NAND2_X1 U1034 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1035 ( .A(KEYINPUT23), .B(n1269), .ZN(n1331) );
XNOR2_X1 U1036 ( .A(G146), .B(n1229), .ZN(n1330) );
XOR2_X1 U1037 ( .A(n1332), .B(KEYINPUT22), .Z(n1328) );
NAND2_X1 U1038 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XNOR2_X1 U1039 ( .A(KEYINPUT23), .B(G128), .ZN(n1334) );
XNOR2_X1 U1040 ( .A(G143), .B(G146), .ZN(n1333) );
NAND2_X1 U1041 ( .A1(KEYINPUT13), .A2(n1118), .ZN(n1327) );
XNOR2_X1 U1042 ( .A(n1335), .B(n1336), .ZN(n1118) );
XNOR2_X1 U1043 ( .A(G137), .B(n1337), .ZN(n1336) );
XNOR2_X1 U1044 ( .A(KEYINPUT61), .B(KEYINPUT14), .ZN(n1337) );
XNOR2_X1 U1045 ( .A(G131), .B(G134), .ZN(n1335) );
XOR2_X1 U1046 ( .A(n1338), .B(n1339), .Z(n1325) );
XOR2_X1 U1047 ( .A(n1179), .B(n1340), .Z(n1339) );
NOR2_X1 U1048 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1049 ( .A(n1343), .B(KEYINPUT49), .Z(n1342) );
NAND2_X1 U1050 ( .A1(n1344), .A2(n1178), .ZN(n1343) );
XNOR2_X1 U1051 ( .A(KEYINPUT12), .B(n1182), .ZN(n1344) );
INV_X1 U1052 ( .A(G110), .ZN(n1182) );
NOR2_X1 U1053 ( .A1(G110), .A2(n1345), .ZN(n1341) );
XNOR2_X1 U1054 ( .A(KEYINPUT20), .B(n1178), .ZN(n1345) );
INV_X1 U1055 ( .A(G140), .ZN(n1178) );
AND2_X1 U1056 ( .A1(G227), .A2(n1060), .ZN(n1179) );
INV_X1 U1057 ( .A(G953), .ZN(n1060) );
NAND2_X1 U1058 ( .A1(KEYINPUT11), .A2(n1183), .ZN(n1338) );
XOR2_X1 U1059 ( .A(n1346), .B(n1347), .Z(n1183) );
NOR2_X1 U1060 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1061 ( .A(KEYINPUT41), .B(n1350), .Z(n1349) );
NOR2_X1 U1062 ( .A1(G104), .A2(n1042), .ZN(n1350) );
AND2_X1 U1063 ( .A1(n1042), .A2(G104), .ZN(n1348) );
INV_X1 U1064 ( .A(G107), .ZN(n1042) );
NAND2_X1 U1065 ( .A1(KEYINPUT51), .A2(n1164), .ZN(n1346) );
INV_X1 U1066 ( .A(G101), .ZN(n1164) );
AND2_X1 U1067 ( .A1(n1092), .A2(n1248), .ZN(n1058) );
NOR2_X1 U1068 ( .A1(n1351), .A2(n1096), .ZN(n1248) );
NOR3_X1 U1069 ( .A1(G475), .A2(G902), .A3(n1155), .ZN(n1096) );
INV_X1 U1070 ( .A(n1352), .ZN(n1155) );
XOR2_X1 U1071 ( .A(n1095), .B(KEYINPUT24), .Z(n1351) );
AND2_X1 U1072 ( .A1(G475), .A2(n1353), .ZN(n1095) );
NAND2_X1 U1073 ( .A1(n1246), .A2(n1352), .ZN(n1353) );
NAND3_X1 U1074 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1352) );
NAND2_X1 U1075 ( .A1(KEYINPUT29), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1076 ( .A1(n1358), .A2(n1359), .ZN(n1355) );
XOR2_X1 U1077 ( .A(KEYINPUT1), .B(n1360), .Z(n1359) );
XNOR2_X1 U1078 ( .A(n1240), .B(n1266), .ZN(n1358) );
INV_X1 U1079 ( .A(G125), .ZN(n1240) );
NAND2_X1 U1080 ( .A1(n1361), .A2(n1362), .ZN(n1354) );
XOR2_X1 U1081 ( .A(KEYINPUT5), .B(n1360), .Z(n1362) );
XNOR2_X1 U1082 ( .A(n1363), .B(n1364), .ZN(n1360) );
XNOR2_X1 U1083 ( .A(n1229), .B(G131), .ZN(n1364) );
INV_X1 U1084 ( .A(G143), .ZN(n1229) );
XOR2_X1 U1085 ( .A(n1365), .B(n1366), .Z(n1363) );
AND2_X1 U1086 ( .A1(n1281), .A2(G214), .ZN(n1366) );
NOR2_X1 U1087 ( .A1(G953), .A2(G237), .ZN(n1281) );
OR2_X1 U1088 ( .A1(n1357), .A2(KEYINPUT29), .ZN(n1365) );
XOR2_X1 U1089 ( .A(n1367), .B(n1310), .Z(n1357) );
XOR2_X1 U1090 ( .A(G104), .B(G113), .Z(n1310) );
XNOR2_X1 U1091 ( .A(G122), .B(KEYINPUT26), .ZN(n1367) );
XNOR2_X1 U1092 ( .A(G125), .B(n1266), .ZN(n1361) );
XOR2_X1 U1093 ( .A(G146), .B(G140), .Z(n1266) );
INV_X1 U1094 ( .A(n1249), .ZN(n1092) );
XNOR2_X1 U1095 ( .A(n1368), .B(G478), .ZN(n1249) );
NAND2_X1 U1096 ( .A1(n1151), .A2(n1246), .ZN(n1368) );
INV_X1 U1097 ( .A(G902), .ZN(n1246) );
XNOR2_X1 U1098 ( .A(n1369), .B(n1370), .ZN(n1151) );
XOR2_X1 U1099 ( .A(n1371), .B(n1372), .Z(n1370) );
XOR2_X1 U1100 ( .A(n1373), .B(n1374), .Z(n1372) );
NOR3_X1 U1101 ( .A1(n1293), .A2(G953), .A3(n1141), .ZN(n1374) );
INV_X1 U1102 ( .A(G217), .ZN(n1141) );
INV_X1 U1103 ( .A(G234), .ZN(n1293) );
NAND2_X1 U1104 ( .A1(KEYINPUT2), .A2(n1311), .ZN(n1373) );
INV_X1 U1105 ( .A(G116), .ZN(n1311) );
NAND2_X1 U1106 ( .A1(KEYINPUT60), .A2(n1305), .ZN(n1371) );
XNOR2_X1 U1107 ( .A(n1269), .B(G143), .ZN(n1305) );
INV_X1 U1108 ( .A(G128), .ZN(n1269) );
XOR2_X1 U1109 ( .A(n1375), .B(n1376), .Z(n1369) );
NOR2_X1 U1110 ( .A1(KEYINPUT8), .A2(G107), .ZN(n1376) );
XNOR2_X1 U1111 ( .A(G134), .B(G122), .ZN(n1375) );
endmodule


