//Key = 1010000011011011101100111111101001010011110100101110101101100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;

XNOR2_X1 U755 ( .A(G107), .B(n1058), .ZN(G9) );
NAND4_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(G75) );
NOR3_X1 U757 ( .A1(n1063), .A2(G953), .A3(n1064), .ZN(n1062) );
INV_X1 U758 ( .A(n1065), .ZN(n1064) );
NOR4_X1 U759 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1063) );
INV_X1 U760 ( .A(n1070), .ZN(n1069) );
XNOR2_X1 U761 ( .A(n1071), .B(n1072), .ZN(n1068) );
NAND2_X1 U762 ( .A1(KEYINPUT16), .A2(n1073), .ZN(n1071) );
NAND3_X1 U763 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1067) );
NAND3_X1 U764 ( .A1(G475), .A2(n1077), .A3(n1078), .ZN(n1075) );
INV_X1 U765 ( .A(KEYINPUT4), .ZN(n1078) );
NAND2_X1 U766 ( .A1(KEYINPUT4), .A2(n1079), .ZN(n1074) );
NAND4_X1 U767 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1066) );
XNOR2_X1 U768 ( .A(n1084), .B(n1085), .ZN(n1080) );
NAND2_X1 U769 ( .A1(KEYINPUT12), .A2(n1086), .ZN(n1085) );
NAND2_X1 U770 ( .A1(n1087), .A2(n1088), .ZN(n1060) );
NAND2_X1 U771 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U772 ( .A1(n1070), .A2(n1091), .A3(n1092), .ZN(n1090) );
NAND2_X1 U773 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND2_X1 U774 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U775 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND3_X1 U776 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NAND2_X1 U777 ( .A1(n1102), .A2(n1103), .ZN(n1093) );
INV_X1 U778 ( .A(n1104), .ZN(n1103) );
NAND3_X1 U779 ( .A1(n1095), .A2(n1105), .A3(n1102), .ZN(n1089) );
NAND3_X1 U780 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
OR2_X1 U781 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND3_X1 U782 ( .A1(n1111), .A2(n1112), .A3(n1070), .ZN(n1107) );
NAND2_X1 U783 ( .A1(n1100), .A2(n1081), .ZN(n1112) );
INV_X1 U784 ( .A(KEYINPUT45), .ZN(n1100) );
NAND2_X1 U785 ( .A1(n1113), .A2(n1114), .ZN(n1106) );
XNOR2_X1 U786 ( .A(n1070), .B(KEYINPUT61), .ZN(n1113) );
INV_X1 U787 ( .A(n1115), .ZN(n1087) );
XOR2_X1 U788 ( .A(n1116), .B(n1117), .Z(G72) );
NOR2_X1 U789 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1118) );
NAND2_X1 U791 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
NAND2_X1 U792 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U793 ( .A(KEYINPUT22), .B(n1124), .Z(n1120) );
NOR2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1124) );
NAND2_X1 U795 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND2_X1 U796 ( .A1(G953), .A2(n1127), .ZN(n1126) );
XOR2_X1 U797 ( .A(n1128), .B(n1129), .Z(n1125) );
XNOR2_X1 U798 ( .A(G131), .B(n1130), .ZN(n1129) );
NAND2_X1 U799 ( .A1(KEYINPUT58), .A2(n1131), .ZN(n1130) );
NAND2_X1 U800 ( .A1(n1132), .A2(n1133), .ZN(n1128) );
NAND2_X1 U801 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U802 ( .A(KEYINPUT26), .B(n1136), .Z(n1134) );
NAND2_X1 U803 ( .A1(G140), .A2(n1137), .ZN(n1132) );
XNOR2_X1 U804 ( .A(n1136), .B(KEYINPUT39), .ZN(n1137) );
XOR2_X1 U805 ( .A(G125), .B(n1138), .Z(n1136) );
NOR2_X1 U806 ( .A1(KEYINPUT51), .A2(n1139), .ZN(n1138) );
AND2_X1 U807 ( .A1(n1140), .A2(n1119), .ZN(n1122) );
NAND2_X1 U808 ( .A1(n1059), .A2(n1141), .ZN(n1140) );
XNOR2_X1 U809 ( .A(KEYINPUT19), .B(n1065), .ZN(n1141) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(G69) );
NAND2_X1 U811 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
OR2_X1 U812 ( .A1(n1119), .A2(G224), .ZN(n1144) );
NAND3_X1 U813 ( .A1(G953), .A2(n1146), .A3(n1147), .ZN(n1142) );
INV_X1 U814 ( .A(n1145), .ZN(n1147) );
NAND2_X1 U815 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
OR4_X1 U816 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(KEYINPUT44), .ZN(n1149) );
NOR2_X1 U817 ( .A1(n1119), .A2(G898), .ZN(n1152) );
NAND4_X1 U818 ( .A1(n1150), .A2(n1119), .A3(n1153), .A4(n1154), .ZN(n1148) );
NAND2_X1 U819 ( .A1(KEYINPUT1), .A2(n1151), .ZN(n1154) );
OR3_X1 U820 ( .A1(KEYINPUT1), .A2(KEYINPUT44), .A3(n1151), .ZN(n1153) );
XNOR2_X1 U821 ( .A(n1155), .B(KEYINPUT38), .ZN(n1151) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XNOR2_X1 U824 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1162), .ZN(G63) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U828 ( .A1(n1165), .A2(n1161), .ZN(n1163) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1166), .ZN(G60) );
NOR3_X1 U830 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
AND2_X1 U831 ( .A1(n1170), .A2(KEYINPUT20), .ZN(n1169) );
NOR3_X1 U832 ( .A1(KEYINPUT20), .A2(n1171), .A3(n1170), .ZN(n1168) );
NOR3_X1 U833 ( .A1(n1161), .A2(KEYINPUT7), .A3(n1079), .ZN(n1171) );
NOR3_X1 U834 ( .A1(n1161), .A2(n1172), .A3(n1079), .ZN(n1167) );
NOR2_X1 U835 ( .A1(n1173), .A2(KEYINPUT20), .ZN(n1172) );
NOR2_X1 U836 ( .A1(KEYINPUT7), .A2(n1174), .ZN(n1173) );
XOR2_X1 U837 ( .A(G104), .B(n1175), .Z(G6) );
NOR2_X1 U838 ( .A1(n1156), .A2(n1176), .ZN(G57) );
XOR2_X1 U839 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U840 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
OR2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U842 ( .A1(n1183), .A2(n1181), .ZN(n1179) );
XNOR2_X1 U843 ( .A(n1184), .B(n1185), .ZN(n1181) );
NOR2_X1 U844 ( .A1(KEYINPUT32), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U845 ( .A(n1187), .B(KEYINPUT34), .ZN(n1186) );
XOR2_X1 U846 ( .A(KEYINPUT47), .B(n1182), .Z(n1183) );
NOR2_X1 U847 ( .A1(n1161), .A2(n1188), .ZN(n1182) );
INV_X1 U848 ( .A(G472), .ZN(n1188) );
NAND2_X1 U849 ( .A1(KEYINPUT14), .A2(n1189), .ZN(n1177) );
NOR2_X1 U850 ( .A1(n1156), .A2(n1190), .ZN(G54) );
NOR2_X1 U851 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U852 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U853 ( .A1(n1086), .A2(n1161), .ZN(n1194) );
INV_X1 U854 ( .A(G469), .ZN(n1086) );
NOR2_X1 U855 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
XOR2_X1 U856 ( .A(n1197), .B(n1198), .Z(n1196) );
INV_X1 U857 ( .A(KEYINPUT0), .ZN(n1195) );
NOR2_X1 U858 ( .A1(KEYINPUT0), .A2(n1199), .ZN(n1191) );
XNOR2_X1 U859 ( .A(n1198), .B(n1197), .ZN(n1199) );
XNOR2_X1 U860 ( .A(n1200), .B(KEYINPUT29), .ZN(n1198) );
NAND2_X1 U861 ( .A1(KEYINPUT57), .A2(n1135), .ZN(n1200) );
NOR2_X1 U862 ( .A1(n1156), .A2(n1201), .ZN(G51) );
XOR2_X1 U863 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U864 ( .A(n1204), .B(n1155), .Z(n1203) );
NOR2_X1 U865 ( .A1(n1072), .A2(n1161), .ZN(n1204) );
NAND2_X1 U866 ( .A1(G902), .A2(n1205), .ZN(n1161) );
NAND3_X1 U867 ( .A1(n1059), .A2(n1065), .A3(n1061), .ZN(n1205) );
INV_X1 U868 ( .A(n1150), .ZN(n1061) );
NAND4_X1 U869 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1150) );
AND4_X1 U870 ( .A1(n1058), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1209) );
NAND3_X1 U871 ( .A1(n1213), .A2(n1070), .A3(n1214), .ZN(n1058) );
NOR2_X1 U872 ( .A1(n1175), .A2(n1215), .ZN(n1208) );
NOR3_X1 U873 ( .A1(n1216), .A2(n1217), .A3(n1076), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1218), .A2(n1219), .A3(n1070), .ZN(n1216) );
NAND2_X1 U875 ( .A1(KEYINPUT50), .A2(n1220), .ZN(n1219) );
NAND2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
INV_X1 U877 ( .A(KEYINPUT50), .ZN(n1222) );
NAND3_X1 U878 ( .A1(n1223), .A2(n1097), .A3(n1092), .ZN(n1221) );
AND3_X1 U879 ( .A1(n1214), .A2(n1070), .A3(n1224), .ZN(n1175) );
AND4_X1 U880 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1059) );
NOR2_X1 U881 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NOR2_X1 U882 ( .A1(n1110), .A2(n1231), .ZN(n1230) );
NOR2_X1 U883 ( .A1(n1232), .A2(n1233), .ZN(n1110) );
NOR3_X1 U884 ( .A1(n1234), .A2(n1104), .A3(n1097), .ZN(n1229) );
NOR2_X1 U885 ( .A1(n1224), .A2(n1213), .ZN(n1104) );
XOR2_X1 U886 ( .A(n1235), .B(KEYINPUT24), .Z(n1202) );
NAND2_X1 U887 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U888 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
OR2_X1 U889 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U890 ( .A(KEYINPUT52), .B(n1242), .Z(n1236) );
NOR3_X1 U891 ( .A1(n1238), .A2(n1241), .A3(n1240), .ZN(n1242) );
XOR2_X1 U892 ( .A(n1243), .B(KEYINPUT46), .Z(n1240) );
NAND2_X1 U893 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NOR2_X1 U894 ( .A1(n1245), .A2(n1244), .ZN(n1241) );
NOR2_X1 U895 ( .A1(n1119), .A2(G952), .ZN(n1156) );
XNOR2_X1 U896 ( .A(n1246), .B(n1247), .ZN(G48) );
NOR4_X1 U897 ( .A1(KEYINPUT36), .A2(n1097), .A3(n1248), .A4(n1234), .ZN(n1247) );
NAND2_X1 U898 ( .A1(n1249), .A2(n1250), .ZN(G45) );
NAND2_X1 U899 ( .A1(G143), .A2(n1065), .ZN(n1250) );
XOR2_X1 U900 ( .A(KEYINPUT23), .B(n1251), .Z(n1249) );
NOR2_X1 U901 ( .A1(G143), .A2(n1065), .ZN(n1251) );
NAND3_X1 U902 ( .A1(n1233), .A2(n1252), .A3(n1253), .ZN(n1065) );
NOR3_X1 U903 ( .A1(n1097), .A2(n1217), .A3(n1076), .ZN(n1253) );
INV_X1 U904 ( .A(n1254), .ZN(n1097) );
XNOR2_X1 U905 ( .A(n1135), .B(n1255), .ZN(G42) );
NOR2_X1 U906 ( .A1(n1231), .A2(n1256), .ZN(n1255) );
XOR2_X1 U907 ( .A(KEYINPUT2), .B(n1232), .Z(n1256) );
XNOR2_X1 U908 ( .A(G137), .B(n1226), .ZN(G39) );
NAND3_X1 U909 ( .A1(n1257), .A2(n1095), .A3(n1102), .ZN(n1226) );
NAND2_X1 U910 ( .A1(n1258), .A2(n1259), .ZN(G36) );
NAND2_X1 U911 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U912 ( .A(n1227), .B(KEYINPUT11), .Z(n1260) );
NAND2_X1 U913 ( .A1(n1262), .A2(G134), .ZN(n1258) );
XNOR2_X1 U914 ( .A(KEYINPUT33), .B(n1227), .ZN(n1262) );
NAND4_X1 U915 ( .A1(n1102), .A2(n1233), .A3(n1252), .A4(n1213), .ZN(n1227) );
XNOR2_X1 U916 ( .A(n1263), .B(n1264), .ZN(G33) );
NOR2_X1 U917 ( .A1(n1265), .A2(n1231), .ZN(n1264) );
NAND3_X1 U918 ( .A1(n1224), .A2(n1252), .A3(n1102), .ZN(n1231) );
AND2_X1 U919 ( .A1(n1099), .A2(n1082), .ZN(n1102) );
NAND2_X1 U920 ( .A1(n1266), .A2(n1267), .ZN(G30) );
NAND2_X1 U921 ( .A1(G128), .A2(n1268), .ZN(n1267) );
XOR2_X1 U922 ( .A(KEYINPUT49), .B(n1269), .Z(n1266) );
NOR2_X1 U923 ( .A1(G128), .A2(n1268), .ZN(n1269) );
NAND3_X1 U924 ( .A1(n1213), .A2(n1254), .A3(n1257), .ZN(n1268) );
INV_X1 U925 ( .A(n1234), .ZN(n1257) );
NAND3_X1 U926 ( .A1(n1270), .A2(n1271), .A3(n1252), .ZN(n1234) );
AND2_X1 U927 ( .A1(n1114), .A2(n1272), .ZN(n1252) );
XNOR2_X1 U928 ( .A(G101), .B(n1206), .ZN(G3) );
NAND3_X1 U929 ( .A1(n1233), .A2(n1214), .A3(n1095), .ZN(n1206) );
XNOR2_X1 U930 ( .A(G125), .B(n1225), .ZN(G27) );
NAND4_X1 U931 ( .A1(n1254), .A2(n1272), .A3(n1232), .A4(n1273), .ZN(n1225) );
NOR2_X1 U932 ( .A1(n1109), .A2(n1248), .ZN(n1273) );
INV_X1 U933 ( .A(n1224), .ZN(n1248) );
NAND2_X1 U934 ( .A1(n1115), .A2(n1274), .ZN(n1272) );
NAND4_X1 U935 ( .A1(G953), .A2(G902), .A3(n1127), .A4(n1275), .ZN(n1274) );
XOR2_X1 U936 ( .A(KEYINPUT55), .B(G900), .Z(n1127) );
XNOR2_X1 U937 ( .A(G122), .B(n1276), .ZN(G24) );
NAND4_X1 U938 ( .A1(n1277), .A2(n1070), .A3(n1278), .A4(n1279), .ZN(n1276) );
NOR2_X1 U939 ( .A1(n1271), .A2(n1270), .ZN(n1070) );
XNOR2_X1 U940 ( .A(G119), .B(n1207), .ZN(G21) );
NAND4_X1 U941 ( .A1(n1277), .A2(n1095), .A3(n1270), .A4(n1271), .ZN(n1207) );
XOR2_X1 U942 ( .A(n1212), .B(n1280), .Z(G18) );
NOR2_X1 U943 ( .A1(G116), .A2(KEYINPUT56), .ZN(n1280) );
NAND3_X1 U944 ( .A1(n1233), .A2(n1213), .A3(n1277), .ZN(n1212) );
NOR2_X1 U945 ( .A1(n1279), .A2(n1076), .ZN(n1213) );
INV_X1 U946 ( .A(n1278), .ZN(n1076) );
XNOR2_X1 U947 ( .A(G113), .B(n1211), .ZN(G15) );
NAND3_X1 U948 ( .A1(n1224), .A2(n1233), .A3(n1277), .ZN(n1211) );
INV_X1 U949 ( .A(n1220), .ZN(n1277) );
NAND3_X1 U950 ( .A1(n1254), .A2(n1223), .A3(n1092), .ZN(n1220) );
INV_X1 U951 ( .A(n1109), .ZN(n1092) );
NAND2_X1 U952 ( .A1(n1111), .A2(n1081), .ZN(n1109) );
INV_X1 U953 ( .A(n1265), .ZN(n1233) );
NAND2_X1 U954 ( .A1(n1281), .A2(n1271), .ZN(n1265) );
NOR2_X1 U955 ( .A1(n1278), .A2(n1217), .ZN(n1224) );
INV_X1 U956 ( .A(n1279), .ZN(n1217) );
XOR2_X1 U957 ( .A(n1210), .B(n1282), .Z(G12) );
XOR2_X1 U958 ( .A(KEYINPUT9), .B(G110), .Z(n1282) );
NAND3_X1 U959 ( .A1(n1095), .A2(n1214), .A3(n1232), .ZN(n1210) );
NOR2_X1 U960 ( .A1(n1271), .A2(n1281), .ZN(n1232) );
INV_X1 U961 ( .A(n1270), .ZN(n1281) );
XOR2_X1 U962 ( .A(n1283), .B(n1160), .Z(n1270) );
NAND2_X1 U963 ( .A1(G217), .A2(n1284), .ZN(n1160) );
NAND2_X1 U964 ( .A1(n1158), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U965 ( .A(n1286), .B(n1287), .ZN(n1158) );
XOR2_X1 U966 ( .A(KEYINPUT59), .B(G137), .Z(n1287) );
XNOR2_X1 U967 ( .A(n1288), .B(n1289), .ZN(n1286) );
NOR3_X1 U968 ( .A1(n1290), .A2(KEYINPUT5), .A3(n1291), .ZN(n1289) );
INV_X1 U969 ( .A(G221), .ZN(n1291) );
NOR2_X1 U970 ( .A1(KEYINPUT3), .A2(n1292), .ZN(n1288) );
XOR2_X1 U971 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U972 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U973 ( .A(n1245), .B(n1297), .ZN(n1296) );
XNOR2_X1 U974 ( .A(G128), .B(n1298), .ZN(n1293) );
XNOR2_X1 U975 ( .A(KEYINPUT6), .B(KEYINPUT18), .ZN(n1298) );
XNOR2_X1 U976 ( .A(n1299), .B(G472), .ZN(n1271) );
NAND2_X1 U977 ( .A1(n1300), .A2(n1285), .ZN(n1299) );
XOR2_X1 U978 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U979 ( .A(n1189), .B(n1187), .ZN(n1302) );
XNOR2_X1 U980 ( .A(n1303), .B(n1304), .ZN(n1187) );
XNOR2_X1 U981 ( .A(G113), .B(G116), .ZN(n1303) );
XOR2_X1 U982 ( .A(n1305), .B(G101), .Z(n1189) );
NAND2_X1 U983 ( .A1(n1306), .A2(G210), .ZN(n1305) );
XNOR2_X1 U984 ( .A(n1307), .B(KEYINPUT43), .ZN(n1301) );
NAND2_X1 U985 ( .A1(KEYINPUT35), .A2(n1184), .ZN(n1307) );
XNOR2_X1 U986 ( .A(n1308), .B(n1309), .ZN(n1184) );
INV_X1 U987 ( .A(n1244), .ZN(n1309) );
AND3_X1 U988 ( .A1(n1114), .A2(n1223), .A3(n1254), .ZN(n1214) );
NOR2_X1 U989 ( .A1(n1099), .A2(n1101), .ZN(n1254) );
INV_X1 U990 ( .A(n1082), .ZN(n1101) );
NAND2_X1 U991 ( .A1(G214), .A2(n1310), .ZN(n1082) );
XOR2_X1 U992 ( .A(n1311), .B(n1072), .Z(n1099) );
NAND2_X1 U993 ( .A1(G210), .A2(n1310), .ZN(n1072) );
NAND2_X1 U994 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
INV_X1 U995 ( .A(G237), .ZN(n1313) );
XNOR2_X1 U996 ( .A(G902), .B(KEYINPUT31), .ZN(n1312) );
NAND2_X1 U997 ( .A1(KEYINPUT30), .A2(n1073), .ZN(n1311) );
NAND2_X1 U998 ( .A1(n1314), .A2(n1285), .ZN(n1073) );
XOR2_X1 U999 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1000 ( .A(n1238), .B(n1317), .Z(n1316) );
NOR2_X1 U1001 ( .A1(KEYINPUT10), .A2(n1155), .ZN(n1317) );
XNOR2_X1 U1002 ( .A(n1318), .B(n1319), .ZN(n1155) );
XOR2_X1 U1003 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1004 ( .A(G101), .B(G122), .ZN(n1321) );
NAND2_X1 U1005 ( .A1(KEYINPUT28), .A2(n1322), .ZN(n1320) );
INV_X1 U1006 ( .A(G116), .ZN(n1322) );
XOR2_X1 U1007 ( .A(n1323), .B(n1324), .Z(n1318) );
XOR2_X1 U1008 ( .A(n1325), .B(n1295), .Z(n1323) );
XOR2_X1 U1009 ( .A(G110), .B(n1304), .Z(n1295) );
XOR2_X1 U1010 ( .A(G119), .B(KEYINPUT13), .Z(n1304) );
NAND2_X1 U1011 ( .A1(KEYINPUT62), .A2(n1326), .ZN(n1325) );
INV_X1 U1012 ( .A(G113), .ZN(n1326) );
NAND2_X1 U1013 ( .A1(G224), .A2(n1119), .ZN(n1238) );
NAND2_X1 U1014 ( .A1(n1327), .A2(n1328), .ZN(n1315) );
NAND2_X1 U1015 ( .A1(G125), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1016 ( .A(n1330), .B(KEYINPUT60), .Z(n1327) );
OR2_X1 U1017 ( .A1(n1329), .A2(G125), .ZN(n1330) );
XOR2_X1 U1018 ( .A(n1244), .B(KEYINPUT54), .Z(n1329) );
XOR2_X1 U1019 ( .A(G146), .B(n1331), .Z(n1244) );
NAND2_X1 U1020 ( .A1(n1115), .A2(n1332), .ZN(n1223) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1275), .A4(n1333), .ZN(n1332) );
INV_X1 U1022 ( .A(G898), .ZN(n1333) );
NAND3_X1 U1023 ( .A1(n1275), .A2(n1119), .A3(G952), .ZN(n1115) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1275) );
NOR2_X1 U1025 ( .A1(n1334), .A2(n1111), .ZN(n1114) );
XOR2_X1 U1026 ( .A(G469), .B(n1335), .Z(n1111) );
NOR2_X1 U1027 ( .A1(n1084), .A2(KEYINPUT37), .ZN(n1335) );
AND2_X1 U1028 ( .A1(n1336), .A2(n1285), .ZN(n1084) );
XOR2_X1 U1029 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1030 ( .A(n1135), .B(n1197), .ZN(n1338) );
XNOR2_X1 U1031 ( .A(n1339), .B(n1340), .ZN(n1197) );
XOR2_X1 U1032 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1033 ( .A(G110), .B(n1343), .Z(n1342) );
NOR2_X1 U1034 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1035 ( .A(n1346), .B(KEYINPUT8), .Z(n1345) );
NAND2_X1 U1036 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
INV_X1 U1037 ( .A(G101), .ZN(n1348) );
XOR2_X1 U1038 ( .A(KEYINPUT27), .B(n1324), .Z(n1347) );
AND2_X1 U1039 ( .A1(n1324), .A2(G101), .ZN(n1344) );
XOR2_X1 U1040 ( .A(G104), .B(G107), .Z(n1324) );
AND2_X1 U1041 ( .A1(n1119), .A2(G227), .ZN(n1341) );
XNOR2_X1 U1042 ( .A(n1308), .B(n1139), .ZN(n1339) );
XOR2_X1 U1043 ( .A(n1349), .B(n1350), .Z(n1139) );
NOR2_X1 U1044 ( .A1(KEYINPUT17), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1045 ( .A(G128), .B(G146), .ZN(n1349) );
XNOR2_X1 U1046 ( .A(G131), .B(n1131), .ZN(n1308) );
XOR2_X1 U1047 ( .A(G137), .B(G134), .Z(n1131) );
INV_X1 U1048 ( .A(G140), .ZN(n1135) );
XOR2_X1 U1049 ( .A(KEYINPUT41), .B(KEYINPUT40), .Z(n1337) );
XNOR2_X1 U1050 ( .A(n1081), .B(KEYINPUT21), .ZN(n1334) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1284), .ZN(n1081) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1285), .ZN(n1284) );
NOR2_X1 U1053 ( .A1(n1278), .A2(n1279), .ZN(n1095) );
NAND2_X1 U1054 ( .A1(n1083), .A2(n1352), .ZN(n1279) );
NAND2_X1 U1055 ( .A1(G475), .A2(n1077), .ZN(n1352) );
NAND2_X1 U1056 ( .A1(n1174), .A2(n1285), .ZN(n1077) );
NAND3_X1 U1057 ( .A1(n1079), .A2(n1285), .A3(n1174), .ZN(n1083) );
INV_X1 U1058 ( .A(n1170), .ZN(n1174) );
XNOR2_X1 U1059 ( .A(n1353), .B(n1354), .ZN(n1170) );
XNOR2_X1 U1060 ( .A(n1355), .B(n1356), .ZN(n1354) );
NOR2_X1 U1061 ( .A1(KEYINPUT63), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1062 ( .A1(KEYINPUT15), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1063 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
NAND2_X1 U1064 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XNOR2_X1 U1065 ( .A(n1263), .B(n1363), .ZN(n1362) );
INV_X1 U1066 ( .A(G131), .ZN(n1263) );
XNOR2_X1 U1067 ( .A(n1364), .B(n1297), .ZN(n1361) );
XOR2_X1 U1068 ( .A(n1365), .B(KEYINPUT42), .Z(n1359) );
NAND2_X1 U1069 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
XNOR2_X1 U1070 ( .A(G131), .B(n1363), .ZN(n1367) );
NOR2_X1 U1071 ( .A1(KEYINPUT53), .A2(n1368), .ZN(n1363) );
XNOR2_X1 U1072 ( .A(G143), .B(n1369), .ZN(n1368) );
NAND2_X1 U1073 ( .A1(n1306), .A2(G214), .ZN(n1369) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1306) );
XOR2_X1 U1075 ( .A(n1364), .B(n1297), .Z(n1366) );
XNOR2_X1 U1076 ( .A(n1246), .B(G140), .ZN(n1297) );
INV_X1 U1077 ( .A(G146), .ZN(n1246) );
NAND2_X1 U1078 ( .A1(KEYINPUT48), .A2(n1245), .ZN(n1364) );
INV_X1 U1079 ( .A(G125), .ZN(n1245) );
XNOR2_X1 U1080 ( .A(G104), .B(G113), .ZN(n1353) );
INV_X1 U1081 ( .A(G902), .ZN(n1285) );
INV_X1 U1082 ( .A(G475), .ZN(n1079) );
XOR2_X1 U1083 ( .A(n1370), .B(n1165), .Z(n1278) );
INV_X1 U1084 ( .A(G478), .ZN(n1165) );
OR2_X1 U1085 ( .A1(n1164), .A2(G902), .ZN(n1370) );
XNOR2_X1 U1086 ( .A(n1371), .B(n1372), .ZN(n1164) );
XOR2_X1 U1087 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1088 ( .A(n1357), .B(G116), .ZN(n1374) );
INV_X1 U1089 ( .A(G122), .ZN(n1357) );
XNOR2_X1 U1090 ( .A(KEYINPUT25), .B(n1261), .ZN(n1373) );
INV_X1 U1091 ( .A(G134), .ZN(n1261) );
XOR2_X1 U1092 ( .A(n1375), .B(n1331), .Z(n1371) );
XNOR2_X1 U1093 ( .A(G128), .B(n1351), .ZN(n1331) );
INV_X1 U1094 ( .A(G143), .ZN(n1351) );
XOR2_X1 U1095 ( .A(n1376), .B(G107), .Z(n1375) );
NAND2_X1 U1096 ( .A1(G217), .A2(n1377), .ZN(n1376) );
INV_X1 U1097 ( .A(n1290), .ZN(n1377) );
NAND2_X1 U1098 ( .A1(G234), .A2(n1119), .ZN(n1290) );
INV_X1 U1099 ( .A(G953), .ZN(n1119) );
endmodule


