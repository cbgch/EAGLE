//Key = 1010110111100011111001000111001010011110000010101111111111011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;

XOR2_X1 U753 ( .A(G107), .B(n1036), .Z(G9) );
NOR2_X1 U754 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR4_X1 U756 ( .A1(G953), .A2(n1039), .A3(n1041), .A4(n1042), .ZN(n1037) );
INV_X1 U757 ( .A(n1043), .ZN(n1042) );
NOR3_X1 U758 ( .A1(n1044), .A2(KEYINPUT20), .A3(n1045), .ZN(n1041) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR4_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NOR3_X1 U761 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1049) );
NOR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1048) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR3_X1 U765 ( .A1(n1052), .A2(n1061), .A3(n1058), .ZN(n1046) );
NOR2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U767 ( .A1(n1064), .A2(n1050), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U770 ( .A1(n1069), .A2(n1051), .ZN(n1062) );
NOR2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
INV_X1 U773 ( .A(n1074), .ZN(n1044) );
AND4_X1 U774 ( .A1(n1075), .A2(n1055), .A3(n1076), .A4(n1077), .ZN(n1039) );
NOR4_X1 U775 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U777 ( .A(KEYINPUT1), .B(G472), .Z(n1083) );
NAND2_X1 U778 ( .A1(KEYINPUT49), .A2(n1084), .ZN(n1082) );
INV_X1 U779 ( .A(n1085), .ZN(n1079) );
NOR2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1076) );
XNOR2_X1 U781 ( .A(n1088), .B(KEYINPUT37), .ZN(n1087) );
XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(n1086) );
XOR2_X1 U783 ( .A(KEYINPUT10), .B(G478), .Z(n1090) );
XOR2_X1 U784 ( .A(n1091), .B(n1092), .Z(n1075) );
XOR2_X1 U785 ( .A(n1093), .B(n1094), .Z(G72) );
XOR2_X1 U786 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U787 ( .A1(n1097), .A2(n1098), .A3(KEYINPUT9), .ZN(n1096) );
OR2_X1 U788 ( .A1(n1099), .A2(G227), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1099), .ZN(n1095) );
XOR2_X1 U790 ( .A(KEYINPUT2), .B(n1101), .Z(n1100) );
NOR2_X1 U791 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XNOR2_X1 U792 ( .A(KEYINPUT46), .B(n1104), .ZN(n1103) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1098), .ZN(n1093) );
OR2_X1 U794 ( .A1(n1099), .A2(G900), .ZN(n1098) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U797 ( .A1(KEYINPUT54), .A2(n1110), .ZN(n1109) );
AND2_X1 U798 ( .A1(KEYINPUT32), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U799 ( .A(n1111), .B(n1112), .ZN(n1110) );
XOR2_X1 U800 ( .A(KEYINPUT52), .B(G131), .Z(n1112) );
XNOR2_X1 U801 ( .A(n1113), .B(n1114), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
INV_X1 U804 ( .A(G137), .ZN(n1118) );
NOR2_X1 U805 ( .A1(KEYINPUT61), .A2(n1119), .ZN(n1117) );
NOR2_X1 U806 ( .A1(KEYINPUT33), .A2(n1120), .ZN(n1119) );
NOR2_X1 U807 ( .A1(G134), .A2(n1121), .ZN(n1115) );
NOR2_X1 U808 ( .A1(n1122), .A2(KEYINPUT33), .ZN(n1121) );
NOR2_X1 U809 ( .A1(KEYINPUT61), .A2(G137), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1123), .B(G140), .Z(n1106) );
XOR2_X1 U811 ( .A(n1124), .B(n1125), .Z(G69) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U814 ( .A1(G953), .A2(n1130), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1131), .B(n1132), .Z(n1128) );
XOR2_X1 U816 ( .A(n1133), .B(KEYINPUT21), .Z(n1132) );
INV_X1 U817 ( .A(G113), .ZN(n1133) );
NAND2_X1 U818 ( .A1(n1134), .A2(n1099), .ZN(n1126) );
XOR2_X1 U819 ( .A(n1135), .B(KEYINPUT39), .Z(n1134) );
NOR2_X1 U820 ( .A1(n1136), .A2(n1099), .ZN(n1124) );
NOR2_X1 U821 ( .A1(n1137), .A2(n1130), .ZN(n1136) );
INV_X1 U822 ( .A(G898), .ZN(n1130) );
NOR2_X1 U823 ( .A1(n1138), .A2(n1139), .ZN(G66) );
NOR3_X1 U824 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
AND3_X1 U825 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
INV_X1 U826 ( .A(n1146), .ZN(n1144) );
NOR2_X1 U827 ( .A1(n1147), .A2(n1143), .ZN(n1141) );
NOR2_X1 U828 ( .A1(n1043), .A2(n1146), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1138), .A2(n1148), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1149), .B(n1150), .ZN(n1148) );
AND2_X1 U831 ( .A1(G478), .A2(n1145), .ZN(n1149) );
NOR3_X1 U832 ( .A1(n1138), .A2(n1151), .A3(n1152), .ZN(G60) );
NOR3_X1 U833 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NOR2_X1 U834 ( .A1(KEYINPUT44), .A2(n1156), .ZN(n1155) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1158), .ZN(n1151) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1159), .ZN(n1157) );
INV_X1 U837 ( .A(KEYINPUT44), .ZN(n1159) );
XOR2_X1 U838 ( .A(n1154), .B(KEYINPUT11), .Z(n1156) );
AND2_X1 U839 ( .A1(n1145), .A2(G475), .ZN(n1154) );
XOR2_X1 U840 ( .A(G104), .B(n1160), .Z(G6) );
NOR2_X1 U841 ( .A1(n1138), .A2(n1161), .ZN(G57) );
XOR2_X1 U842 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U843 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U844 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U845 ( .A(n1168), .B(KEYINPUT5), .Z(n1167) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U847 ( .A1(n1171), .A2(G210), .ZN(n1170) );
AND3_X1 U848 ( .A1(n1171), .A2(G210), .A3(G101), .ZN(n1166) );
NAND3_X1 U849 ( .A1(n1145), .A2(G472), .A3(KEYINPUT48), .ZN(n1164) );
NOR3_X1 U850 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(G54) );
AND2_X1 U851 ( .A1(KEYINPUT36), .A2(n1138), .ZN(n1174) );
NOR2_X1 U852 ( .A1(KEYINPUT36), .A2(n1040), .ZN(n1173) );
XOR2_X1 U853 ( .A(n1175), .B(n1176), .Z(n1172) );
XOR2_X1 U854 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U855 ( .A(n1179), .B(n1180), .Z(n1178) );
AND2_X1 U856 ( .A1(G469), .A2(n1145), .ZN(n1180) );
NOR2_X1 U857 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
XOR2_X1 U858 ( .A(KEYINPUT12), .B(n1183), .Z(n1182) );
AND2_X1 U859 ( .A1(n1113), .A2(n1184), .ZN(n1183) );
NOR2_X1 U860 ( .A1(n1184), .A2(n1113), .ZN(n1181) );
XOR2_X1 U861 ( .A(n1185), .B(n1186), .Z(n1175) );
XOR2_X1 U862 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U863 ( .A(G140), .B(KEYINPUT6), .ZN(n1185) );
NOR2_X1 U864 ( .A1(n1138), .A2(n1189), .ZN(G51) );
NOR2_X1 U865 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U866 ( .A(KEYINPUT31), .B(n1192), .Z(n1191) );
NOR2_X1 U867 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
AND2_X1 U868 ( .A1(n1194), .A2(n1193), .ZN(n1190) );
NAND2_X1 U869 ( .A1(n1145), .A2(n1092), .ZN(n1194) );
NOR2_X1 U870 ( .A1(n1195), .A2(n1043), .ZN(n1145) );
NOR3_X1 U871 ( .A1(n1102), .A2(n1135), .A3(n1104), .ZN(n1043) );
OR3_X1 U872 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1104) );
AND2_X1 U873 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U874 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND2_X1 U875 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND2_X1 U876 ( .A1(n1205), .A2(n1206), .ZN(n1201) );
NAND4_X1 U877 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1135) );
NOR3_X1 U878 ( .A1(n1160), .A2(n1211), .A3(n1036), .ZN(n1210) );
AND3_X1 U879 ( .A1(n1053), .A2(n1212), .A3(n1213), .ZN(n1036) );
AND3_X1 U880 ( .A1(n1212), .A2(n1054), .A3(n1213), .ZN(n1160) );
NAND2_X1 U881 ( .A1(n1214), .A2(n1215), .ZN(n1209) );
NAND3_X1 U882 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND2_X1 U883 ( .A1(n1219), .A2(n1212), .ZN(n1218) );
INV_X1 U884 ( .A(n1050), .ZN(n1212) );
OR3_X1 U885 ( .A1(n1220), .A2(KEYINPUT30), .A3(n1058), .ZN(n1217) );
NAND3_X1 U886 ( .A1(n1221), .A2(n1222), .A3(n1073), .ZN(n1216) );
NAND2_X1 U887 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U888 ( .A1(KEYINPUT30), .A2(n1204), .ZN(n1223) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1072), .ZN(n1221) );
XOR2_X1 U890 ( .A(KEYINPUT14), .B(n1053), .Z(n1225) );
INV_X1 U891 ( .A(n1226), .ZN(n1207) );
NAND3_X1 U892 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1102) );
NAND2_X1 U893 ( .A1(n1066), .A2(n1230), .ZN(n1229) );
NAND2_X1 U894 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
OR3_X1 U895 ( .A1(n1233), .A2(n1234), .A3(n1052), .ZN(n1232) );
NAND2_X1 U896 ( .A1(n1203), .A2(n1053), .ZN(n1231) );
INV_X1 U897 ( .A(n1235), .ZN(n1203) );
NOR2_X1 U898 ( .A1(n1099), .A2(G952), .ZN(n1138) );
NAND2_X1 U899 ( .A1(n1236), .A2(n1237), .ZN(G48) );
NAND2_X1 U900 ( .A1(n1196), .A2(n1238), .ZN(n1237) );
XOR2_X1 U901 ( .A(KEYINPUT55), .B(n1239), .Z(n1236) );
NOR2_X1 U902 ( .A1(n1196), .A2(n1238), .ZN(n1239) );
NOR3_X1 U903 ( .A1(n1240), .A2(n1241), .A3(n1235), .ZN(n1196) );
XOR2_X1 U904 ( .A(n1242), .B(n1197), .Z(G45) );
AND3_X1 U905 ( .A1(n1243), .A2(n1066), .A3(n1219), .ZN(n1197) );
INV_X1 U906 ( .A(n1240), .ZN(n1066) );
NAND2_X1 U907 ( .A1(KEYINPUT57), .A2(n1244), .ZN(n1242) );
XNOR2_X1 U908 ( .A(G140), .B(n1245), .ZN(G42) );
NAND4_X1 U909 ( .A1(KEYINPUT51), .A2(n1205), .A3(n1206), .A4(n1246), .ZN(n1245) );
XOR2_X1 U910 ( .A(KEYINPUT24), .B(n1199), .Z(n1246) );
XOR2_X1 U911 ( .A(G137), .B(n1247), .Z(G39) );
NOR4_X1 U912 ( .A1(KEYINPUT19), .A2(n1058), .A3(n1235), .A4(n1051), .ZN(n1247) );
INV_X1 U913 ( .A(n1199), .ZN(n1051) );
XNOR2_X1 U914 ( .A(n1248), .B(n1227), .ZN(G36) );
NAND3_X1 U915 ( .A1(n1243), .A2(n1053), .A3(n1199), .ZN(n1227) );
NAND2_X1 U916 ( .A1(KEYINPUT63), .A2(n1120), .ZN(n1248) );
NAND2_X1 U917 ( .A1(n1249), .A2(n1250), .ZN(G33) );
OR2_X1 U918 ( .A1(n1228), .A2(G131), .ZN(n1250) );
XOR2_X1 U919 ( .A(n1251), .B(KEYINPUT62), .Z(n1249) );
NAND2_X1 U920 ( .A1(G131), .A2(n1228), .ZN(n1251) );
NAND3_X1 U921 ( .A1(n1243), .A2(n1054), .A3(n1199), .ZN(n1228) );
NOR2_X1 U922 ( .A1(n1067), .A2(n1078), .ZN(n1199) );
INV_X1 U923 ( .A(n1068), .ZN(n1078) );
AND2_X1 U924 ( .A1(n1206), .A2(n1071), .ZN(n1243) );
XOR2_X1 U925 ( .A(G128), .B(n1252), .Z(G30) );
NOR3_X1 U926 ( .A1(n1235), .A2(n1253), .A3(n1254), .ZN(n1252) );
XOR2_X1 U927 ( .A(n1240), .B(KEYINPUT47), .Z(n1253) );
NAND2_X1 U928 ( .A1(n1220), .A2(n1206), .ZN(n1235) );
NOR3_X1 U929 ( .A1(n1059), .A2(n1255), .A3(n1234), .ZN(n1206) );
XOR2_X1 U930 ( .A(G101), .B(n1211), .Z(G3) );
AND3_X1 U931 ( .A1(n1071), .A2(n1213), .A3(n1204), .ZN(n1211) );
XOR2_X1 U932 ( .A(n1123), .B(n1256), .Z(G27) );
NAND3_X1 U933 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NOR3_X1 U934 ( .A1(n1233), .A2(KEYINPUT29), .A3(n1234), .ZN(n1259) );
NAND2_X1 U935 ( .A1(n1260), .A2(n1261), .ZN(n1234) );
NAND2_X1 U936 ( .A1(G900), .A2(G953), .ZN(n1261) );
INV_X1 U937 ( .A(n1205), .ZN(n1233) );
NOR3_X1 U938 ( .A1(n1241), .A2(n1072), .A3(n1073), .ZN(n1205) );
INV_X1 U939 ( .A(n1262), .ZN(n1073) );
XOR2_X1 U940 ( .A(n1052), .B(KEYINPUT59), .Z(n1258) );
XOR2_X1 U941 ( .A(n1240), .B(KEYINPUT60), .Z(n1257) );
XNOR2_X1 U942 ( .A(G122), .B(n1263), .ZN(G24) );
NAND4_X1 U943 ( .A1(n1264), .A2(n1055), .A3(n1265), .A4(n1219), .ZN(n1263) );
AND2_X1 U944 ( .A1(n1266), .A2(n1267), .ZN(n1219) );
XNOR2_X1 U945 ( .A(KEYINPUT18), .B(n1088), .ZN(n1266) );
NOR2_X1 U946 ( .A1(n1268), .A2(n1050), .ZN(n1265) );
NAND2_X1 U947 ( .A1(n1072), .A2(n1262), .ZN(n1050) );
INV_X1 U948 ( .A(n1052), .ZN(n1055) );
XOR2_X1 U949 ( .A(n1240), .B(KEYINPUT8), .Z(n1264) );
XOR2_X1 U950 ( .A(n1269), .B(n1270), .Z(G21) );
NAND3_X1 U951 ( .A1(n1204), .A2(n1220), .A3(n1214), .ZN(n1270) );
NOR2_X1 U952 ( .A1(n1262), .A2(n1072), .ZN(n1220) );
INV_X1 U953 ( .A(n1224), .ZN(n1072) );
XOR2_X1 U954 ( .A(G116), .B(n1271), .Z(G18) );
NOR2_X1 U955 ( .A1(n1254), .A2(n1272), .ZN(n1271) );
INV_X1 U956 ( .A(n1053), .ZN(n1254) );
NOR2_X1 U957 ( .A1(n1088), .A2(n1273), .ZN(n1053) );
XOR2_X1 U958 ( .A(G113), .B(n1226), .Z(G15) );
NOR2_X1 U959 ( .A1(n1272), .A2(n1241), .ZN(n1226) );
INV_X1 U960 ( .A(n1054), .ZN(n1241) );
NAND2_X1 U961 ( .A1(n1274), .A2(n1275), .ZN(n1054) );
OR2_X1 U962 ( .A1(n1058), .A2(KEYINPUT18), .ZN(n1275) );
INV_X1 U963 ( .A(n1204), .ZN(n1058) );
NAND3_X1 U964 ( .A1(n1273), .A2(n1088), .A3(KEYINPUT18), .ZN(n1274) );
INV_X1 U965 ( .A(n1267), .ZN(n1273) );
NAND2_X1 U966 ( .A1(n1214), .A2(n1071), .ZN(n1272) );
NOR2_X1 U967 ( .A1(n1224), .A2(n1262), .ZN(n1071) );
NOR3_X1 U968 ( .A1(n1240), .A2(n1268), .A3(n1052), .ZN(n1214) );
NAND2_X1 U969 ( .A1(n1059), .A2(n1060), .ZN(n1052) );
XOR2_X1 U970 ( .A(n1187), .B(n1208), .Z(G12) );
NAND4_X1 U971 ( .A1(n1204), .A2(n1213), .A3(n1262), .A4(n1224), .ZN(n1208) );
NAND3_X1 U972 ( .A1(n1276), .A2(n1277), .A3(n1085), .ZN(n1224) );
NAND2_X1 U973 ( .A1(n1140), .A2(n1146), .ZN(n1085) );
NAND2_X1 U974 ( .A1(n1080), .A2(n1278), .ZN(n1277) );
INV_X1 U975 ( .A(KEYINPUT41), .ZN(n1278) );
NOR2_X1 U976 ( .A1(n1146), .A2(n1140), .ZN(n1080) );
NAND2_X1 U977 ( .A1(G217), .A2(n1279), .ZN(n1146) );
NAND2_X1 U978 ( .A1(KEYINPUT41), .A2(n1140), .ZN(n1276) );
NOR2_X1 U979 ( .A1(n1143), .A2(G902), .ZN(n1140) );
XNOR2_X1 U980 ( .A(n1280), .B(n1281), .ZN(n1143) );
XOR2_X1 U981 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U982 ( .A(n1284), .B(n1285), .Z(n1283) );
NOR2_X1 U983 ( .A1(KEYINPUT34), .A2(n1286), .ZN(n1285) );
XOR2_X1 U984 ( .A(G110), .B(n1287), .Z(n1286) );
XOR2_X1 U985 ( .A(G128), .B(G119), .Z(n1287) );
NAND2_X1 U986 ( .A1(n1288), .A2(G221), .ZN(n1284) );
XOR2_X1 U987 ( .A(n1123), .B(n1289), .Z(n1280) );
XOR2_X1 U988 ( .A(KEYINPUT28), .B(G137), .Z(n1289) );
XOR2_X1 U989 ( .A(n1084), .B(G472), .Z(n1262) );
NAND2_X1 U990 ( .A1(n1290), .A2(n1195), .ZN(n1084) );
XOR2_X1 U991 ( .A(n1162), .B(n1291), .Z(n1290) );
XOR2_X1 U992 ( .A(n1169), .B(n1292), .Z(n1291) );
NAND3_X1 U993 ( .A1(n1171), .A2(G210), .A3(n1293), .ZN(n1292) );
XNOR2_X1 U994 ( .A(KEYINPUT4), .B(KEYINPUT27), .ZN(n1293) );
XOR2_X1 U995 ( .A(n1294), .B(n1295), .Z(n1162) );
XNOR2_X1 U996 ( .A(G116), .B(n1296), .ZN(n1295) );
NAND2_X1 U997 ( .A1(KEYINPUT7), .A2(n1269), .ZN(n1296) );
INV_X1 U998 ( .A(G119), .ZN(n1269) );
XNOR2_X1 U999 ( .A(n1297), .B(n1298), .ZN(n1294) );
NOR4_X1 U1000 ( .A1(n1240), .A2(n1268), .A3(n1059), .A4(n1255), .ZN(n1213) );
INV_X1 U1001 ( .A(n1060), .ZN(n1255) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1279), .ZN(n1060) );
NAND2_X1 U1003 ( .A1(G234), .A2(n1195), .ZN(n1279) );
XOR2_X1 U1004 ( .A(n1299), .B(G469), .Z(n1059) );
NAND2_X1 U1005 ( .A1(n1300), .A2(n1195), .ZN(n1299) );
XOR2_X1 U1006 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1007 ( .A(n1177), .B(n1113), .Z(n1302) );
XOR2_X1 U1008 ( .A(n1238), .B(n1303), .Z(n1113) );
XOR2_X1 U1009 ( .A(n1298), .B(KEYINPUT50), .Z(n1177) );
XNOR2_X1 U1010 ( .A(n1304), .B(n1305), .ZN(n1298) );
NOR2_X1 U1011 ( .A1(KEYINPUT23), .A2(G131), .ZN(n1305) );
XOR2_X1 U1012 ( .A(n1120), .B(G137), .Z(n1304) );
INV_X1 U1013 ( .A(G134), .ZN(n1120) );
XOR2_X1 U1014 ( .A(n1306), .B(n1307), .Z(n1301) );
XOR2_X1 U1015 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1016 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1017 ( .A(KEYINPUT13), .B(n1312), .Z(n1311) );
NOR2_X1 U1018 ( .A1(G140), .A2(n1187), .ZN(n1312) );
AND2_X1 U1019 ( .A1(n1187), .A2(G140), .ZN(n1310) );
NOR2_X1 U1020 ( .A1(KEYINPUT22), .A2(n1188), .ZN(n1308) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1099), .ZN(n1188) );
NOR2_X1 U1022 ( .A1(KEYINPUT58), .A2(n1184), .ZN(n1306) );
XNOR2_X1 U1023 ( .A(n1313), .B(n1314), .ZN(n1184) );
XOR2_X1 U1024 ( .A(n1169), .B(KEYINPUT0), .Z(n1313) );
INV_X1 U1025 ( .A(G101), .ZN(n1169) );
NAND2_X1 U1026 ( .A1(n1260), .A2(n1315), .ZN(n1268) );
NAND2_X1 U1027 ( .A1(G898), .A2(G953), .ZN(n1315) );
AND3_X1 U1028 ( .A1(n1074), .A2(n1040), .A3(n1316), .ZN(n1260) );
NAND2_X1 U1029 ( .A1(G953), .A2(n1195), .ZN(n1316) );
OR2_X1 U1030 ( .A1(G952), .A2(G953), .ZN(n1040) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1074) );
NAND2_X1 U1032 ( .A1(n1067), .A2(n1068), .ZN(n1240) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1317), .ZN(n1068) );
XOR2_X1 U1034 ( .A(n1318), .B(n1092), .Z(n1067) );
AND2_X1 U1035 ( .A1(G210), .A2(n1317), .ZN(n1092) );
NAND2_X1 U1036 ( .A1(n1319), .A2(n1195), .ZN(n1317) );
INV_X1 U1037 ( .A(G237), .ZN(n1319) );
NAND2_X1 U1038 ( .A1(KEYINPUT17), .A2(n1091), .ZN(n1318) );
NAND2_X1 U1039 ( .A1(n1320), .A2(n1195), .ZN(n1091) );
XOR2_X1 U1040 ( .A(n1193), .B(n1321), .Z(n1320) );
XNOR2_X1 U1041 ( .A(KEYINPUT42), .B(KEYINPUT26), .ZN(n1321) );
XOR2_X1 U1042 ( .A(n1322), .B(n1323), .Z(n1193) );
XOR2_X1 U1043 ( .A(G125), .B(n1324), .Z(n1323) );
NOR2_X1 U1044 ( .A1(G953), .A2(n1137), .ZN(n1324) );
INV_X1 U1045 ( .A(G224), .ZN(n1137) );
XOR2_X1 U1046 ( .A(n1131), .B(n1297), .Z(n1322) );
XOR2_X1 U1047 ( .A(n1325), .B(n1303), .Z(n1297) );
XOR2_X1 U1048 ( .A(n1326), .B(G113), .Z(n1325) );
NAND2_X1 U1049 ( .A1(KEYINPUT25), .A2(n1238), .ZN(n1326) );
XOR2_X1 U1050 ( .A(n1327), .B(n1328), .Z(n1131) );
XNOR2_X1 U1051 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1052 ( .A1(KEYINPUT3), .A2(n1314), .ZN(n1330) );
XNOR2_X1 U1053 ( .A(G104), .B(G107), .ZN(n1314) );
NAND2_X1 U1054 ( .A1(KEYINPUT53), .A2(G110), .ZN(n1329) );
XOR2_X1 U1055 ( .A(n1331), .B(n1332), .Z(n1327) );
XOR2_X1 U1056 ( .A(G122), .B(G101), .Z(n1332) );
NAND2_X1 U1057 ( .A1(n1333), .A2(KEYINPUT15), .ZN(n1331) );
XNOR2_X1 U1058 ( .A(G116), .B(n1334), .ZN(n1333) );
NOR2_X1 U1059 ( .A1(G119), .A2(KEYINPUT45), .ZN(n1334) );
NOR2_X1 U1060 ( .A1(n1267), .A2(n1088), .ZN(n1204) );
XNOR2_X1 U1061 ( .A(n1335), .B(G475), .ZN(n1088) );
NAND2_X1 U1062 ( .A1(n1153), .A2(n1195), .ZN(n1335) );
INV_X1 U1063 ( .A(G902), .ZN(n1195) );
INV_X1 U1064 ( .A(n1158), .ZN(n1153) );
XOR2_X1 U1065 ( .A(n1336), .B(KEYINPUT56), .Z(n1158) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1067 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1068 ( .A(G122), .B(G113), .Z(n1340) );
XOR2_X1 U1069 ( .A(G143), .B(G131), .Z(n1339) );
XOR2_X1 U1070 ( .A(n1341), .B(n1342), .Z(n1337) );
XOR2_X1 U1071 ( .A(n1343), .B(n1282), .Z(n1342) );
XOR2_X1 U1072 ( .A(n1238), .B(G140), .Z(n1282) );
INV_X1 U1073 ( .A(G146), .ZN(n1238) );
NAND2_X1 U1074 ( .A1(KEYINPUT16), .A2(n1123), .ZN(n1343) );
INV_X1 U1075 ( .A(G125), .ZN(n1123) );
XOR2_X1 U1076 ( .A(n1344), .B(G104), .Z(n1341) );
NAND2_X1 U1077 ( .A1(n1171), .A2(G214), .ZN(n1344) );
NOR2_X1 U1078 ( .A1(G237), .A2(G953), .ZN(n1171) );
NAND2_X1 U1079 ( .A1(n1345), .A2(n1346), .ZN(n1267) );
NAND2_X1 U1080 ( .A1(G478), .A2(n1089), .ZN(n1346) );
XOR2_X1 U1081 ( .A(KEYINPUT38), .B(n1347), .Z(n1345) );
NOR2_X1 U1082 ( .A1(G478), .A2(n1089), .ZN(n1347) );
NAND2_X1 U1083 ( .A1(n1150), .A2(n1348), .ZN(n1089) );
XOR2_X1 U1084 ( .A(KEYINPUT35), .B(G902), .Z(n1348) );
XOR2_X1 U1085 ( .A(n1349), .B(n1350), .Z(n1150) );
XOR2_X1 U1086 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1087 ( .A(n1353), .B(n1354), .ZN(n1352) );
NOR2_X1 U1088 ( .A1(KEYINPUT43), .A2(n1303), .ZN(n1354) );
XOR2_X1 U1089 ( .A(G128), .B(n1244), .Z(n1303) );
INV_X1 U1090 ( .A(G143), .ZN(n1244) );
NOR2_X1 U1091 ( .A1(G107), .A2(KEYINPUT40), .ZN(n1353) );
NAND2_X1 U1092 ( .A1(G217), .A2(n1288), .ZN(n1351) );
AND2_X1 U1093 ( .A1(G234), .A2(n1099), .ZN(n1288) );
INV_X1 U1094 ( .A(G953), .ZN(n1099) );
XNOR2_X1 U1095 ( .A(G116), .B(n1355), .ZN(n1349) );
XOR2_X1 U1096 ( .A(G134), .B(G122), .Z(n1355) );
INV_X1 U1097 ( .A(G110), .ZN(n1187) );
endmodule


