//Key = 0000010101100101100010001010011001011101010110101101001011011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U744 ( .A(G107), .B(n1033), .Z(G9) );
NOR2_X1 U745 ( .A1(KEYINPUT3), .A2(n1034), .ZN(n1033) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U747 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U750 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1048) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR3_X1 U757 ( .A1(n1057), .A2(n1060), .A3(n1051), .ZN(n1043) );
NOR2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U759 ( .A1(n1063), .A2(n1045), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1047), .ZN(n1061) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR3_X1 U764 ( .A1(n1040), .A2(G952), .A3(n1037), .ZN(n1035) );
AND4_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1037) );
NOR4_X1 U766 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1075) );
NAND2_X1 U768 ( .A1(KEYINPUT5), .A2(n1081), .ZN(n1079) );
NOR3_X1 U769 ( .A1(n1082), .A2(n1083), .A3(n1067), .ZN(n1073) );
NOR3_X1 U770 ( .A1(n1084), .A2(KEYINPUT4), .A3(n1085), .ZN(n1082) );
INV_X1 U771 ( .A(n1086), .ZN(n1085) );
NAND2_X1 U772 ( .A1(n1087), .A2(n1088), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NAND2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
OR2_X1 U775 ( .A1(n1084), .A2(KEYINPUT4), .ZN(n1091) );
NAND2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1089) );
NAND2_X1 U777 ( .A1(G478), .A2(n1095), .ZN(n1071) );
XOR2_X1 U778 ( .A(n1096), .B(n1097), .Z(G72) );
NOR2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR3_X1 U780 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
XOR2_X1 U781 ( .A(KEYINPUT12), .B(n1103), .Z(n1102) );
NOR2_X1 U782 ( .A1(n1104), .A2(G953), .ZN(n1103) );
NOR2_X1 U783 ( .A1(G900), .A2(n1105), .ZN(n1101) );
INV_X1 U784 ( .A(n1106), .ZN(n1100) );
NOR3_X1 U785 ( .A1(n1106), .A2(G953), .A3(n1104), .ZN(n1098) );
XNOR2_X1 U786 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U787 ( .A1(KEYINPUT2), .A2(n1109), .ZN(n1108) );
XNOR2_X1 U788 ( .A(n1110), .B(G125), .ZN(n1109) );
NAND2_X1 U789 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
NAND2_X1 U790 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U791 ( .A(KEYINPUT62), .B(n1115), .Z(n1111) );
NOR2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(n1115) );
AND2_X1 U793 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U795 ( .A(G134), .B(n1120), .ZN(n1118) );
NAND2_X1 U796 ( .A1(n1121), .A2(G131), .ZN(n1116) );
XNOR2_X1 U797 ( .A(n1120), .B(n1122), .ZN(n1121) );
INV_X1 U798 ( .A(G134), .ZN(n1122) );
NAND2_X1 U799 ( .A1(KEYINPUT24), .A2(n1123), .ZN(n1120) );
NAND3_X1 U800 ( .A1(G953), .A2(n1124), .A3(KEYINPUT51), .ZN(n1096) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1124) );
XOR2_X1 U802 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U803 ( .A1(n1127), .A2(n1105), .ZN(n1126) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1130), .A2(n1105), .ZN(n1129) );
XNOR2_X1 U807 ( .A(n1131), .B(n1132), .ZN(n1130) );
NAND3_X1 U808 ( .A1(G898), .A2(n1132), .A3(G953), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U810 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U811 ( .A1(n1137), .A2(G217), .ZN(n1135) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1138), .ZN(G63) );
XOR2_X1 U813 ( .A(n1139), .B(n1093), .Z(n1138) );
NAND2_X1 U814 ( .A1(n1137), .A2(G478), .ZN(n1139) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1140), .ZN(G60) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U817 ( .A(KEYINPUT7), .B(n1092), .ZN(n1142) );
NAND3_X1 U818 ( .A1(n1137), .A2(G475), .A3(KEYINPUT33), .ZN(n1141) );
XNOR2_X1 U819 ( .A(n1143), .B(n1144), .ZN(G6) );
NOR3_X1 U820 ( .A1(n1133), .A2(n1145), .A3(n1146), .ZN(G57) );
NOR2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U822 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U823 ( .A1(KEYINPUT31), .A2(n1151), .ZN(n1150) );
INV_X1 U824 ( .A(n1152), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1145) );
XOR2_X1 U826 ( .A(n1149), .B(n1155), .Z(n1154) );
NOR2_X1 U827 ( .A1(KEYINPUT31), .A2(n1152), .ZN(n1155) );
XOR2_X1 U828 ( .A(n1156), .B(n1157), .Z(n1152) );
NAND2_X1 U829 ( .A1(KEYINPUT15), .A2(n1158), .ZN(n1156) );
INV_X1 U830 ( .A(n1159), .ZN(n1158) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1149) );
XNOR2_X1 U832 ( .A(G101), .B(n1162), .ZN(n1161) );
NAND2_X1 U833 ( .A1(n1137), .A2(G472), .ZN(n1160) );
NOR2_X1 U834 ( .A1(n1133), .A2(n1163), .ZN(G54) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U836 ( .A(n1110), .B(n1166), .ZN(n1165) );
NOR2_X1 U837 ( .A1(KEYINPUT40), .A2(n1167), .ZN(n1166) );
XOR2_X1 U838 ( .A(n1168), .B(n1114), .Z(n1167) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1164) );
NAND3_X1 U840 ( .A1(n1137), .A2(G469), .A3(KEYINPUT36), .ZN(n1169) );
NOR2_X1 U841 ( .A1(n1133), .A2(n1171), .ZN(G51) );
XOR2_X1 U842 ( .A(n1172), .B(n1173), .Z(n1171) );
XNOR2_X1 U843 ( .A(n1174), .B(n1132), .ZN(n1173) );
NOR2_X1 U844 ( .A1(KEYINPUT32), .A2(n1175), .ZN(n1174) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(n1172) );
XNOR2_X1 U846 ( .A(G125), .B(n1178), .ZN(n1177) );
NAND2_X1 U847 ( .A1(n1137), .A2(n1080), .ZN(n1178) );
AND2_X1 U848 ( .A1(G902), .A2(n1039), .ZN(n1137) );
NAND2_X1 U849 ( .A1(n1131), .A2(n1104), .ZN(n1039) );
AND4_X1 U850 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1104) );
AND4_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NAND2_X1 U852 ( .A1(n1187), .A2(n1053), .ZN(n1181) );
XNOR2_X1 U853 ( .A(n1188), .B(KEYINPUT56), .ZN(n1187) );
NAND3_X1 U854 ( .A1(n1070), .A2(n1189), .A3(n1190), .ZN(n1180) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1058), .A2(n1193), .ZN(n1192) );
XNOR2_X1 U857 ( .A(KEYINPUT61), .B(n1057), .ZN(n1193) );
INV_X1 U858 ( .A(n1194), .ZN(n1057) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1059), .ZN(n1191) );
XNOR2_X1 U860 ( .A(n1194), .B(KEYINPUT39), .ZN(n1195) );
NAND3_X1 U861 ( .A1(n1196), .A2(n1197), .A3(n1194), .ZN(n1179) );
AND4_X1 U862 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1131) );
NOR4_X1 U863 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1144), .ZN(n1201) );
AND2_X1 U864 ( .A1(n1070), .A2(n1205), .ZN(n1144) );
INV_X1 U865 ( .A(n1034), .ZN(n1204) );
NAND2_X1 U866 ( .A1(n1069), .A2(n1205), .ZN(n1034) );
AND3_X1 U867 ( .A1(n1206), .A2(n1207), .A3(n1065), .ZN(n1205) );
OR2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1200) );
NAND4_X1 U869 ( .A1(n1197), .A2(n1065), .A3(n1206), .A4(n1059), .ZN(n1199) );
NAND2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1198) );
NAND2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND2_X1 U872 ( .A1(n1214), .A2(n1069), .ZN(n1213) );
XNOR2_X1 U873 ( .A(n1058), .B(KEYINPUT13), .ZN(n1214) );
NAND2_X1 U874 ( .A1(n1215), .A2(n1197), .ZN(n1212) );
NAND2_X1 U875 ( .A1(KEYINPUT44), .A2(n1159), .ZN(n1176) );
NOR2_X1 U876 ( .A1(n1105), .A2(G952), .ZN(n1133) );
XNOR2_X1 U877 ( .A(G146), .B(n1216), .ZN(G48) );
NAND2_X1 U878 ( .A1(n1188), .A2(n1053), .ZN(n1216) );
AND2_X1 U879 ( .A1(n1196), .A2(n1070), .ZN(n1188) );
XNOR2_X1 U880 ( .A(G143), .B(n1186), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1190), .A2(n1058), .A3(n1217), .A4(n1218), .ZN(n1186) );
NOR2_X1 U882 ( .A1(n1219), .A2(n1209), .ZN(n1217) );
XNOR2_X1 U883 ( .A(n1110), .B(n1220), .ZN(G42) );
NOR2_X1 U884 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
INV_X1 U885 ( .A(n1059), .ZN(n1221) );
XNOR2_X1 U886 ( .A(G137), .B(n1223), .ZN(G39) );
NAND3_X1 U887 ( .A1(n1196), .A2(n1197), .A3(n1224), .ZN(n1223) );
XNOR2_X1 U888 ( .A(n1194), .B(KEYINPUT16), .ZN(n1224) );
XNOR2_X1 U889 ( .A(G134), .B(n1185), .ZN(G36) );
NAND4_X1 U890 ( .A1(n1194), .A2(n1190), .A3(n1058), .A4(n1069), .ZN(n1185) );
XNOR2_X1 U891 ( .A(n1119), .B(n1225), .ZN(G33) );
NOR2_X1 U892 ( .A1(n1226), .A2(n1222), .ZN(n1225) );
NAND3_X1 U893 ( .A1(n1190), .A2(n1070), .A3(n1194), .ZN(n1222) );
NOR2_X1 U894 ( .A1(n1054), .A2(n1083), .ZN(n1194) );
INV_X1 U895 ( .A(n1055), .ZN(n1083) );
INV_X1 U896 ( .A(G131), .ZN(n1119) );
XNOR2_X1 U897 ( .A(G128), .B(n1184), .ZN(G30) );
NAND3_X1 U898 ( .A1(n1069), .A2(n1053), .A3(n1196), .ZN(n1184) );
AND2_X1 U899 ( .A1(n1190), .A2(n1215), .ZN(n1196) );
AND2_X1 U900 ( .A1(n1065), .A2(n1227), .ZN(n1190) );
XNOR2_X1 U901 ( .A(G101), .B(n1228), .ZN(G3) );
NAND2_X1 U902 ( .A1(n1229), .A2(n1053), .ZN(n1228) );
XOR2_X1 U903 ( .A(n1208), .B(KEYINPUT9), .Z(n1229) );
NAND4_X1 U904 ( .A1(n1197), .A2(n1058), .A3(n1065), .A4(n1230), .ZN(n1208) );
XNOR2_X1 U905 ( .A(n1231), .B(n1183), .ZN(G27) );
NAND4_X1 U906 ( .A1(n1070), .A2(n1232), .A3(n1233), .A4(n1059), .ZN(n1183) );
AND2_X1 U907 ( .A1(n1227), .A2(n1053), .ZN(n1233) );
NAND2_X1 U908 ( .A1(n1234), .A2(n1042), .ZN(n1227) );
NAND4_X1 U909 ( .A1(G953), .A2(G902), .A3(n1235), .A4(n1236), .ZN(n1234) );
INV_X1 U910 ( .A(G900), .ZN(n1236) );
NOR2_X1 U911 ( .A1(KEYINPUT58), .A2(n1237), .ZN(n1231) );
XNOR2_X1 U912 ( .A(G125), .B(KEYINPUT38), .ZN(n1237) );
XNOR2_X1 U913 ( .A(n1203), .B(n1238), .ZN(G24) );
NAND2_X1 U914 ( .A1(KEYINPUT26), .A2(G122), .ZN(n1238) );
NOR4_X1 U915 ( .A1(n1239), .A2(n1240), .A3(n1051), .A4(n1219), .ZN(n1203) );
INV_X1 U916 ( .A(n1207), .ZN(n1051) );
NAND2_X1 U917 ( .A1(n1241), .A2(n1242), .ZN(n1207) );
OR3_X1 U918 ( .A1(n1077), .A2(n1078), .A3(KEYINPUT21), .ZN(n1242) );
NAND2_X1 U919 ( .A1(KEYINPUT21), .A2(n1059), .ZN(n1241) );
XOR2_X1 U920 ( .A(G119), .B(n1243), .Z(G21) );
NOR3_X1 U921 ( .A1(n1244), .A2(n1240), .A3(n1045), .ZN(n1243) );
XOR2_X1 U922 ( .A(KEYINPUT20), .B(n1215), .Z(n1244) );
AND2_X1 U923 ( .A1(n1078), .A2(n1077), .ZN(n1215) );
XNOR2_X1 U924 ( .A(G116), .B(n1245), .ZN(G18) );
NAND4_X1 U925 ( .A1(n1058), .A2(n1069), .A3(n1206), .A4(n1246), .ZN(n1245) );
XNOR2_X1 U926 ( .A(KEYINPUT8), .B(n1047), .ZN(n1246) );
NOR2_X1 U927 ( .A1(n1218), .A2(n1219), .ZN(n1069) );
XOR2_X1 U928 ( .A(G113), .B(n1202), .Z(G15) );
AND3_X1 U929 ( .A1(n1070), .A2(n1058), .A3(n1210), .ZN(n1202) );
INV_X1 U930 ( .A(n1240), .ZN(n1210) );
NAND2_X1 U931 ( .A1(n1232), .A2(n1206), .ZN(n1240) );
INV_X1 U932 ( .A(n1047), .ZN(n1232) );
NAND2_X1 U933 ( .A1(n1066), .A2(n1247), .ZN(n1047) );
INV_X1 U934 ( .A(n1226), .ZN(n1058) );
NAND2_X1 U935 ( .A1(n1248), .A2(n1078), .ZN(n1226) );
XNOR2_X1 U936 ( .A(KEYINPUT21), .B(n1077), .ZN(n1248) );
AND2_X1 U937 ( .A1(n1218), .A2(n1249), .ZN(n1070) );
INV_X1 U938 ( .A(n1239), .ZN(n1218) );
XNOR2_X1 U939 ( .A(n1250), .B(n1251), .ZN(G12) );
NOR2_X1 U940 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NOR2_X1 U941 ( .A1(KEYINPUT45), .A2(n1254), .ZN(n1253) );
INV_X1 U942 ( .A(n1255), .ZN(n1254) );
NOR2_X1 U943 ( .A1(KEYINPUT57), .A2(n1255), .ZN(n1252) );
NAND4_X1 U944 ( .A1(n1197), .A2(n1206), .A3(n1059), .A4(n1256), .ZN(n1255) );
XOR2_X1 U945 ( .A(KEYINPUT52), .B(n1065), .Z(n1256) );
NOR2_X1 U946 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U947 ( .A(n1247), .ZN(n1067) );
NAND2_X1 U948 ( .A1(G221), .A2(n1257), .ZN(n1247) );
NAND2_X1 U949 ( .A1(G234), .A2(n1088), .ZN(n1257) );
XNOR2_X1 U950 ( .A(n1076), .B(KEYINPUT63), .ZN(n1066) );
XNOR2_X1 U951 ( .A(n1258), .B(G469), .ZN(n1076) );
NAND2_X1 U952 ( .A1(n1259), .A2(n1088), .ZN(n1258) );
XOR2_X1 U953 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U954 ( .A(n1168), .B(n1170), .Z(n1261) );
XNOR2_X1 U955 ( .A(n1250), .B(n1262), .ZN(n1170) );
AND2_X1 U956 ( .A1(n1105), .A2(G227), .ZN(n1262) );
XOR2_X1 U957 ( .A(n1263), .B(n1264), .Z(n1168) );
XOR2_X1 U958 ( .A(n1265), .B(n1157), .Z(n1264) );
NAND2_X1 U959 ( .A1(KEYINPUT37), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U960 ( .A(G107), .B(n1267), .ZN(n1263) );
NOR2_X1 U961 ( .A1(KEYINPUT42), .A2(n1143), .ZN(n1267) );
INV_X1 U962 ( .A(G104), .ZN(n1143) );
XNOR2_X1 U963 ( .A(n1268), .B(n1269), .ZN(n1260) );
XOR2_X1 U964 ( .A(KEYINPUT18), .B(n1270), .Z(n1269) );
NOR2_X1 U965 ( .A1(n1078), .A2(n1271), .ZN(n1059) );
INV_X1 U966 ( .A(n1077), .ZN(n1271) );
NAND3_X1 U967 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1077) );
OR2_X1 U968 ( .A1(n1275), .A2(n1136), .ZN(n1274) );
NAND3_X1 U969 ( .A1(n1136), .A2(n1275), .A3(n1088), .ZN(n1273) );
NAND2_X1 U970 ( .A1(G217), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U971 ( .A(n1277), .B(n1278), .ZN(n1136) );
XOR2_X1 U972 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U973 ( .A(G137), .B(n1281), .ZN(n1280) );
NOR2_X1 U974 ( .A1(KEYINPUT47), .A2(n1282), .ZN(n1281) );
XOR2_X1 U975 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U976 ( .A(G110), .B(G128), .ZN(n1283) );
NAND2_X1 U977 ( .A1(KEYINPUT29), .A2(n1285), .ZN(n1279) );
XOR2_X1 U978 ( .A(n1286), .B(n1270), .Z(n1277) );
XNOR2_X1 U979 ( .A(n1110), .B(G146), .ZN(n1270) );
NAND2_X1 U980 ( .A1(G221), .A2(n1287), .ZN(n1286) );
NAND2_X1 U981 ( .A1(G902), .A2(G217), .ZN(n1272) );
XNOR2_X1 U982 ( .A(n1288), .B(G472), .ZN(n1078) );
NAND2_X1 U983 ( .A1(n1088), .A2(n1289), .ZN(n1288) );
NAND2_X1 U984 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U985 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U986 ( .A(n1266), .B(n1294), .ZN(n1293) );
INV_X1 U987 ( .A(G101), .ZN(n1266) );
XNOR2_X1 U988 ( .A(n1295), .B(n1147), .ZN(n1292) );
INV_X1 U989 ( .A(n1153), .ZN(n1147) );
XOR2_X1 U990 ( .A(n1296), .B(KEYINPUT55), .Z(n1290) );
NAND2_X1 U991 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XNOR2_X1 U992 ( .A(n1295), .B(n1153), .ZN(n1298) );
XOR2_X1 U993 ( .A(n1299), .B(n1300), .Z(n1153) );
NOR2_X1 U994 ( .A1(KEYINPUT53), .A2(n1301), .ZN(n1300) );
NAND2_X1 U995 ( .A1(n1302), .A2(n1303), .ZN(n1295) );
NAND2_X1 U996 ( .A1(n1157), .A2(n1159), .ZN(n1303) );
XOR2_X1 U997 ( .A(KEYINPUT41), .B(n1304), .Z(n1302) );
NOR2_X1 U998 ( .A1(n1157), .A2(n1159), .ZN(n1304) );
XOR2_X1 U999 ( .A(n1305), .B(KEYINPUT49), .Z(n1157) );
NAND2_X1 U1000 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1001 ( .A1(G131), .A2(n1308), .ZN(n1307) );
XOR2_X1 U1002 ( .A(KEYINPUT59), .B(n1309), .Z(n1306) );
NOR2_X1 U1003 ( .A1(G131), .A2(n1308), .ZN(n1309) );
XNOR2_X1 U1004 ( .A(n1123), .B(G134), .ZN(n1308) );
INV_X1 U1005 ( .A(G137), .ZN(n1123) );
XNOR2_X1 U1006 ( .A(G101), .B(n1294), .ZN(n1297) );
NOR2_X1 U1007 ( .A1(KEYINPUT50), .A2(n1162), .ZN(n1294) );
NAND3_X1 U1008 ( .A1(n1310), .A2(n1105), .A3(G210), .ZN(n1162) );
AND2_X1 U1009 ( .A1(n1053), .A2(n1230), .ZN(n1206) );
NAND2_X1 U1010 ( .A1(n1042), .A2(n1311), .ZN(n1230) );
NAND4_X1 U1011 ( .A1(G953), .A2(G902), .A3(n1235), .A4(n1312), .ZN(n1311) );
INV_X1 U1012 ( .A(G898), .ZN(n1312) );
NAND3_X1 U1013 ( .A1(n1313), .A2(n1235), .A3(n1314), .ZN(n1042) );
XNOR2_X1 U1014 ( .A(G952), .B(KEYINPUT35), .ZN(n1314) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1235) );
INV_X1 U1016 ( .A(n1040), .ZN(n1313) );
XOR2_X1 U1017 ( .A(G953), .B(KEYINPUT11), .Z(n1040) );
INV_X1 U1018 ( .A(n1209), .ZN(n1053) );
NAND2_X1 U1019 ( .A1(n1054), .A2(n1055), .ZN(n1209) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1315), .ZN(n1055) );
NAND2_X1 U1021 ( .A1(n1316), .A2(n1317), .ZN(n1054) );
OR2_X1 U1022 ( .A1(n1081), .A2(n1080), .ZN(n1317) );
XOR2_X1 U1023 ( .A(n1318), .B(KEYINPUT22), .Z(n1316) );
NAND2_X1 U1024 ( .A1(n1080), .A2(n1081), .ZN(n1318) );
NAND2_X1 U1025 ( .A1(n1319), .A2(n1088), .ZN(n1081) );
XNOR2_X1 U1026 ( .A(n1132), .B(n1320), .ZN(n1319) );
XNOR2_X1 U1027 ( .A(n1321), .B(n1175), .ZN(n1320) );
NAND2_X1 U1028 ( .A1(G224), .A2(n1105), .ZN(n1175) );
NOR2_X1 U1029 ( .A1(KEYINPUT23), .A2(n1322), .ZN(n1321) );
NOR2_X1 U1030 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1031 ( .A(n1325), .B(KEYINPUT30), .Z(n1324) );
NAND2_X1 U1032 ( .A1(n1326), .A2(G125), .ZN(n1325) );
NOR2_X1 U1033 ( .A1(G125), .A2(n1326), .ZN(n1323) );
XNOR2_X1 U1034 ( .A(n1159), .B(KEYINPUT0), .ZN(n1326) );
NAND2_X1 U1035 ( .A1(n1327), .A2(n1328), .ZN(n1159) );
NAND2_X1 U1036 ( .A1(n1114), .A2(n1329), .ZN(n1328) );
INV_X1 U1037 ( .A(KEYINPUT19), .ZN(n1329) );
XOR2_X1 U1038 ( .A(G146), .B(n1268), .Z(n1114) );
NAND3_X1 U1039 ( .A1(G128), .A2(n1330), .A3(KEYINPUT19), .ZN(n1327) );
XNOR2_X1 U1040 ( .A(G146), .B(n1331), .ZN(n1330) );
XOR2_X1 U1041 ( .A(n1332), .B(n1333), .Z(n1132) );
XOR2_X1 U1042 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1043 ( .A(n1336), .B(n1337), .ZN(n1335) );
INV_X1 U1044 ( .A(n1299), .ZN(n1337) );
XOR2_X1 U1045 ( .A(G113), .B(n1284), .Z(n1299) );
XOR2_X1 U1046 ( .A(G119), .B(KEYINPUT46), .Z(n1284) );
NOR2_X1 U1047 ( .A1(KEYINPUT25), .A2(n1338), .ZN(n1336) );
XNOR2_X1 U1048 ( .A(n1301), .B(KEYINPUT10), .ZN(n1338) );
XOR2_X1 U1049 ( .A(G116), .B(KEYINPUT27), .Z(n1301) );
XNOR2_X1 U1050 ( .A(G101), .B(n1339), .ZN(n1332) );
XNOR2_X1 U1051 ( .A(n1250), .B(G104), .ZN(n1339) );
AND2_X1 U1052 ( .A1(G210), .A2(n1315), .ZN(n1080) );
NAND2_X1 U1053 ( .A1(n1088), .A2(n1310), .ZN(n1315) );
INV_X1 U1054 ( .A(n1045), .ZN(n1197) );
NAND2_X1 U1055 ( .A1(n1249), .A2(n1239), .ZN(n1045) );
XOR2_X1 U1056 ( .A(n1084), .B(n1340), .Z(n1239) );
NOR2_X1 U1057 ( .A1(KEYINPUT14), .A2(n1086), .ZN(n1340) );
NAND2_X1 U1058 ( .A1(n1088), .A2(n1092), .ZN(n1086) );
NAND2_X1 U1059 ( .A1(n1341), .A2(n1342), .ZN(n1092) );
NAND2_X1 U1060 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1061 ( .A(KEYINPUT54), .B(n1345), .Z(n1341) );
NOR2_X1 U1062 ( .A1(n1344), .A2(n1343), .ZN(n1345) );
XOR2_X1 U1063 ( .A(n1346), .B(n1347), .Z(n1343) );
XNOR2_X1 U1064 ( .A(G131), .B(n1348), .ZN(n1347) );
XOR2_X1 U1065 ( .A(KEYINPUT1), .B(G146), .Z(n1348) );
XOR2_X1 U1066 ( .A(n1349), .B(n1350), .Z(n1346) );
XNOR2_X1 U1067 ( .A(n1285), .B(n1351), .ZN(n1350) );
NOR2_X1 U1068 ( .A1(KEYINPUT34), .A2(n1352), .ZN(n1351) );
XNOR2_X1 U1069 ( .A(G143), .B(n1353), .ZN(n1352) );
AND3_X1 U1070 ( .A1(G214), .A2(n1105), .A3(n1310), .ZN(n1353) );
INV_X1 U1071 ( .A(G237), .ZN(n1310) );
INV_X1 U1072 ( .A(G953), .ZN(n1105) );
INV_X1 U1073 ( .A(G125), .ZN(n1285) );
NAND2_X1 U1074 ( .A1(KEYINPUT48), .A2(n1110), .ZN(n1349) );
INV_X1 U1075 ( .A(G140), .ZN(n1110) );
XNOR2_X1 U1076 ( .A(n1354), .B(n1355), .ZN(n1344) );
XOR2_X1 U1077 ( .A(KEYINPUT28), .B(G122), .Z(n1355) );
XNOR2_X1 U1078 ( .A(G113), .B(G104), .ZN(n1354) );
XOR2_X1 U1079 ( .A(G475), .B(KEYINPUT60), .Z(n1084) );
XNOR2_X1 U1080 ( .A(n1219), .B(KEYINPUT43), .ZN(n1249) );
XOR2_X1 U1081 ( .A(n1094), .B(n1356), .Z(n1219) );
NOR2_X1 U1082 ( .A1(KEYINPUT17), .A2(n1095), .ZN(n1356) );
NAND2_X1 U1083 ( .A1(n1093), .A2(n1088), .ZN(n1095) );
INV_X1 U1084 ( .A(G902), .ZN(n1088) );
XOR2_X1 U1085 ( .A(n1357), .B(n1358), .Z(n1093) );
NOR2_X1 U1086 ( .A1(KEYINPUT6), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1087 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1088 ( .A(n1334), .B(n1268), .ZN(n1361) );
XNOR2_X1 U1089 ( .A(G128), .B(n1331), .ZN(n1268) );
INV_X1 U1090 ( .A(G143), .ZN(n1331) );
XOR2_X1 U1091 ( .A(G107), .B(G122), .Z(n1334) );
XNOR2_X1 U1092 ( .A(G116), .B(G134), .ZN(n1360) );
NAND2_X1 U1093 ( .A1(G217), .A2(n1287), .ZN(n1357) );
NOR2_X1 U1094 ( .A1(n1276), .A2(G953), .ZN(n1287) );
INV_X1 U1095 ( .A(G234), .ZN(n1276) );
INV_X1 U1096 ( .A(G478), .ZN(n1094) );
INV_X1 U1097 ( .A(G110), .ZN(n1250) );
endmodule


