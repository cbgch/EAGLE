//Key = 0010011011101010110001001110101001110001110111001000101001000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426;

NAND3_X1 U776 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(G9) );
NAND2_X1 U777 ( .A1(KEYINPUT42), .A2(n1076), .ZN(n1075) );
NAND2_X1 U778 ( .A1(G107), .A2(n1077), .ZN(n1076) );
NAND3_X1 U779 ( .A1(n1078), .A2(n1079), .A3(G107), .ZN(n1074) );
INV_X1 U780 ( .A(KEYINPUT42), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND3_X1 U782 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1073) );
INV_X1 U783 ( .A(KEYINPUT58), .ZN(n1081) );
INV_X1 U784 ( .A(n1077), .ZN(n1080) );
NAND3_X1 U785 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1077) );
XNOR2_X1 U786 ( .A(n1086), .B(KEYINPUT63), .ZN(n1085) );
NOR2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(G75) );
NOR4_X1 U788 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
NOR2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR3_X1 U790 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1093) );
AND2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR3_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1096) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR3_X1 U795 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1105) );
NOR3_X1 U796 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
INV_X1 U797 ( .A(KEYINPUT48), .ZN(n1110) );
NOR2_X1 U798 ( .A1(KEYINPUT48), .A2(n1113), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1113), .ZN(n1103) );
NOR2_X1 U800 ( .A1(n1084), .A2(n1115), .ZN(n1114) );
XOR2_X1 U801 ( .A(KEYINPUT19), .B(n1116), .Z(n1095) );
NOR2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR3_X1 U803 ( .A1(n1118), .A2(n1119), .A3(n1102), .ZN(n1091) );
INV_X1 U804 ( .A(n1086), .ZN(n1102) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1122), .B(KEYINPUT26), .Z(n1121) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U808 ( .A1(KEYINPUT51), .A2(n1125), .ZN(n1120) );
INV_X1 U809 ( .A(n1099), .ZN(n1118) );
NAND3_X1 U810 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1089) );
NAND3_X1 U811 ( .A1(n1129), .A2(n1130), .A3(KEYINPUT51), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1099), .A2(n1086), .ZN(n1130) );
NOR3_X1 U813 ( .A1(n1113), .A2(n1106), .A3(n1100), .ZN(n1099) );
INV_X1 U814 ( .A(n1131), .ZN(n1106) );
INV_X1 U815 ( .A(n1132), .ZN(n1113) );
NOR3_X1 U816 ( .A1(n1133), .A2(G953), .A3(G952), .ZN(n1087) );
INV_X1 U817 ( .A(n1126), .ZN(n1133) );
NAND4_X1 U818 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1126) );
NOR4_X1 U819 ( .A1(n1094), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1137) );
XNOR2_X1 U820 ( .A(n1141), .B(n1142), .ZN(n1140) );
XNOR2_X1 U821 ( .A(n1143), .B(n1144), .ZN(n1139) );
XNOR2_X1 U822 ( .A(G475), .B(KEYINPUT11), .ZN(n1144) );
AND3_X1 U823 ( .A1(n1145), .A2(n1146), .A3(n1111), .ZN(n1136) );
XNOR2_X1 U824 ( .A(KEYINPUT44), .B(n1147), .ZN(n1134) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(G72) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U827 ( .A1(G953), .A2(n1152), .ZN(n1151) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1152) );
NAND2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NAND2_X1 U830 ( .A1(G953), .A2(n1155), .ZN(n1154) );
XOR2_X1 U831 ( .A(n1156), .B(n1157), .Z(n1153) );
XNOR2_X1 U832 ( .A(G131), .B(n1158), .ZN(n1157) );
NAND2_X1 U833 ( .A1(KEYINPUT2), .A2(n1159), .ZN(n1158) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1156) );
AND2_X1 U835 ( .A1(n1162), .A2(n1127), .ZN(n1148) );
NAND2_X1 U836 ( .A1(n1163), .A2(n1164), .ZN(G69) );
NAND3_X1 U837 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U839 ( .A1(KEYINPUT25), .A2(n1170), .ZN(n1168) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1163) );
NAND2_X1 U841 ( .A1(n1165), .A2(n1166), .ZN(n1172) );
XNOR2_X1 U842 ( .A(KEYINPUT7), .B(G953), .ZN(n1165) );
XOR2_X1 U843 ( .A(n1173), .B(n1169), .Z(n1171) );
AND2_X1 U844 ( .A1(n1174), .A2(n1175), .ZN(n1169) );
NAND2_X1 U845 ( .A1(G953), .A2(n1176), .ZN(n1175) );
NAND2_X1 U846 ( .A1(KEYINPUT25), .A2(n1177), .ZN(n1173) );
XNOR2_X1 U847 ( .A(KEYINPUT46), .B(n1170), .ZN(n1177) );
NAND3_X1 U848 ( .A1(n1178), .A2(n1174), .A3(n1179), .ZN(n1170) );
INV_X1 U849 ( .A(n1180), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1181), .A2(n1182), .ZN(G66) );
NOR3_X1 U851 ( .A1(n1141), .A2(n1183), .A3(n1184), .ZN(n1182) );
NOR3_X1 U852 ( .A1(n1185), .A2(n1142), .A3(n1186), .ZN(n1184) );
INV_X1 U853 ( .A(n1187), .ZN(n1185) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1187), .ZN(n1183) );
NOR2_X1 U855 ( .A1(n1189), .A2(n1142), .ZN(n1188) );
NOR2_X1 U856 ( .A1(n1181), .A2(n1190), .ZN(G63) );
XOR2_X1 U857 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND3_X1 U858 ( .A1(n1193), .A2(n1194), .A3(G478), .ZN(n1191) );
NAND2_X1 U859 ( .A1(n1186), .A2(n1195), .ZN(n1194) );
INV_X1 U860 ( .A(KEYINPUT60), .ZN(n1195) );
NAND2_X1 U861 ( .A1(KEYINPUT60), .A2(n1196), .ZN(n1193) );
NAND2_X1 U862 ( .A1(n1189), .A2(G902), .ZN(n1196) );
NOR2_X1 U863 ( .A1(n1181), .A2(n1197), .ZN(G60) );
NOR3_X1 U864 ( .A1(n1143), .A2(n1198), .A3(n1199), .ZN(n1197) );
NOR3_X1 U865 ( .A1(n1200), .A2(n1201), .A3(n1186), .ZN(n1199) );
INV_X1 U866 ( .A(n1202), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1203), .A2(n1202), .ZN(n1198) );
NOR2_X1 U868 ( .A1(n1189), .A2(n1201), .ZN(n1203) );
INV_X1 U869 ( .A(G475), .ZN(n1201) );
XOR2_X1 U870 ( .A(G104), .B(n1204), .Z(G6) );
NOR2_X1 U871 ( .A1(n1125), .A2(n1205), .ZN(n1204) );
NOR2_X1 U872 ( .A1(n1181), .A2(n1206), .ZN(G57) );
XOR2_X1 U873 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U874 ( .A(n1209), .B(n1210), .ZN(n1208) );
XOR2_X1 U875 ( .A(n1211), .B(n1212), .Z(n1207) );
NOR2_X1 U876 ( .A1(n1213), .A2(n1186), .ZN(n1212) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
XOR2_X1 U878 ( .A(n1216), .B(KEYINPUT22), .Z(n1214) );
NOR2_X1 U879 ( .A1(n1181), .A2(n1217), .ZN(G54) );
XOR2_X1 U880 ( .A(n1218), .B(n1219), .Z(n1217) );
XNOR2_X1 U881 ( .A(n1220), .B(n1210), .ZN(n1219) );
XOR2_X1 U882 ( .A(n1221), .B(n1222), .Z(n1218) );
NOR2_X1 U883 ( .A1(KEYINPUT3), .A2(n1223), .ZN(n1222) );
XOR2_X1 U884 ( .A(n1224), .B(n1225), .Z(n1221) );
NOR2_X1 U885 ( .A1(n1226), .A2(n1186), .ZN(n1225) );
NOR2_X1 U886 ( .A1(n1181), .A2(n1227), .ZN(G51) );
XOR2_X1 U887 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U888 ( .A1(n1230), .A2(n1186), .ZN(n1229) );
NAND2_X1 U889 ( .A1(G902), .A2(n1090), .ZN(n1186) );
INV_X1 U890 ( .A(n1189), .ZN(n1090) );
NOR2_X1 U891 ( .A1(n1162), .A2(n1166), .ZN(n1189) );
NAND4_X1 U892 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1166) );
NOR4_X1 U893 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1234) );
INV_X1 U894 ( .A(n1239), .ZN(n1236) );
NAND2_X1 U895 ( .A1(n1240), .A2(n1241), .ZN(n1233) );
NAND2_X1 U896 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XNOR2_X1 U897 ( .A(n1115), .B(KEYINPUT20), .ZN(n1242) );
NAND3_X1 U898 ( .A1(n1084), .A2(n1086), .A3(n1083), .ZN(n1232) );
NAND2_X1 U899 ( .A1(n1129), .A2(n1244), .ZN(n1231) );
XNOR2_X1 U900 ( .A(KEYINPUT49), .B(n1205), .ZN(n1244) );
NAND4_X1 U901 ( .A1(n1115), .A2(n1086), .A3(n1245), .A4(n1246), .ZN(n1205) );
NAND4_X1 U902 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1162) );
NOR4_X1 U903 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
INV_X1 U904 ( .A(n1255), .ZN(n1251) );
NAND2_X1 U905 ( .A1(n1129), .A2(n1256), .ZN(n1249) );
NAND2_X1 U906 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND3_X1 U907 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
NAND2_X1 U908 ( .A1(n1132), .A2(n1262), .ZN(n1257) );
NAND3_X1 U909 ( .A1(n1261), .A2(n1084), .A3(n1263), .ZN(n1247) );
XNOR2_X1 U910 ( .A(n1264), .B(KEYINPUT57), .ZN(n1263) );
INV_X1 U911 ( .A(n1265), .ZN(n1261) );
INV_X1 U912 ( .A(G210), .ZN(n1230) );
NOR2_X1 U913 ( .A1(n1266), .A2(n1267), .ZN(n1228) );
XOR2_X1 U914 ( .A(KEYINPUT59), .B(n1268), .Z(n1267) );
AND2_X1 U915 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NOR2_X1 U916 ( .A1(n1270), .A2(n1269), .ZN(n1266) );
NAND2_X1 U917 ( .A1(n1271), .A2(n1272), .ZN(n1269) );
NAND2_X1 U918 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
NOR2_X1 U919 ( .A1(n1127), .A2(G952), .ZN(n1181) );
XNOR2_X1 U920 ( .A(G146), .B(n1248), .ZN(G48) );
NAND4_X1 U921 ( .A1(n1115), .A2(n1275), .A3(n1129), .A4(n1107), .ZN(n1248) );
XOR2_X1 U922 ( .A(G143), .B(n1276), .Z(G45) );
NOR4_X1 U923 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(n1276) );
XOR2_X1 U924 ( .A(n1281), .B(KEYINPUT39), .Z(n1280) );
NAND3_X1 U925 ( .A1(n1259), .A2(n1129), .A3(n1098), .ZN(n1277) );
XOR2_X1 U926 ( .A(G140), .B(n1254), .Z(G42) );
AND3_X1 U927 ( .A1(n1264), .A2(n1107), .A3(n1262), .ZN(n1254) );
XOR2_X1 U928 ( .A(G137), .B(n1253), .Z(G39) );
AND4_X1 U929 ( .A1(n1131), .A2(n1275), .A3(n1264), .A4(n1107), .ZN(n1253) );
INV_X1 U930 ( .A(n1094), .ZN(n1264) );
XOR2_X1 U931 ( .A(n1282), .B(n1283), .Z(G36) );
NOR3_X1 U932 ( .A1(n1265), .A2(n1243), .A3(n1094), .ZN(n1283) );
INV_X1 U933 ( .A(n1084), .ZN(n1243) );
NOR2_X1 U934 ( .A1(KEYINPUT29), .A2(n1284), .ZN(n1282) );
XNOR2_X1 U935 ( .A(n1285), .B(n1252), .ZN(G33) );
NOR3_X1 U936 ( .A1(n1265), .A2(n1094), .A3(n1286), .ZN(n1252) );
INV_X1 U937 ( .A(n1115), .ZN(n1286) );
NAND2_X1 U938 ( .A1(n1124), .A2(n1287), .ZN(n1094) );
NAND3_X1 U939 ( .A1(n1107), .A2(n1281), .A3(n1098), .ZN(n1265) );
XNOR2_X1 U940 ( .A(G128), .B(n1255), .ZN(G30) );
NAND4_X1 U941 ( .A1(n1275), .A2(n1084), .A3(n1245), .A4(n1129), .ZN(n1255) );
AND3_X1 U942 ( .A1(n1138), .A2(n1281), .A3(n1288), .ZN(n1275) );
XNOR2_X1 U943 ( .A(n1289), .B(n1238), .ZN(G3) );
AND3_X1 U944 ( .A1(n1098), .A2(n1083), .A3(n1131), .ZN(n1238) );
XNOR2_X1 U945 ( .A(G125), .B(n1290), .ZN(G27) );
NAND3_X1 U946 ( .A1(n1262), .A2(n1291), .A3(n1132), .ZN(n1290) );
XNOR2_X1 U947 ( .A(KEYINPUT36), .B(n1125), .ZN(n1291) );
INV_X1 U948 ( .A(n1129), .ZN(n1125) );
AND3_X1 U949 ( .A1(n1115), .A2(n1281), .A3(n1292), .ZN(n1262) );
NAND2_X1 U950 ( .A1(n1100), .A2(n1293), .ZN(n1281) );
NAND4_X1 U951 ( .A1(G902), .A2(G953), .A3(n1294), .A4(n1155), .ZN(n1293) );
INV_X1 U952 ( .A(G900), .ZN(n1155) );
XOR2_X1 U953 ( .A(G122), .B(n1237), .Z(G24) );
AND4_X1 U954 ( .A1(n1259), .A2(n1295), .A3(n1086), .A4(n1260), .ZN(n1237) );
NOR2_X1 U955 ( .A1(n1138), .A2(n1288), .ZN(n1086) );
XNOR2_X1 U956 ( .A(G119), .B(n1239), .ZN(G21) );
NAND4_X1 U957 ( .A1(n1295), .A2(n1131), .A3(n1288), .A4(n1138), .ZN(n1239) );
XNOR2_X1 U958 ( .A(G116), .B(n1296), .ZN(G18) );
NAND2_X1 U959 ( .A1(n1240), .A2(n1084), .ZN(n1296) );
NOR2_X1 U960 ( .A1(n1259), .A2(n1279), .ZN(n1084) );
INV_X1 U961 ( .A(n1260), .ZN(n1279) );
XNOR2_X1 U962 ( .A(G113), .B(n1297), .ZN(G15) );
NAND2_X1 U963 ( .A1(n1298), .A2(n1240), .ZN(n1297) );
AND2_X1 U964 ( .A1(n1295), .A2(n1098), .ZN(n1240) );
NOR2_X1 U965 ( .A1(n1288), .A2(n1299), .ZN(n1098) );
AND3_X1 U966 ( .A1(n1129), .A2(n1246), .A3(n1132), .ZN(n1295) );
NOR2_X1 U967 ( .A1(n1112), .A2(n1300), .ZN(n1132) );
XNOR2_X1 U968 ( .A(n1115), .B(KEYINPUT16), .ZN(n1298) );
NOR2_X1 U969 ( .A1(n1260), .A2(n1301), .ZN(n1115) );
XNOR2_X1 U970 ( .A(n1302), .B(n1235), .ZN(G12) );
AND3_X1 U971 ( .A1(n1131), .A2(n1083), .A3(n1292), .ZN(n1235) );
INV_X1 U972 ( .A(n1117), .ZN(n1292) );
NAND2_X1 U973 ( .A1(n1299), .A2(n1288), .ZN(n1117) );
XOR2_X1 U974 ( .A(n1141), .B(n1303), .Z(n1288) );
NOR2_X1 U975 ( .A1(KEYINPUT23), .A2(n1142), .ZN(n1303) );
NAND2_X1 U976 ( .A1(G217), .A2(n1304), .ZN(n1142) );
NOR2_X1 U977 ( .A1(n1187), .A2(G902), .ZN(n1141) );
XNOR2_X1 U978 ( .A(n1305), .B(n1306), .ZN(n1187) );
XOR2_X1 U979 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U980 ( .A(n1302), .B(n1309), .ZN(n1308) );
NOR2_X1 U981 ( .A1(KEYINPUT47), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U982 ( .A(G146), .B(n1311), .ZN(n1310) );
NAND2_X1 U983 ( .A1(KEYINPUT40), .A2(n1312), .ZN(n1311) );
AND3_X1 U984 ( .A1(G221), .A2(n1127), .A3(G234), .ZN(n1307) );
XNOR2_X1 U985 ( .A(G119), .B(n1313), .ZN(n1305) );
XNOR2_X1 U986 ( .A(G137), .B(n1314), .ZN(n1313) );
INV_X1 U987 ( .A(G128), .ZN(n1314) );
INV_X1 U988 ( .A(n1138), .ZN(n1299) );
XOR2_X1 U989 ( .A(n1315), .B(n1213), .Z(n1138) );
INV_X1 U990 ( .A(G472), .ZN(n1213) );
NAND2_X1 U991 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U992 ( .A(n1318), .B(n1319), .Z(n1316) );
AND2_X1 U993 ( .A1(n1216), .A2(n1215), .ZN(n1319) );
NAND3_X1 U994 ( .A1(G101), .A2(G210), .A3(n1320), .ZN(n1215) );
NAND2_X1 U995 ( .A1(n1321), .A2(n1289), .ZN(n1216) );
NAND2_X1 U996 ( .A1(n1320), .A2(G210), .ZN(n1321) );
NOR2_X1 U997 ( .A1(KEYINPUT4), .A2(n1322), .ZN(n1318) );
XNOR2_X1 U998 ( .A(n1323), .B(n1324), .ZN(n1322) );
INV_X1 U999 ( .A(n1209), .ZN(n1324) );
XOR2_X1 U1000 ( .A(n1325), .B(n1326), .Z(n1209) );
NOR3_X1 U1001 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1326) );
NOR2_X1 U1002 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NOR2_X1 U1003 ( .A1(n1332), .A2(n1333), .ZN(n1330) );
XNOR2_X1 U1004 ( .A(KEYINPUT18), .B(n1334), .ZN(n1333) );
INV_X1 U1005 ( .A(KEYINPUT8), .ZN(n1332) );
AND3_X1 U1006 ( .A1(n1331), .A2(n1334), .A3(KEYINPUT8), .ZN(n1328) );
XOR2_X1 U1007 ( .A(G116), .B(n1335), .Z(n1331) );
INV_X1 U1008 ( .A(G119), .ZN(n1335) );
NOR2_X1 U1009 ( .A1(KEYINPUT8), .A2(n1334), .ZN(n1327) );
NAND2_X1 U1010 ( .A1(KEYINPUT12), .A2(n1336), .ZN(n1323) );
INV_X1 U1011 ( .A(n1210), .ZN(n1336) );
AND3_X1 U1012 ( .A1(n1245), .A2(n1246), .A3(n1129), .ZN(n1083) );
NOR2_X1 U1013 ( .A1(n1124), .A2(n1123), .ZN(n1129) );
INV_X1 U1014 ( .A(n1287), .ZN(n1123) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1337), .ZN(n1287) );
XOR2_X1 U1016 ( .A(n1338), .B(n1339), .Z(n1124) );
AND2_X1 U1017 ( .A1(n1337), .A2(G210), .ZN(n1339) );
NAND2_X1 U1018 ( .A1(n1340), .A2(n1317), .ZN(n1337) );
XNOR2_X1 U1019 ( .A(G237), .B(KEYINPUT55), .ZN(n1340) );
NAND2_X1 U1020 ( .A1(n1341), .A2(n1317), .ZN(n1338) );
XNOR2_X1 U1021 ( .A(n1270), .B(n1342), .ZN(n1341) );
NAND3_X1 U1022 ( .A1(n1343), .A2(n1344), .A3(n1272), .ZN(n1342) );
OR2_X1 U1023 ( .A1(n1274), .A2(n1273), .ZN(n1272) );
OR2_X1 U1024 ( .A1(n1274), .A2(KEYINPUT17), .ZN(n1344) );
NAND3_X1 U1025 ( .A1(n1273), .A2(n1274), .A3(KEYINPUT17), .ZN(n1343) );
XNOR2_X1 U1026 ( .A(G125), .B(n1345), .ZN(n1274) );
INV_X1 U1027 ( .A(n1325), .ZN(n1345) );
XNOR2_X1 U1028 ( .A(n1346), .B(KEYINPUT32), .ZN(n1325) );
NOR2_X1 U1029 ( .A1(n1176), .A2(G953), .ZN(n1273) );
INV_X1 U1030 ( .A(G224), .ZN(n1176) );
AND3_X1 U1031 ( .A1(n1347), .A2(n1348), .A3(n1178), .ZN(n1270) );
NAND2_X1 U1032 ( .A1(n1349), .A2(n1350), .ZN(n1178) );
NAND2_X1 U1033 ( .A1(KEYINPUT61), .A2(n1351), .ZN(n1348) );
NAND3_X1 U1034 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
INV_X1 U1035 ( .A(n1349), .ZN(n1354) );
NOR2_X1 U1036 ( .A1(n1355), .A2(n1356), .ZN(n1349) );
NAND2_X1 U1037 ( .A1(n1350), .A2(n1357), .ZN(n1353) );
NAND3_X1 U1038 ( .A1(n1358), .A2(n1355), .A3(n1356), .ZN(n1352) );
OR2_X1 U1039 ( .A1(n1179), .A2(KEYINPUT61), .ZN(n1347) );
AND2_X1 U1040 ( .A1(n1359), .A2(n1360), .ZN(n1179) );
NAND2_X1 U1041 ( .A1(n1361), .A2(n1356), .ZN(n1360) );
INV_X1 U1042 ( .A(n1357), .ZN(n1356) );
XNOR2_X1 U1043 ( .A(n1350), .B(n1355), .ZN(n1361) );
INV_X1 U1044 ( .A(n1358), .ZN(n1350) );
NAND3_X1 U1045 ( .A1(n1358), .A2(n1355), .A3(n1357), .ZN(n1359) );
XOR2_X1 U1046 ( .A(G110), .B(n1362), .Z(n1357) );
XOR2_X1 U1047 ( .A(KEYINPUT53), .B(G122), .Z(n1362) );
XNOR2_X1 U1048 ( .A(n1363), .B(n1289), .ZN(n1355) );
NAND3_X1 U1049 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1363) );
NAND2_X1 U1050 ( .A1(KEYINPUT31), .A2(G107), .ZN(n1366) );
NAND3_X1 U1051 ( .A1(n1082), .A2(n1367), .A3(n1368), .ZN(n1365) );
NAND2_X1 U1052 ( .A1(n1369), .A2(n1370), .ZN(n1364) );
NAND2_X1 U1053 ( .A1(n1371), .A2(n1367), .ZN(n1370) );
INV_X1 U1054 ( .A(KEYINPUT31), .ZN(n1367) );
XNOR2_X1 U1055 ( .A(KEYINPUT35), .B(n1082), .ZN(n1371) );
XNOR2_X1 U1056 ( .A(n1372), .B(n1373), .ZN(n1358) );
NOR2_X1 U1057 ( .A1(G113), .A2(KEYINPUT15), .ZN(n1373) );
XNOR2_X1 U1058 ( .A(G119), .B(n1374), .ZN(n1372) );
NOR2_X1 U1059 ( .A1(G116), .A2(KEYINPUT13), .ZN(n1374) );
NAND2_X1 U1060 ( .A1(n1100), .A2(n1375), .ZN(n1246) );
NAND3_X1 U1061 ( .A1(n1180), .A2(n1294), .A3(G902), .ZN(n1375) );
NOR2_X1 U1062 ( .A1(G898), .A2(n1127), .ZN(n1180) );
NAND3_X1 U1063 ( .A1(n1294), .A2(n1127), .A3(G952), .ZN(n1100) );
NAND2_X1 U1064 ( .A1(G234), .A2(G237), .ZN(n1294) );
XNOR2_X1 U1065 ( .A(n1107), .B(KEYINPUT41), .ZN(n1245) );
INV_X1 U1066 ( .A(n1278), .ZN(n1107) );
NAND2_X1 U1067 ( .A1(n1376), .A2(n1112), .ZN(n1278) );
NAND2_X1 U1068 ( .A1(n1135), .A2(n1147), .ZN(n1112) );
NAND3_X1 U1069 ( .A1(n1226), .A2(n1317), .A3(n1377), .ZN(n1147) );
INV_X1 U1070 ( .A(G469), .ZN(n1226) );
NAND2_X1 U1071 ( .A1(G469), .A2(n1378), .ZN(n1135) );
NAND2_X1 U1072 ( .A1(n1377), .A2(n1317), .ZN(n1378) );
XOR2_X1 U1073 ( .A(n1379), .B(n1380), .Z(n1377) );
XOR2_X1 U1074 ( .A(n1381), .B(n1382), .Z(n1380) );
XNOR2_X1 U1075 ( .A(n1383), .B(KEYINPUT54), .ZN(n1382) );
NAND2_X1 U1076 ( .A1(KEYINPUT5), .A2(n1384), .ZN(n1383) );
XNOR2_X1 U1077 ( .A(KEYINPUT56), .B(n1385), .ZN(n1384) );
INV_X1 U1078 ( .A(n1220), .ZN(n1385) );
XNOR2_X1 U1079 ( .A(n1386), .B(n1387), .ZN(n1220) );
XOR2_X1 U1080 ( .A(n1388), .B(n1160), .Z(n1387) );
XOR2_X1 U1081 ( .A(n1346), .B(KEYINPUT62), .Z(n1160) );
XOR2_X1 U1082 ( .A(n1389), .B(G146), .Z(n1346) );
NAND2_X1 U1083 ( .A1(KEYINPUT43), .A2(n1368), .ZN(n1388) );
INV_X1 U1084 ( .A(n1369), .ZN(n1368) );
XOR2_X1 U1085 ( .A(G104), .B(KEYINPUT9), .Z(n1369) );
XNOR2_X1 U1086 ( .A(n1390), .B(n1082), .ZN(n1386) );
NAND2_X1 U1087 ( .A1(KEYINPUT6), .A2(n1289), .ZN(n1390) );
INV_X1 U1088 ( .A(G101), .ZN(n1289) );
NOR2_X1 U1089 ( .A1(KEYINPUT38), .A2(n1224), .ZN(n1381) );
NAND2_X1 U1090 ( .A1(G227), .A2(n1127), .ZN(n1224) );
XNOR2_X1 U1091 ( .A(n1223), .B(n1210), .ZN(n1379) );
XOR2_X1 U1092 ( .A(n1391), .B(n1285), .Z(n1210) );
NAND2_X1 U1093 ( .A1(KEYINPUT10), .A2(n1161), .ZN(n1391) );
XNOR2_X1 U1094 ( .A(n1284), .B(G137), .ZN(n1161) );
XNOR2_X1 U1095 ( .A(G140), .B(n1302), .ZN(n1223) );
XOR2_X1 U1096 ( .A(KEYINPUT34), .B(n1300), .Z(n1376) );
INV_X1 U1097 ( .A(n1111), .ZN(n1300) );
NAND2_X1 U1098 ( .A1(G221), .A2(n1304), .ZN(n1111) );
NAND2_X1 U1099 ( .A1(G234), .A2(n1317), .ZN(n1304) );
NOR2_X1 U1100 ( .A1(n1260), .A2(n1259), .ZN(n1131) );
INV_X1 U1101 ( .A(n1301), .ZN(n1259) );
XNOR2_X1 U1102 ( .A(n1392), .B(n1393), .ZN(n1301) );
NOR2_X1 U1103 ( .A1(KEYINPUT1), .A2(n1394), .ZN(n1393) );
INV_X1 U1104 ( .A(n1143), .ZN(n1394) );
NOR2_X1 U1105 ( .A1(n1202), .A2(G902), .ZN(n1143) );
XNOR2_X1 U1106 ( .A(n1395), .B(n1396), .ZN(n1202) );
XOR2_X1 U1107 ( .A(G104), .B(n1397), .Z(n1396) );
NOR2_X1 U1108 ( .A1(KEYINPUT0), .A2(n1398), .ZN(n1397) );
XNOR2_X1 U1109 ( .A(n1334), .B(n1399), .ZN(n1398) );
XOR2_X1 U1110 ( .A(KEYINPUT30), .B(G122), .Z(n1399) );
INV_X1 U1111 ( .A(G113), .ZN(n1334) );
NAND3_X1 U1112 ( .A1(n1400), .A2(n1401), .A3(KEYINPUT33), .ZN(n1395) );
NAND3_X1 U1113 ( .A1(n1402), .A2(n1403), .A3(n1404), .ZN(n1401) );
INV_X1 U1114 ( .A(KEYINPUT28), .ZN(n1404) );
XNOR2_X1 U1115 ( .A(n1405), .B(n1406), .ZN(n1402) );
NAND2_X1 U1116 ( .A1(n1407), .A2(KEYINPUT28), .ZN(n1400) );
XNOR2_X1 U1117 ( .A(n1408), .B(n1406), .ZN(n1407) );
XNOR2_X1 U1118 ( .A(G146), .B(n1159), .ZN(n1406) );
INV_X1 U1119 ( .A(n1312), .ZN(n1159) );
XOR2_X1 U1120 ( .A(G125), .B(G140), .Z(n1312) );
NAND2_X1 U1121 ( .A1(n1403), .A2(n1405), .ZN(n1408) );
INV_X1 U1122 ( .A(KEYINPUT27), .ZN(n1405) );
XNOR2_X1 U1123 ( .A(n1409), .B(n1285), .ZN(n1403) );
INV_X1 U1124 ( .A(G131), .ZN(n1285) );
NAND2_X1 U1125 ( .A1(KEYINPUT14), .A2(n1410), .ZN(n1409) );
XNOR2_X1 U1126 ( .A(n1411), .B(n1412), .ZN(n1410) );
NAND2_X1 U1127 ( .A1(n1320), .A2(G214), .ZN(n1411) );
NOR2_X1 U1128 ( .A1(G953), .A2(G237), .ZN(n1320) );
XNOR2_X1 U1129 ( .A(G475), .B(KEYINPUT52), .ZN(n1392) );
NAND2_X1 U1130 ( .A1(n1413), .A2(n1145), .ZN(n1260) );
NAND2_X1 U1131 ( .A1(n1414), .A2(n1415), .ZN(n1145) );
NAND2_X1 U1132 ( .A1(n1192), .A2(n1317), .ZN(n1415) );
XNOR2_X1 U1133 ( .A(KEYINPUT24), .B(n1146), .ZN(n1413) );
NAND3_X1 U1134 ( .A1(n1192), .A2(n1317), .A3(n1416), .ZN(n1146) );
INV_X1 U1135 ( .A(n1414), .ZN(n1416) );
XOR2_X1 U1136 ( .A(G478), .B(KEYINPUT37), .Z(n1414) );
INV_X1 U1137 ( .A(G902), .ZN(n1317) );
NAND2_X1 U1138 ( .A1(n1417), .A2(n1418), .ZN(n1192) );
NAND2_X1 U1139 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
INV_X1 U1140 ( .A(n1421), .ZN(n1420) );
XOR2_X1 U1141 ( .A(KEYINPUT45), .B(n1422), .Z(n1419) );
NAND2_X1 U1142 ( .A1(n1423), .A2(n1421), .ZN(n1417) );
XNOR2_X1 U1143 ( .A(n1424), .B(n1425), .ZN(n1421) );
XOR2_X1 U1144 ( .A(G116), .B(n1426), .Z(n1425) );
XNOR2_X1 U1145 ( .A(n1284), .B(G122), .ZN(n1426) );
INV_X1 U1146 ( .A(G134), .ZN(n1284) );
XNOR2_X1 U1147 ( .A(n1389), .B(n1082), .ZN(n1424) );
INV_X1 U1148 ( .A(G107), .ZN(n1082) );
XNOR2_X1 U1149 ( .A(G128), .B(n1412), .ZN(n1389) );
XOR2_X1 U1150 ( .A(G143), .B(KEYINPUT21), .Z(n1412) );
XOR2_X1 U1151 ( .A(KEYINPUT50), .B(n1422), .Z(n1423) );
AND3_X1 U1152 ( .A1(G234), .A2(n1127), .A3(G217), .ZN(n1422) );
INV_X1 U1153 ( .A(G953), .ZN(n1127) );
INV_X1 U1154 ( .A(G110), .ZN(n1302) );
endmodule


