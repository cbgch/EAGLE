//Key = 1010010111110100101001101000101000010001100010101111101010011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381;

XNOR2_X1 U759 ( .A(G107), .B(n1051), .ZN(G9) );
NAND2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(G75) );
NOR4_X1 U762 ( .A1(G953), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U765 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
AND3_X1 U769 ( .A1(KEYINPUT7), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1066) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR3_X1 U772 ( .A1(n1069), .A2(n1078), .A3(n1075), .ZN(n1061) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1081), .A2(n1065), .ZN(n1080) );
INV_X1 U775 ( .A(n1052), .ZN(n1065) );
NOR3_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR2_X1 U777 ( .A1(KEYINPUT7), .A2(n1063), .ZN(n1084) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1063), .ZN(n1079) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR3_X1 U781 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1054) );
AND4_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1056) );
NOR4_X1 U783 ( .A1(n1073), .A2(n1094), .A3(n1063), .A4(n1095), .ZN(n1093) );
XOR2_X1 U784 ( .A(G472), .B(n1096), .Z(n1095) );
NOR2_X1 U785 ( .A1(KEYINPUT19), .A2(n1097), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1098), .B(G475), .Z(n1092) );
XOR2_X1 U787 ( .A(n1099), .B(G478), .Z(n1091) );
XOR2_X1 U788 ( .A(n1100), .B(n1101), .Z(n1090) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(G72) );
XOR2_X1 U790 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U792 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XOR2_X1 U793 ( .A(n1109), .B(KEYINPUT26), .Z(n1106) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U797 ( .A1(KEYINPUT39), .A2(n1116), .ZN(n1115) );
INV_X1 U798 ( .A(n1117), .ZN(n1116) );
INV_X1 U799 ( .A(KEYINPUT63), .ZN(n1114) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1110) );
NAND2_X1 U801 ( .A1(KEYINPUT39), .A2(n1119), .ZN(n1118) );
OR2_X1 U802 ( .A1(n1112), .A2(KEYINPUT63), .ZN(n1119) );
XNOR2_X1 U803 ( .A(n1120), .B(KEYINPUT27), .ZN(n1112) );
XNOR2_X1 U804 ( .A(n1121), .B(n1122), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1123), .B(KEYINPUT59), .Z(n1121) );
NAND2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U807 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U808 ( .A(KEYINPUT44), .B(n1128), .Z(n1124) );
NOR2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1128) );
NAND2_X1 U810 ( .A1(n1129), .A2(n1130), .ZN(n1104) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U812 ( .A(KEYINPUT40), .B(n1133), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1134), .A2(n1129), .ZN(n1102) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1108), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(G69) );
NAND2_X1 U816 ( .A1(n1138), .A2(n1129), .ZN(n1137) );
XNOR2_X1 U817 ( .A(n1139), .B(n1140), .ZN(n1138) );
NAND2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
XNOR2_X1 U819 ( .A(n1143), .B(KEYINPUT49), .ZN(n1141) );
NAND2_X1 U820 ( .A1(n1144), .A2(G953), .ZN(n1136) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1140), .A2(n1147), .ZN(n1146) );
NAND2_X1 U823 ( .A1(G224), .A2(n1148), .ZN(n1145) );
NAND2_X1 U824 ( .A1(G898), .A2(n1140), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1149), .A2(n1150), .ZN(n1140) );
NAND2_X1 U826 ( .A1(G953), .A2(n1151), .ZN(n1150) );
XOR2_X1 U827 ( .A(n1152), .B(n1153), .Z(n1149) );
NAND2_X1 U828 ( .A1(KEYINPUT8), .A2(n1154), .ZN(n1152) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XNOR2_X1 U830 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1161), .ZN(G63) );
XNOR2_X1 U833 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1160), .ZN(n1162) );
INV_X1 U835 ( .A(G478), .ZN(n1164) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1165), .ZN(G60) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U839 ( .A1(n1170), .A2(n1160), .ZN(n1169) );
AND2_X1 U840 ( .A1(n1171), .A2(KEYINPUT18), .ZN(n1168) );
NOR2_X1 U841 ( .A1(KEYINPUT18), .A2(n1171), .ZN(n1166) );
XNOR2_X1 U842 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U843 ( .A1(n1173), .A2(KEYINPUT57), .ZN(n1172) );
INV_X1 U844 ( .A(n1174), .ZN(n1173) );
NOR3_X1 U845 ( .A1(n1155), .A2(n1175), .A3(n1176), .ZN(G57) );
NOR2_X1 U846 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U847 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U848 ( .A1(KEYINPUT6), .A2(n1181), .ZN(n1180) );
NOR2_X1 U849 ( .A1(G101), .A2(n1182), .ZN(n1175) );
XOR2_X1 U850 ( .A(n1179), .B(n1183), .Z(n1182) );
NOR2_X1 U851 ( .A1(n1184), .A2(KEYINPUT6), .ZN(n1183) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1179) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1185) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1160), .ZN(n1188) );
INV_X1 U855 ( .A(G472), .ZN(n1189) );
NAND2_X1 U856 ( .A1(KEYINPUT2), .A2(n1190), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1155), .A2(n1191), .ZN(G54) );
XOR2_X1 U858 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U859 ( .A1(n1100), .A2(n1160), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NAND4_X1 U861 ( .A1(KEYINPUT54), .A2(KEYINPUT22), .A3(n1196), .A4(n1197), .ZN(n1195) );
NAND2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1194) );
NAND2_X1 U863 ( .A1(n1197), .A2(n1200), .ZN(n1199) );
OR2_X1 U864 ( .A1(n1196), .A2(KEYINPUT54), .ZN(n1200) );
XOR2_X1 U865 ( .A(n1201), .B(n1202), .Z(n1197) );
XOR2_X1 U866 ( .A(KEYINPUT4), .B(n1203), .Z(n1202) );
NAND2_X1 U867 ( .A1(KEYINPUT22), .A2(n1196), .ZN(n1198) );
XNOR2_X1 U868 ( .A(n1204), .B(n1122), .ZN(n1196) );
XOR2_X1 U869 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U870 ( .A1(KEYINPUT12), .A2(n1207), .ZN(n1206) );
NOR2_X1 U871 ( .A1(n1208), .A2(n1209), .ZN(G51) );
XOR2_X1 U872 ( .A(KEYINPUT3), .B(n1155), .Z(n1209) );
NOR2_X1 U873 ( .A1(n1129), .A2(G952), .ZN(n1155) );
XOR2_X1 U874 ( .A(n1210), .B(n1211), .Z(n1208) );
XOR2_X1 U875 ( .A(n1212), .B(n1213), .Z(n1210) );
NOR2_X1 U876 ( .A1(n1214), .A2(n1160), .ZN(n1213) );
NAND2_X1 U877 ( .A1(G902), .A2(n1058), .ZN(n1160) );
NAND4_X1 U878 ( .A1(n1143), .A2(n1131), .A3(n1142), .A4(n1133), .ZN(n1058) );
NAND2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1133) );
AND4_X1 U880 ( .A1(n1217), .A2(n1174), .A3(n1218), .A4(n1219), .ZN(n1142) );
NAND3_X1 U881 ( .A1(n1052), .A2(n1220), .A3(n1077), .ZN(n1174) );
NAND2_X1 U882 ( .A1(n1053), .A2(n1221), .ZN(n1217) );
XOR2_X1 U883 ( .A(KEYINPUT42), .B(n1052), .Z(n1221) );
AND2_X1 U884 ( .A1(n1220), .A2(n1076), .ZN(n1053) );
AND4_X1 U885 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1131) );
NOR4_X1 U886 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NAND3_X1 U887 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1222) );
XOR2_X1 U888 ( .A(KEYINPUT15), .B(n1071), .Z(n1230) );
AND4_X1 U889 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1143) );
NAND2_X1 U890 ( .A1(n1237), .A2(n1083), .ZN(n1233) );
XOR2_X1 U891 ( .A(n1238), .B(KEYINPUT51), .Z(n1237) );
NAND3_X1 U892 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1212) );
INV_X1 U893 ( .A(n1242), .ZN(n1241) );
NAND3_X1 U894 ( .A1(G125), .A2(n1190), .A3(n1243), .ZN(n1240) );
OR2_X1 U895 ( .A1(n1243), .A2(G125), .ZN(n1239) );
INV_X1 U896 ( .A(KEYINPUT20), .ZN(n1243) );
XOR2_X1 U897 ( .A(G146), .B(n1229), .Z(G48) );
AND2_X1 U898 ( .A1(n1244), .A2(n1077), .ZN(n1229) );
XNOR2_X1 U899 ( .A(n1228), .B(n1245), .ZN(G45) );
XOR2_X1 U900 ( .A(n1246), .B(KEYINPUT31), .Z(n1245) );
AND4_X1 U901 ( .A1(n1247), .A2(n1089), .A3(n1248), .A4(n1249), .ZN(n1228) );
NOR2_X1 U902 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
XOR2_X1 U903 ( .A(n1252), .B(n1253), .Z(G42) );
NOR2_X1 U904 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U905 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND4_X1 U906 ( .A1(n1247), .A2(n1088), .A3(n1077), .A4(n1063), .ZN(n1257) );
INV_X1 U907 ( .A(KEYINPUT55), .ZN(n1256) );
NOR2_X1 U908 ( .A1(KEYINPUT55), .A2(n1224), .ZN(n1254) );
NAND3_X1 U909 ( .A1(n1088), .A2(n1077), .A3(n1215), .ZN(n1224) );
XOR2_X1 U910 ( .A(n1258), .B(n1259), .Z(G39) );
NAND2_X1 U911 ( .A1(KEYINPUT28), .A2(G137), .ZN(n1259) );
NAND4_X1 U912 ( .A1(n1260), .A2(n1216), .A3(n1261), .A4(n1071), .ZN(n1258) );
XOR2_X1 U913 ( .A(n1231), .B(KEYINPUT33), .Z(n1260) );
XNOR2_X1 U914 ( .A(G134), .B(n1223), .ZN(G36) );
NAND3_X1 U915 ( .A1(n1089), .A2(n1076), .A3(n1215), .ZN(n1223) );
NOR2_X1 U916 ( .A1(n1262), .A2(n1063), .ZN(n1215) );
INV_X1 U917 ( .A(n1261), .ZN(n1063) );
NAND2_X1 U918 ( .A1(n1263), .A2(n1264), .ZN(G33) );
NAND2_X1 U919 ( .A1(G131), .A2(n1265), .ZN(n1264) );
NAND2_X1 U920 ( .A1(n1232), .A2(n1247), .ZN(n1265) );
INV_X1 U921 ( .A(n1266), .ZN(n1232) );
XOR2_X1 U922 ( .A(KEYINPUT60), .B(n1267), .Z(n1263) );
NOR3_X1 U923 ( .A1(n1266), .A2(G131), .A3(n1262), .ZN(n1267) );
NAND3_X1 U924 ( .A1(n1089), .A2(n1261), .A3(n1077), .ZN(n1266) );
NOR2_X1 U925 ( .A1(n1086), .A2(n1268), .ZN(n1261) );
XOR2_X1 U926 ( .A(G128), .B(n1227), .Z(G30) );
AND2_X1 U927 ( .A1(n1244), .A2(n1076), .ZN(n1227) );
AND4_X1 U928 ( .A1(n1247), .A2(n1083), .A3(n1269), .A4(n1094), .ZN(n1244) );
INV_X1 U929 ( .A(n1262), .ZN(n1247) );
NAND2_X1 U930 ( .A1(n1071), .A2(n1231), .ZN(n1262) );
XOR2_X1 U931 ( .A(n1177), .B(n1218), .Z(G3) );
NAND3_X1 U932 ( .A1(n1089), .A2(n1220), .A3(n1270), .ZN(n1218) );
XOR2_X1 U933 ( .A(G125), .B(n1226), .Z(G27) );
AND4_X1 U934 ( .A1(n1088), .A2(n1077), .A3(n1271), .A4(n1272), .ZN(n1226) );
AND2_X1 U935 ( .A1(n1231), .A2(n1083), .ZN(n1271) );
NAND2_X1 U936 ( .A1(n1060), .A2(n1273), .ZN(n1231) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1274), .A4(n1108), .ZN(n1273) );
INV_X1 U938 ( .A(G900), .ZN(n1108) );
XOR2_X1 U939 ( .A(G122), .B(n1275), .Z(G24) );
NOR2_X1 U940 ( .A1(n1250), .A2(n1238), .ZN(n1275) );
NAND4_X1 U941 ( .A1(n1276), .A2(n1277), .A3(n1052), .A4(n1278), .ZN(n1238) );
NOR2_X1 U942 ( .A1(n1075), .A2(n1279), .ZN(n1278) );
NOR2_X1 U943 ( .A1(n1094), .A2(n1269), .ZN(n1052) );
XOR2_X1 U944 ( .A(n1280), .B(n1234), .Z(G21) );
NAND2_X1 U945 ( .A1(n1216), .A2(n1281), .ZN(n1234) );
AND3_X1 U946 ( .A1(n1269), .A2(n1094), .A3(n1270), .ZN(n1216) );
INV_X1 U947 ( .A(n1282), .ZN(n1094) );
XNOR2_X1 U948 ( .A(G116), .B(n1235), .ZN(G18) );
NAND3_X1 U949 ( .A1(n1281), .A2(n1076), .A3(n1089), .ZN(n1235) );
NOR2_X1 U950 ( .A1(n1251), .A2(n1249), .ZN(n1076) );
XNOR2_X1 U951 ( .A(G113), .B(n1236), .ZN(G15) );
NAND3_X1 U952 ( .A1(n1089), .A2(n1281), .A3(n1077), .ZN(n1236) );
NOR2_X1 U953 ( .A1(n1279), .A2(n1276), .ZN(n1077) );
AND3_X1 U954 ( .A1(n1083), .A2(n1277), .A3(n1272), .ZN(n1281) );
INV_X1 U955 ( .A(n1075), .ZN(n1272) );
NAND2_X1 U956 ( .A1(n1072), .A2(n1283), .ZN(n1075) );
AND2_X1 U957 ( .A1(n1282), .A2(n1269), .ZN(n1089) );
XNOR2_X1 U958 ( .A(G110), .B(n1219), .ZN(G12) );
NAND3_X1 U959 ( .A1(n1270), .A2(n1220), .A3(n1088), .ZN(n1219) );
NOR2_X1 U960 ( .A1(n1269), .A2(n1282), .ZN(n1088) );
XNOR2_X1 U961 ( .A(n1284), .B(n1159), .ZN(n1282) );
NAND2_X1 U962 ( .A1(G217), .A2(n1285), .ZN(n1159) );
NAND2_X1 U963 ( .A1(n1158), .A2(n1286), .ZN(n1284) );
XOR2_X1 U964 ( .A(n1287), .B(n1288), .Z(n1158) );
XOR2_X1 U965 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U966 ( .A(n1291), .B(n1292), .Z(n1290) );
NOR2_X1 U967 ( .A1(KEYINPUT14), .A2(G125), .ZN(n1292) );
NAND2_X1 U968 ( .A1(G221), .A2(n1293), .ZN(n1291) );
XOR2_X1 U969 ( .A(n1294), .B(n1295), .Z(n1287) );
NOR2_X1 U970 ( .A1(KEYINPUT45), .A2(n1296), .ZN(n1295) );
XOR2_X1 U971 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U972 ( .A(G110), .B(G128), .ZN(n1298) );
NAND2_X1 U973 ( .A1(KEYINPUT24), .A2(n1280), .ZN(n1297) );
INV_X1 U974 ( .A(G119), .ZN(n1280) );
XOR2_X1 U975 ( .A(G137), .B(n1252), .Z(n1294) );
XNOR2_X1 U976 ( .A(n1097), .B(G472), .ZN(n1269) );
NAND2_X1 U977 ( .A1(n1299), .A2(n1286), .ZN(n1097) );
XOR2_X1 U978 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U979 ( .A(n1302), .B(n1184), .Z(n1301) );
INV_X1 U980 ( .A(n1181), .ZN(n1184) );
NAND3_X1 U981 ( .A1(n1303), .A2(n1129), .A3(G210), .ZN(n1181) );
NOR2_X1 U982 ( .A1(G101), .A2(KEYINPUT47), .ZN(n1302) );
XNOR2_X1 U983 ( .A(n1186), .B(n1190), .ZN(n1300) );
XNOR2_X1 U984 ( .A(n1304), .B(n1305), .ZN(n1186) );
XOR2_X1 U985 ( .A(G119), .B(n1306), .Z(n1305) );
NOR2_X1 U986 ( .A1(G113), .A2(KEYINPUT38), .ZN(n1306) );
XOR2_X1 U987 ( .A(n1307), .B(n1308), .Z(n1304) );
NOR2_X1 U988 ( .A1(G116), .A2(KEYINPUT17), .ZN(n1308) );
AND3_X1 U989 ( .A1(n1083), .A2(n1277), .A3(n1071), .ZN(n1220) );
NOR2_X1 U990 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U991 ( .A(n1283), .ZN(n1073) );
NAND2_X1 U992 ( .A1(n1309), .A2(n1285), .ZN(n1283) );
NAND2_X1 U993 ( .A1(G234), .A2(n1310), .ZN(n1285) );
XOR2_X1 U994 ( .A(KEYINPUT41), .B(G221), .Z(n1309) );
XNOR2_X1 U995 ( .A(n1311), .B(n1101), .ZN(n1072) );
AND2_X1 U996 ( .A1(n1286), .A2(n1312), .ZN(n1101) );
XOR2_X1 U997 ( .A(n1313), .B(n1314), .Z(n1312) );
NAND2_X1 U998 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U999 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1000 ( .A1(KEYINPUT35), .A2(n1319), .ZN(n1318) );
OR2_X1 U1001 ( .A1(n1207), .A2(KEYINPUT1), .ZN(n1319) );
NAND2_X1 U1002 ( .A1(n1207), .A2(n1320), .ZN(n1315) );
NAND2_X1 U1003 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1004 ( .A1(KEYINPUT35), .A2(n1323), .ZN(n1322) );
INV_X1 U1005 ( .A(n1317), .ZN(n1323) );
XOR2_X1 U1006 ( .A(n1205), .B(n1324), .Z(n1317) );
NOR2_X1 U1007 ( .A1(KEYINPUT32), .A2(n1122), .ZN(n1324) );
XOR2_X1 U1008 ( .A(n1289), .B(n1325), .Z(n1122) );
XOR2_X1 U1009 ( .A(G128), .B(n1326), .Z(n1325) );
NOR2_X1 U1010 ( .A1(KEYINPUT53), .A2(n1246), .ZN(n1326) );
INV_X1 U1011 ( .A(G143), .ZN(n1246) );
XOR2_X1 U1012 ( .A(n1177), .B(n1327), .Z(n1205) );
INV_X1 U1013 ( .A(KEYINPUT1), .ZN(n1321) );
XOR2_X1 U1014 ( .A(n1307), .B(KEYINPUT16), .Z(n1207) );
XNOR2_X1 U1015 ( .A(n1328), .B(n1126), .ZN(n1307) );
XNOR2_X1 U1016 ( .A(G134), .B(G137), .ZN(n1126) );
NAND2_X1 U1017 ( .A1(KEYINPUT30), .A2(n1127), .ZN(n1328) );
INV_X1 U1018 ( .A(G131), .ZN(n1127) );
NAND2_X1 U1019 ( .A1(n1329), .A2(n1330), .ZN(n1313) );
NAND2_X1 U1020 ( .A1(n1331), .A2(n1201), .ZN(n1330) );
XOR2_X1 U1021 ( .A(KEYINPUT9), .B(n1332), .Z(n1329) );
NOR2_X1 U1022 ( .A1(n1331), .A2(n1201), .ZN(n1332) );
XOR2_X1 U1023 ( .A(G110), .B(n1333), .Z(n1201) );
XOR2_X1 U1024 ( .A(KEYINPUT5), .B(G140), .Z(n1333) );
XNOR2_X1 U1025 ( .A(KEYINPUT61), .B(n1203), .ZN(n1331) );
NOR2_X1 U1026 ( .A1(n1135), .A2(G953), .ZN(n1203) );
INV_X1 U1027 ( .A(G227), .ZN(n1135) );
NAND2_X1 U1028 ( .A1(KEYINPUT0), .A2(n1100), .ZN(n1311) );
INV_X1 U1029 ( .A(G469), .ZN(n1100) );
NAND2_X1 U1030 ( .A1(n1060), .A2(n1334), .ZN(n1277) );
NAND4_X1 U1031 ( .A1(G953), .A2(G902), .A3(n1274), .A4(n1151), .ZN(n1334) );
INV_X1 U1032 ( .A(G898), .ZN(n1151) );
NAND3_X1 U1033 ( .A1(n1274), .A2(n1129), .A3(G952), .ZN(n1060) );
NAND2_X1 U1034 ( .A1(G237), .A2(G234), .ZN(n1274) );
INV_X1 U1035 ( .A(n1250), .ZN(n1083) );
NAND2_X1 U1036 ( .A1(n1335), .A2(n1086), .ZN(n1250) );
XOR2_X1 U1037 ( .A(n1336), .B(n1214), .Z(n1086) );
NAND2_X1 U1038 ( .A1(G210), .A2(n1337), .ZN(n1214) );
NAND2_X1 U1039 ( .A1(n1286), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1040 ( .A(n1339), .B(n1211), .Z(n1338) );
XNOR2_X1 U1041 ( .A(n1154), .B(n1340), .ZN(n1211) );
XOR2_X1 U1042 ( .A(n1341), .B(n1153), .Z(n1340) );
XNOR2_X1 U1043 ( .A(n1342), .B(n1343), .ZN(n1153) );
XOR2_X1 U1044 ( .A(G113), .B(n1344), .Z(n1343) );
NOR2_X1 U1045 ( .A1(KEYINPUT43), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1046 ( .A(G116), .B(n1346), .Z(n1345) );
XOR2_X1 U1047 ( .A(KEYINPUT56), .B(G119), .Z(n1346) );
NAND3_X1 U1048 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1342) );
OR2_X1 U1049 ( .A1(n1350), .A2(G101), .ZN(n1349) );
NAND2_X1 U1050 ( .A1(n1351), .A2(n1352), .ZN(n1348) );
INV_X1 U1051 ( .A(KEYINPUT21), .ZN(n1352) );
NAND2_X1 U1052 ( .A1(n1353), .A2(n1350), .ZN(n1351) );
XOR2_X1 U1053 ( .A(KEYINPUT13), .B(n1177), .Z(n1353) );
INV_X1 U1054 ( .A(G101), .ZN(n1177) );
NAND2_X1 U1055 ( .A1(KEYINPUT21), .A2(n1354), .ZN(n1347) );
NAND2_X1 U1056 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
OR2_X1 U1057 ( .A1(G101), .A2(KEYINPUT13), .ZN(n1356) );
NAND3_X1 U1058 ( .A1(G101), .A2(n1350), .A3(KEYINPUT13), .ZN(n1355) );
XNOR2_X1 U1059 ( .A(n1327), .B(KEYINPUT10), .ZN(n1350) );
XOR2_X1 U1060 ( .A(G104), .B(G107), .Z(n1327) );
NOR2_X1 U1061 ( .A1(G953), .A2(n1147), .ZN(n1341) );
INV_X1 U1062 ( .A(G224), .ZN(n1147) );
XNOR2_X1 U1063 ( .A(G110), .B(n1357), .ZN(n1154) );
XOR2_X1 U1064 ( .A(KEYINPUT46), .B(G122), .Z(n1357) );
NOR2_X1 U1065 ( .A1(n1242), .A2(n1358), .ZN(n1339) );
XOR2_X1 U1066 ( .A(n1359), .B(KEYINPUT48), .Z(n1358) );
NAND2_X1 U1067 ( .A1(G125), .A2(n1190), .ZN(n1359) );
NOR2_X1 U1068 ( .A1(n1190), .A2(G125), .ZN(n1242) );
XNOR2_X1 U1069 ( .A(n1360), .B(n1361), .ZN(n1190) );
XOR2_X1 U1070 ( .A(G143), .B(G128), .Z(n1361) );
NAND2_X1 U1071 ( .A1(KEYINPUT11), .A2(n1289), .ZN(n1360) );
XNOR2_X1 U1072 ( .A(n1268), .B(KEYINPUT58), .ZN(n1335) );
INV_X1 U1073 ( .A(n1085), .ZN(n1268) );
NAND2_X1 U1074 ( .A1(G214), .A2(n1337), .ZN(n1085) );
NAND2_X1 U1075 ( .A1(n1310), .A2(n1303), .ZN(n1337) );
INV_X1 U1076 ( .A(n1069), .ZN(n1270) );
NAND2_X1 U1077 ( .A1(n1279), .A2(n1251), .ZN(n1069) );
INV_X1 U1078 ( .A(n1276), .ZN(n1251) );
XOR2_X1 U1079 ( .A(n1099), .B(n1362), .Z(n1276) );
NOR2_X1 U1080 ( .A1(G478), .A2(KEYINPUT23), .ZN(n1362) );
NAND2_X1 U1081 ( .A1(n1163), .A2(n1286), .ZN(n1099) );
XOR2_X1 U1082 ( .A(n1363), .B(n1364), .Z(n1163) );
XOR2_X1 U1083 ( .A(n1365), .B(n1366), .Z(n1364) );
XOR2_X1 U1084 ( .A(G134), .B(G128), .Z(n1366) );
XOR2_X1 U1085 ( .A(KEYINPUT29), .B(G143), .Z(n1365) );
XOR2_X1 U1086 ( .A(n1367), .B(n1368), .Z(n1363) );
XOR2_X1 U1087 ( .A(G116), .B(G107), .Z(n1368) );
XOR2_X1 U1088 ( .A(n1369), .B(n1370), .Z(n1367) );
NOR2_X1 U1089 ( .A1(KEYINPUT36), .A2(G122), .ZN(n1370) );
NAND2_X1 U1090 ( .A1(n1293), .A2(G217), .ZN(n1369) );
AND2_X1 U1091 ( .A1(G234), .A2(n1129), .ZN(n1293) );
INV_X1 U1092 ( .A(n1249), .ZN(n1279) );
XNOR2_X1 U1093 ( .A(n1371), .B(n1098), .ZN(n1249) );
NAND2_X1 U1094 ( .A1(n1286), .A2(n1171), .ZN(n1098) );
XNOR2_X1 U1095 ( .A(n1372), .B(KEYINPUT25), .ZN(n1171) );
XOR2_X1 U1096 ( .A(n1373), .B(n1374), .Z(n1372) );
XOR2_X1 U1097 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1098 ( .A(G122), .B(G104), .Z(n1376) );
XOR2_X1 U1099 ( .A(G143), .B(G131), .Z(n1375) );
XOR2_X1 U1100 ( .A(n1377), .B(n1378), .Z(n1373) );
XOR2_X1 U1101 ( .A(n1379), .B(n1120), .Z(n1378) );
XNOR2_X1 U1102 ( .A(n1252), .B(G125), .ZN(n1120) );
INV_X1 U1103 ( .A(G140), .ZN(n1252) );
NOR2_X1 U1104 ( .A1(G113), .A2(KEYINPUT37), .ZN(n1379) );
XOR2_X1 U1105 ( .A(n1380), .B(n1381), .Z(n1377) );
AND3_X1 U1106 ( .A1(G214), .A2(n1129), .A3(n1303), .ZN(n1381) );
INV_X1 U1107 ( .A(G237), .ZN(n1303) );
INV_X1 U1108 ( .A(G953), .ZN(n1129) );
NAND2_X1 U1109 ( .A1(KEYINPUT50), .A2(n1289), .ZN(n1380) );
XNOR2_X1 U1110 ( .A(G146), .B(KEYINPUT34), .ZN(n1289) );
XOR2_X1 U1111 ( .A(n1310), .B(KEYINPUT62), .Z(n1286) );
INV_X1 U1112 ( .A(G902), .ZN(n1310) );
NAND2_X1 U1113 ( .A1(KEYINPUT52), .A2(n1170), .ZN(n1371) );
INV_X1 U1114 ( .A(G475), .ZN(n1170) );
endmodule


