//Key = 0001111010010101110111110111001000001101010110000010101000001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XNOR2_X1 U723 ( .A(n1005), .B(n1006), .ZN(G9) );
NAND3_X1 U724 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(G75) );
NAND2_X1 U725 ( .A1(G952), .A2(n1010), .ZN(n1009) );
NAND2_X1 U726 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U727 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U728 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND4_X1 U729 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NAND2_X1 U730 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NAND2_X1 U731 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U732 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1021) );
XNOR2_X1 U734 ( .A(n1029), .B(n1030), .ZN(n1028) );
NAND3_X1 U735 ( .A1(n1023), .A2(n1031), .A3(n1027), .ZN(n1015) );
NAND2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U737 ( .A1(n1034), .A2(n1035), .A3(n1017), .ZN(n1033) );
NAND2_X1 U738 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U739 ( .A1(n1038), .A2(n1039), .A3(n1020), .ZN(n1034) );
NAND2_X1 U740 ( .A1(n1040), .A2(n1018), .ZN(n1032) );
NAND4_X1 U741 ( .A1(n1023), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1007) );
NOR4_X1 U742 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U743 ( .A(KEYINPUT32), .B(n1048), .Z(n1047) );
XNOR2_X1 U744 ( .A(n1049), .B(n1050), .ZN(n1046) );
XOR2_X1 U745 ( .A(n1051), .B(n1052), .Z(n1045) );
NAND2_X1 U746 ( .A1(n1053), .A2(KEYINPUT62), .ZN(n1052) );
XOR2_X1 U747 ( .A(n1054), .B(KEYINPUT11), .Z(n1053) );
XNOR2_X1 U748 ( .A(n1055), .B(n1056), .ZN(n1044) );
NOR2_X1 U749 ( .A1(KEYINPUT51), .A2(n1057), .ZN(n1056) );
NOR2_X1 U750 ( .A1(n1036), .A2(n1058), .ZN(n1042) );
XNOR2_X1 U751 ( .A(n1059), .B(n1060), .ZN(n1041) );
XOR2_X1 U752 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n1060) );
XOR2_X1 U753 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U754 ( .A1(n1063), .A2(n1008), .ZN(n1062) );
AND2_X1 U755 ( .A1(G227), .A2(G900), .ZN(n1063) );
NAND2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NAND2_X1 U757 ( .A1(n1066), .A2(n1008), .ZN(n1065) );
XOR2_X1 U758 ( .A(n1067), .B(n1068), .Z(n1066) );
NAND3_X1 U759 ( .A1(G900), .A2(n1068), .A3(G953), .ZN(n1064) );
XOR2_X1 U760 ( .A(n1069), .B(n1070), .Z(n1068) );
XOR2_X1 U761 ( .A(n1071), .B(n1072), .Z(n1069) );
NAND2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U764 ( .A(KEYINPUT42), .B(G134), .Z(n1076) );
XNOR2_X1 U765 ( .A(KEYINPUT17), .B(G137), .ZN(n1075) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
XOR2_X1 U767 ( .A(KEYINPUT21), .B(G134), .Z(n1078) );
XOR2_X1 U768 ( .A(KEYINPUT17), .B(G137), .Z(n1077) );
XOR2_X1 U769 ( .A(n1079), .B(n1080), .Z(G69) );
NOR2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U771 ( .A(n1083), .ZN(n1082) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND2_X1 U773 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NAND2_X1 U774 ( .A1(G898), .A2(G224), .ZN(n1086) );
INV_X1 U775 ( .A(n1087), .ZN(n1084) );
NOR2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1050), .ZN(n1090) );
INV_X1 U779 ( .A(n1094), .ZN(n1050) );
INV_X1 U780 ( .A(n1011), .ZN(n1093) );
XNOR2_X1 U781 ( .A(KEYINPUT0), .B(n1095), .ZN(n1092) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1096), .ZN(G63) );
XNOR2_X1 U783 ( .A(n1097), .B(n1098), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1099), .B(KEYINPUT15), .Z(n1098) );
NAND2_X1 U785 ( .A1(n1100), .A2(G478), .ZN(n1099) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1101), .ZN(G60) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U788 ( .A1(n1100), .A2(G475), .ZN(n1102) );
XOR2_X1 U789 ( .A(G104), .B(n1104), .Z(G6) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(G57) );
XOR2_X1 U791 ( .A(KEYINPUT14), .B(n1088), .Z(n1106) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(n1105) );
XNOR2_X1 U793 ( .A(G101), .B(n1109), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1110), .A2(KEYINPUT6), .ZN(n1107) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1111) );
NOR3_X1 U798 ( .A1(n1117), .A2(KEYINPUT35), .A3(n1057), .ZN(n1116) );
INV_X1 U799 ( .A(G472), .ZN(n1057) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XNOR2_X1 U802 ( .A(KEYINPUT40), .B(n1122), .ZN(n1121) );
XNOR2_X1 U803 ( .A(n1123), .B(KEYINPUT30), .ZN(n1120) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
XNOR2_X1 U805 ( .A(KEYINPUT43), .B(n1126), .ZN(n1125) );
XNOR2_X1 U806 ( .A(KEYINPUT40), .B(n1127), .ZN(n1124) );
NOR3_X1 U807 ( .A1(n1088), .A2(n1128), .A3(n1129), .ZN(G54) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1130) );
NOR2_X1 U810 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
INV_X1 U811 ( .A(KEYINPUT37), .ZN(n1135) );
NOR2_X1 U812 ( .A1(n1136), .A2(n1137), .ZN(n1128) );
XOR2_X1 U813 ( .A(n1132), .B(n1138), .Z(n1137) );
AND2_X1 U814 ( .A1(KEYINPUT37), .A2(n1134), .ZN(n1138) );
XOR2_X1 U815 ( .A(n1139), .B(n1126), .Z(n1134) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
INV_X1 U818 ( .A(KEYINPUT58), .ZN(n1143) );
NAND3_X1 U819 ( .A1(n1144), .A2(n1122), .A3(KEYINPUT58), .ZN(n1140) );
AND2_X1 U820 ( .A1(n1100), .A2(G469), .ZN(n1132) );
INV_X1 U821 ( .A(n1131), .ZN(n1136) );
NAND2_X1 U822 ( .A1(n1145), .A2(KEYINPUT44), .ZN(n1131) );
XNOR2_X1 U823 ( .A(n1146), .B(G110), .ZN(n1145) );
NOR2_X1 U824 ( .A1(n1088), .A2(n1147), .ZN(G51) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U826 ( .A(n1150), .B(n1083), .ZN(n1149) );
OR2_X1 U827 ( .A1(n1117), .A2(n1054), .ZN(n1150) );
INV_X1 U828 ( .A(n1100), .ZN(n1117) );
NOR2_X1 U829 ( .A1(n1095), .A2(n1011), .ZN(n1100) );
NOR2_X1 U830 ( .A1(n1067), .A2(n1087), .ZN(n1011) );
NAND4_X1 U831 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1087) );
NOR4_X1 U832 ( .A1(n1104), .A2(n1006), .A3(n1155), .A4(n1156), .ZN(n1154) );
NOR3_X1 U833 ( .A1(n1026), .A2(n1037), .A3(n1157), .ZN(n1006) );
INV_X1 U834 ( .A(n1158), .ZN(n1026) );
NOR3_X1 U835 ( .A1(n1157), .A2(n1037), .A3(n1025), .ZN(n1104) );
INV_X1 U836 ( .A(n1018), .ZN(n1037) );
NOR2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
INV_X1 U838 ( .A(n1161), .ZN(n1159) );
OR3_X1 U839 ( .A1(n1162), .A2(n1157), .A3(n1038), .ZN(n1151) );
NAND4_X1 U840 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1067) );
NOR4_X1 U841 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U842 ( .A(n1171), .ZN(n1168) );
NOR3_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1165) );
AND2_X1 U844 ( .A1(KEYINPUT8), .A2(n1175), .ZN(n1174) );
NOR3_X1 U845 ( .A1(KEYINPUT8), .A2(n1176), .A3(n1177), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1025), .A2(n1178), .ZN(n1172) );
XNOR2_X1 U847 ( .A(n1179), .B(KEYINPUT1), .ZN(n1148) );
NAND2_X1 U848 ( .A1(KEYINPUT63), .A2(n1180), .ZN(n1179) );
XOR2_X1 U849 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND3_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
NAND2_X1 U851 ( .A1(KEYINPUT12), .A2(n1186), .ZN(n1185) );
NAND3_X1 U852 ( .A1(n1187), .A2(n1188), .A3(n1122), .ZN(n1184) );
INV_X1 U853 ( .A(KEYINPUT12), .ZN(n1188) );
OR2_X1 U854 ( .A1(n1122), .A2(n1187), .ZN(n1183) );
NOR2_X1 U855 ( .A1(KEYINPUT45), .A2(n1186), .ZN(n1187) );
NOR2_X1 U856 ( .A1(n1008), .A2(G952), .ZN(n1088) );
XNOR2_X1 U857 ( .A(G146), .B(n1164), .ZN(G48) );
NAND2_X1 U858 ( .A1(n1189), .A2(n1190), .ZN(n1164) );
XNOR2_X1 U859 ( .A(n1191), .B(n1175), .ZN(G45) );
NOR2_X1 U860 ( .A1(n1177), .A2(n1038), .ZN(n1175) );
NAND4_X1 U861 ( .A1(n1192), .A2(n1040), .A3(n1193), .A4(n1194), .ZN(n1177) );
XOR2_X1 U862 ( .A(G140), .B(n1170), .Z(G42) );
AND3_X1 U863 ( .A1(n1190), .A2(n1195), .A3(n1196), .ZN(n1170) );
XOR2_X1 U864 ( .A(n1197), .B(n1169), .Z(G39) );
AND3_X1 U865 ( .A1(n1196), .A2(n1198), .A3(n1027), .ZN(n1169) );
NAND2_X1 U866 ( .A1(n1199), .A2(KEYINPUT13), .ZN(n1197) );
XNOR2_X1 U867 ( .A(G137), .B(KEYINPUT2), .ZN(n1199) );
XOR2_X1 U868 ( .A(n1200), .B(G134), .Z(G36) );
NAND2_X1 U869 ( .A1(KEYINPUT41), .A2(n1163), .ZN(n1200) );
NAND2_X1 U870 ( .A1(n1201), .A2(n1158), .ZN(n1163) );
XOR2_X1 U871 ( .A(n1202), .B(n1203), .Z(G33) );
XOR2_X1 U872 ( .A(KEYINPUT52), .B(G131), .Z(n1203) );
NAND2_X1 U873 ( .A1(n1201), .A2(n1204), .ZN(n1202) );
XNOR2_X1 U874 ( .A(KEYINPUT7), .B(n1025), .ZN(n1204) );
INV_X1 U875 ( .A(n1190), .ZN(n1025) );
INV_X1 U876 ( .A(n1178), .ZN(n1201) );
NAND2_X1 U877 ( .A1(n1176), .A2(n1196), .ZN(n1178) );
AND3_X1 U878 ( .A1(n1192), .A2(n1020), .A3(n1017), .ZN(n1196) );
XNOR2_X1 U879 ( .A(n1205), .B(n1206), .ZN(G30) );
NOR2_X1 U880 ( .A1(KEYINPUT38), .A2(n1171), .ZN(n1206) );
NAND2_X1 U881 ( .A1(n1189), .A2(n1158), .ZN(n1171) );
AND3_X1 U882 ( .A1(n1198), .A2(n1040), .A3(n1192), .ZN(n1189) );
AND3_X1 U883 ( .A1(n1207), .A2(n1029), .A3(n1030), .ZN(n1192) );
XOR2_X1 U884 ( .A(n1208), .B(n1209), .Z(G3) );
XNOR2_X1 U885 ( .A(KEYINPUT59), .B(n1210), .ZN(n1209) );
NOR4_X1 U886 ( .A1(KEYINPUT49), .A2(n1157), .A3(n1162), .A4(n1038), .ZN(n1208) );
XOR2_X1 U887 ( .A(n1211), .B(n1212), .Z(G27) );
XNOR2_X1 U888 ( .A(G125), .B(KEYINPUT16), .ZN(n1212) );
NAND2_X1 U889 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NAND2_X1 U890 ( .A1(n1167), .A2(n1215), .ZN(n1214) );
INV_X1 U891 ( .A(KEYINPUT10), .ZN(n1215) );
NOR2_X1 U892 ( .A1(n1216), .A2(n1217), .ZN(n1167) );
INV_X1 U893 ( .A(n1040), .ZN(n1217) );
NAND3_X1 U894 ( .A1(n1040), .A2(n1216), .A3(KEYINPUT10), .ZN(n1213) );
NAND4_X1 U895 ( .A1(n1190), .A2(n1023), .A3(n1195), .A4(n1207), .ZN(n1216) );
NAND2_X1 U896 ( .A1(n1218), .A2(n1219), .ZN(n1207) );
NAND4_X1 U897 ( .A1(G902), .A2(G953), .A3(n1014), .A4(n1220), .ZN(n1219) );
INV_X1 U898 ( .A(G900), .ZN(n1220) );
XNOR2_X1 U899 ( .A(G122), .B(n1152), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1221), .A2(n1018), .A3(n1193), .A4(n1194), .ZN(n1152) );
NAND2_X1 U901 ( .A1(n1222), .A2(n1223), .ZN(n1018) );
OR3_X1 U902 ( .A1(n1224), .A2(n1225), .A3(KEYINPUT34), .ZN(n1223) );
NAND2_X1 U903 ( .A1(KEYINPUT34), .A2(n1195), .ZN(n1222) );
XOR2_X1 U904 ( .A(G119), .B(n1160), .Z(G21) );
AND3_X1 U905 ( .A1(n1027), .A2(n1198), .A3(n1221), .ZN(n1160) );
AND2_X1 U906 ( .A1(n1224), .A2(n1225), .ZN(n1198) );
XNOR2_X1 U907 ( .A(G116), .B(n1161), .ZN(G18) );
NAND3_X1 U908 ( .A1(n1176), .A2(n1158), .A3(n1221), .ZN(n1161) );
NOR2_X1 U909 ( .A1(n1193), .A2(n1226), .ZN(n1158) );
XOR2_X1 U910 ( .A(G113), .B(n1156), .Z(G15) );
AND3_X1 U911 ( .A1(n1176), .A2(n1190), .A3(n1221), .ZN(n1156) );
AND2_X1 U912 ( .A1(n1023), .A2(n1227), .ZN(n1221) );
NOR2_X1 U913 ( .A1(n1030), .A2(n1228), .ZN(n1023) );
INV_X1 U914 ( .A(n1029), .ZN(n1228) );
NOR2_X1 U915 ( .A1(n1194), .A2(n1059), .ZN(n1190) );
INV_X1 U916 ( .A(n1193), .ZN(n1059) );
INV_X1 U917 ( .A(n1038), .ZN(n1176) );
NAND2_X1 U918 ( .A1(n1229), .A2(n1225), .ZN(n1038) );
XNOR2_X1 U919 ( .A(KEYINPUT34), .B(n1224), .ZN(n1229) );
INV_X1 U920 ( .A(n1230), .ZN(n1224) );
XNOR2_X1 U921 ( .A(n1231), .B(n1155), .ZN(G12) );
NOR3_X1 U922 ( .A1(n1157), .A2(n1039), .A3(n1162), .ZN(n1155) );
INV_X1 U923 ( .A(n1027), .ZN(n1162) );
NOR2_X1 U924 ( .A1(n1194), .A2(n1193), .ZN(n1027) );
XNOR2_X1 U925 ( .A(n1232), .B(G475), .ZN(n1193) );
NAND2_X1 U926 ( .A1(n1103), .A2(n1095), .ZN(n1232) );
XOR2_X1 U927 ( .A(n1233), .B(G113), .Z(n1103) );
XOR2_X1 U928 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U929 ( .A(n1236), .B(n1070), .Z(n1235) );
XOR2_X1 U930 ( .A(G140), .B(G131), .Z(n1070) );
XOR2_X1 U931 ( .A(KEYINPUT28), .B(G146), .Z(n1236) );
XOR2_X1 U932 ( .A(n1237), .B(n1238), .Z(n1234) );
XOR2_X1 U933 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U934 ( .A1(KEYINPUT25), .A2(n1241), .ZN(n1240) );
NAND2_X1 U935 ( .A1(n1242), .A2(n1243), .ZN(n1239) );
NAND2_X1 U936 ( .A1(n1244), .A2(n1191), .ZN(n1243) );
XOR2_X1 U937 ( .A(KEYINPUT50), .B(n1245), .Z(n1242) );
NOR2_X1 U938 ( .A1(n1191), .A2(n1244), .ZN(n1245) );
NAND3_X1 U939 ( .A1(n1246), .A2(n1247), .A3(G214), .ZN(n1244) );
XNOR2_X1 U940 ( .A(G104), .B(G122), .ZN(n1237) );
INV_X1 U941 ( .A(n1226), .ZN(n1194) );
NOR2_X1 U942 ( .A1(n1048), .A2(n1058), .ZN(n1226) );
AND2_X1 U943 ( .A1(n1248), .A2(G478), .ZN(n1058) );
NOR2_X1 U944 ( .A1(n1248), .A2(G478), .ZN(n1048) );
NAND2_X1 U945 ( .A1(n1097), .A2(n1095), .ZN(n1248) );
XNOR2_X1 U946 ( .A(n1249), .B(n1250), .ZN(n1097) );
XOR2_X1 U947 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U948 ( .A(G107), .B(n1253), .ZN(n1252) );
NOR2_X1 U949 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U950 ( .A(G217), .ZN(n1255) );
NAND2_X1 U951 ( .A1(KEYINPUT4), .A2(G143), .ZN(n1251) );
XOR2_X1 U952 ( .A(n1256), .B(n1257), .Z(n1249) );
XNOR2_X1 U953 ( .A(G134), .B(n1205), .ZN(n1257) );
XNOR2_X1 U954 ( .A(G116), .B(G122), .ZN(n1256) );
INV_X1 U955 ( .A(n1195), .ZN(n1039) );
NOR2_X1 U956 ( .A1(n1225), .A2(n1230), .ZN(n1195) );
XOR2_X1 U957 ( .A(n1258), .B(n1094), .Z(n1230) );
NAND2_X1 U958 ( .A1(G217), .A2(n1259), .ZN(n1094) );
NAND2_X1 U959 ( .A1(n1260), .A2(KEYINPUT54), .ZN(n1258) );
XOR2_X1 U960 ( .A(n1049), .B(KEYINPUT33), .Z(n1260) );
NAND2_X1 U961 ( .A1(n1091), .A2(n1095), .ZN(n1049) );
XOR2_X1 U962 ( .A(n1261), .B(n1262), .Z(n1091) );
NOR2_X1 U963 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U964 ( .A(n1265), .B(KEYINPUT19), .Z(n1264) );
NAND2_X1 U965 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NOR2_X1 U966 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
NAND2_X1 U967 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U968 ( .A1(G146), .A2(n1270), .ZN(n1269) );
XOR2_X1 U969 ( .A(KEYINPUT5), .B(n1271), .Z(n1268) );
NOR2_X1 U970 ( .A1(G146), .A2(n1270), .ZN(n1271) );
XNOR2_X1 U971 ( .A(G140), .B(n1241), .ZN(n1270) );
XNOR2_X1 U972 ( .A(n1231), .B(n1272), .ZN(n1266) );
XNOR2_X1 U973 ( .A(n1205), .B(G119), .ZN(n1272) );
INV_X1 U974 ( .A(G128), .ZN(n1205) );
XNOR2_X1 U975 ( .A(G137), .B(n1273), .ZN(n1261) );
NOR2_X1 U976 ( .A1(n1274), .A2(n1254), .ZN(n1273) );
NAND2_X1 U977 ( .A1(n1275), .A2(n1246), .ZN(n1254) );
XNOR2_X1 U978 ( .A(G234), .B(KEYINPUT27), .ZN(n1275) );
INV_X1 U979 ( .A(G221), .ZN(n1274) );
XNOR2_X1 U980 ( .A(n1055), .B(G472), .ZN(n1225) );
NAND2_X1 U981 ( .A1(n1276), .A2(n1095), .ZN(n1055) );
XOR2_X1 U982 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U983 ( .A(n1279), .B(n1114), .Z(n1278) );
XNOR2_X1 U984 ( .A(G119), .B(KEYINPUT22), .ZN(n1114) );
XNOR2_X1 U985 ( .A(n1280), .B(n1109), .ZN(n1277) );
NAND3_X1 U986 ( .A1(n1246), .A2(n1247), .A3(G210), .ZN(n1109) );
NAND3_X1 U987 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1280) );
NAND2_X1 U988 ( .A1(KEYINPUT48), .A2(n1126), .ZN(n1283) );
NAND3_X1 U989 ( .A1(n1123), .A2(n1284), .A3(n1127), .ZN(n1282) );
NAND2_X1 U990 ( .A1(n1122), .A2(n1285), .ZN(n1281) );
NAND2_X1 U991 ( .A1(n1286), .A2(n1284), .ZN(n1285) );
INV_X1 U992 ( .A(KEYINPUT48), .ZN(n1284) );
XNOR2_X1 U993 ( .A(KEYINPUT46), .B(n1126), .ZN(n1286) );
INV_X1 U994 ( .A(n1127), .ZN(n1122) );
NAND3_X1 U995 ( .A1(n1030), .A2(n1029), .A3(n1227), .ZN(n1157) );
AND2_X1 U996 ( .A1(n1040), .A2(n1287), .ZN(n1227) );
NAND2_X1 U997 ( .A1(n1218), .A2(n1288), .ZN(n1287) );
NAND3_X1 U998 ( .A1(n1081), .A2(n1014), .A3(G902), .ZN(n1288) );
NOR2_X1 U999 ( .A1(n1008), .A2(G898), .ZN(n1081) );
NAND3_X1 U1000 ( .A1(n1289), .A2(n1008), .A3(G952), .ZN(n1218) );
XNOR2_X1 U1001 ( .A(KEYINPUT39), .B(n1014), .ZN(n1289) );
NAND2_X1 U1002 ( .A1(G237), .A2(G234), .ZN(n1014) );
NOR2_X1 U1003 ( .A1(n1017), .A2(n1036), .ZN(n1040) );
INV_X1 U1004 ( .A(n1020), .ZN(n1036) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1290), .ZN(n1020) );
XNOR2_X1 U1006 ( .A(n1051), .B(n1054), .ZN(n1017) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1290), .ZN(n1054) );
NAND2_X1 U1008 ( .A1(n1247), .A2(n1095), .ZN(n1290) );
INV_X1 U1009 ( .A(G237), .ZN(n1247) );
NAND2_X1 U1010 ( .A1(n1291), .A2(n1095), .ZN(n1051) );
XOR2_X1 U1011 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U1012 ( .A(n1294), .B(n1295), .ZN(n1293) );
NOR2_X1 U1013 ( .A1(KEYINPUT9), .A2(n1083), .ZN(n1295) );
XNOR2_X1 U1014 ( .A(n1296), .B(n1297), .ZN(n1083) );
XOR2_X1 U1015 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U1016 ( .A(n1300), .B(G110), .ZN(n1299) );
INV_X1 U1017 ( .A(G122), .ZN(n1300) );
XOR2_X1 U1018 ( .A(KEYINPUT53), .B(KEYINPUT3), .Z(n1298) );
XOR2_X1 U1019 ( .A(n1279), .B(n1301), .Z(n1296) );
XOR2_X1 U1020 ( .A(n1302), .B(n1303), .Z(n1301) );
NOR2_X1 U1021 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1022 ( .A(n1306), .B(KEYINPUT36), .Z(n1305) );
NOR2_X1 U1023 ( .A1(KEYINPUT56), .A2(n1307), .ZN(n1302) );
XOR2_X1 U1024 ( .A(KEYINPUT18), .B(G119), .Z(n1307) );
XNOR2_X1 U1025 ( .A(n1113), .B(n1210), .ZN(n1279) );
INV_X1 U1026 ( .A(G101), .ZN(n1210) );
XOR2_X1 U1027 ( .A(n1308), .B(n1309), .Z(n1113) );
XNOR2_X1 U1028 ( .A(n1310), .B(G113), .ZN(n1309) );
INV_X1 U1029 ( .A(G116), .ZN(n1310) );
XNOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT31), .ZN(n1308) );
NAND2_X1 U1031 ( .A1(KEYINPUT60), .A2(n1072), .ZN(n1294) );
XNOR2_X1 U1032 ( .A(n1241), .B(n1127), .ZN(n1072) );
INV_X1 U1033 ( .A(n1186), .ZN(n1241) );
XOR2_X1 U1034 ( .A(G125), .B(KEYINPUT47), .Z(n1186) );
XNOR2_X1 U1035 ( .A(KEYINPUT29), .B(n1181), .ZN(n1292) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1246), .ZN(n1181) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1259), .ZN(n1029) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1095), .ZN(n1259) );
XNOR2_X1 U1039 ( .A(n1311), .B(G469), .ZN(n1030) );
NAND2_X1 U1040 ( .A1(n1312), .A2(n1095), .ZN(n1311) );
INV_X1 U1041 ( .A(G902), .ZN(n1095) );
XOR2_X1 U1042 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1043 ( .A(n1142), .B(n1126), .ZN(n1314) );
INV_X1 U1044 ( .A(n1123), .ZN(n1126) );
XNOR2_X1 U1045 ( .A(n1315), .B(n1316), .ZN(n1123) );
XOR2_X1 U1046 ( .A(G137), .B(G131), .Z(n1316) );
NAND2_X1 U1047 ( .A1(KEYINPUT20), .A2(G134), .ZN(n1315) );
XNOR2_X1 U1048 ( .A(n1127), .B(n1144), .ZN(n1142) );
XNOR2_X1 U1049 ( .A(n1317), .B(G101), .ZN(n1144) );
NAND2_X1 U1050 ( .A1(n1318), .A2(n1306), .ZN(n1317) );
NAND2_X1 U1051 ( .A1(G104), .A2(n1005), .ZN(n1306) );
XNOR2_X1 U1052 ( .A(n1304), .B(KEYINPUT57), .ZN(n1318) );
NOR2_X1 U1053 ( .A1(n1005), .A2(G104), .ZN(n1304) );
INV_X1 U1054 ( .A(G107), .ZN(n1005) );
XOR2_X1 U1055 ( .A(G128), .B(n1319), .Z(n1127) );
XNOR2_X1 U1056 ( .A(G146), .B(n1191), .ZN(n1319) );
INV_X1 U1057 ( .A(G143), .ZN(n1191) );
NAND2_X1 U1058 ( .A1(n1320), .A2(n1321), .ZN(n1313) );
NAND2_X1 U1059 ( .A1(G110), .A2(n1322), .ZN(n1321) );
NAND2_X1 U1060 ( .A1(n1323), .A2(n1231), .ZN(n1320) );
XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(n1322), .ZN(n1323) );
INV_X1 U1062 ( .A(n1146), .ZN(n1322) );
XNOR2_X1 U1063 ( .A(n1324), .B(G140), .ZN(n1146) );
NAND2_X1 U1064 ( .A1(G227), .A2(n1246), .ZN(n1324) );
XNOR2_X1 U1065 ( .A(n1008), .B(KEYINPUT26), .ZN(n1246) );
INV_X1 U1066 ( .A(G953), .ZN(n1008) );
INV_X1 U1067 ( .A(G110), .ZN(n1231) );
endmodule


