//Key = 0000100110100000000010100000111101000111111100000000100110001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414;

XOR2_X1 U776 ( .A(G107), .B(n1081), .Z(G9) );
NOR2_X1 U777 ( .A1(n1082), .A2(n1083), .ZN(G75) );
NOR4_X1 U778 ( .A1(G953), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1083) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR3_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NOR2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(n1098) );
NOR2_X1 U789 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR3_X1 U791 ( .A1(n1101), .A2(n1112), .A3(n1113), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
AND2_X1 U793 ( .A1(n1096), .A2(KEYINPUT17), .ZN(n1115) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1107), .ZN(n1112) );
NOR2_X1 U795 ( .A1(KEYINPUT17), .A2(n1117), .ZN(n1116) );
NOR4_X1 U796 ( .A1(n1118), .A2(n1119), .A3(n1096), .A4(n1101), .ZN(n1089) );
NOR2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U798 ( .A1(n1122), .A2(n1091), .ZN(n1120) );
XNOR2_X1 U799 ( .A(n1114), .B(KEYINPUT36), .ZN(n1122) );
NOR2_X1 U800 ( .A1(n1123), .A2(n1093), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1117), .A2(n1107), .ZN(n1123) );
NOR3_X1 U802 ( .A1(n1124), .A2(n1125), .A3(n1096), .ZN(n1117) );
NOR3_X1 U803 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1082) );
AND4_X1 U804 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1084) );
NOR3_X1 U805 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
XOR2_X1 U806 ( .A(n1133), .B(KEYINPUT43), .Z(n1131) );
NAND2_X1 U807 ( .A1(G472), .A2(n1134), .ZN(n1133) );
NAND3_X1 U808 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1130) );
XNOR2_X1 U809 ( .A(n1138), .B(KEYINPUT9), .ZN(n1137) );
NAND2_X1 U810 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
INV_X1 U811 ( .A(G478), .ZN(n1140) );
NAND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
OR2_X1 U814 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
INV_X1 U815 ( .A(KEYINPUT41), .ZN(n1144) );
NAND2_X1 U816 ( .A1(n1145), .A2(G478), .ZN(n1135) );
NOR2_X1 U817 ( .A1(n1146), .A2(KEYINPUT0), .ZN(n1145) );
INV_X1 U818 ( .A(n1143), .ZN(n1146) );
NOR3_X1 U819 ( .A1(n1096), .A2(n1147), .A3(n1148), .ZN(n1128) );
INV_X1 U820 ( .A(n1149), .ZN(n1096) );
XNOR2_X1 U821 ( .A(KEYINPUT57), .B(n1104), .ZN(n1127) );
XOR2_X1 U822 ( .A(n1150), .B(n1151), .Z(n1126) );
XNOR2_X1 U823 ( .A(KEYINPUT2), .B(n1152), .ZN(n1151) );
NOR2_X1 U824 ( .A1(G469), .A2(KEYINPUT44), .ZN(n1150) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(G72) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U827 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U828 ( .A(n1159), .B(n1160), .Z(n1158) );
XNOR2_X1 U829 ( .A(n1161), .B(n1162), .ZN(n1160) );
XNOR2_X1 U830 ( .A(G134), .B(n1163), .ZN(n1159) );
NAND2_X1 U831 ( .A1(KEYINPUT56), .A2(n1164), .ZN(n1163) );
NOR2_X1 U832 ( .A1(G900), .A2(n1165), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1155) );
NAND3_X1 U834 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
XOR2_X1 U835 ( .A(n1171), .B(KEYINPUT47), .Z(n1170) );
XNOR2_X1 U836 ( .A(G953), .B(KEYINPUT18), .ZN(n1166) );
NAND2_X1 U837 ( .A1(G953), .A2(n1172), .ZN(n1153) );
NAND2_X1 U838 ( .A1(G900), .A2(G227), .ZN(n1172) );
XOR2_X1 U839 ( .A(n1173), .B(n1174), .Z(G69) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U841 ( .A1(n1177), .A2(KEYINPUT54), .A3(G953), .ZN(n1176) );
NOR2_X1 U842 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
XNOR2_X1 U843 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U844 ( .A1(KEYINPUT35), .A2(n1182), .ZN(n1181) );
NOR2_X1 U845 ( .A1(G898), .A2(n1165), .ZN(n1178) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1165), .ZN(n1173) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1187), .ZN(G66) );
NOR2_X1 U849 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U850 ( .A(n1190), .B(KEYINPUT55), .Z(n1189) );
NAND2_X1 U851 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
NAND4_X1 U853 ( .A1(G217), .A2(n1086), .A3(n1193), .A4(n1194), .ZN(n1192) );
NAND2_X1 U854 ( .A1(G902), .A2(n1195), .ZN(n1194) );
NAND2_X1 U855 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
NAND2_X1 U856 ( .A1(n1195), .A2(n1198), .ZN(n1196) );
INV_X1 U857 ( .A(KEYINPUT4), .ZN(n1195) );
NOR3_X1 U858 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(G63) );
NOR3_X1 U859 ( .A1(n1202), .A2(G953), .A3(G952), .ZN(n1201) );
AND2_X1 U860 ( .A1(n1202), .A2(n1186), .ZN(n1200) );
INV_X1 U861 ( .A(KEYINPUT59), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
XOR2_X1 U863 ( .A(KEYINPUT51), .B(n1205), .Z(n1204) );
NOR2_X1 U864 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
AND2_X1 U865 ( .A1(n1207), .A2(n1206), .ZN(n1203) );
XNOR2_X1 U866 ( .A(n1208), .B(KEYINPUT62), .ZN(n1206) );
NAND2_X1 U867 ( .A1(n1209), .A2(G478), .ZN(n1207) );
NOR2_X1 U868 ( .A1(n1186), .A2(n1210), .ZN(G60) );
XOR2_X1 U869 ( .A(n1211), .B(n1212), .Z(n1210) );
NOR2_X1 U870 ( .A1(n1213), .A2(KEYINPUT50), .ZN(n1211) );
AND2_X1 U871 ( .A1(G475), .A2(n1209), .ZN(n1213) );
XNOR2_X1 U872 ( .A(G104), .B(n1214), .ZN(G6) );
NOR2_X1 U873 ( .A1(n1186), .A2(n1215), .ZN(G57) );
XOR2_X1 U874 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U877 ( .A1(n1222), .A2(n1223), .ZN(n1218) );
XOR2_X1 U878 ( .A(KEYINPUT34), .B(n1224), .Z(n1223) );
NAND2_X1 U879 ( .A1(n1225), .A2(n1226), .ZN(n1216) );
NAND2_X1 U880 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XNOR2_X1 U881 ( .A(KEYINPUT39), .B(n1229), .ZN(n1227) );
OR2_X1 U882 ( .A1(n1229), .A2(n1228), .ZN(n1225) );
NOR2_X1 U883 ( .A1(n1186), .A2(n1230), .ZN(G54) );
XOR2_X1 U884 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U885 ( .A(n1233), .B(n1234), .Z(n1232) );
AND2_X1 U886 ( .A1(G469), .A2(n1209), .ZN(n1234) );
XOR2_X1 U887 ( .A(n1235), .B(n1236), .Z(n1231) );
NOR2_X1 U888 ( .A1(KEYINPUT13), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U889 ( .A(G140), .B(G110), .ZN(n1237) );
NAND2_X1 U890 ( .A1(n1238), .A2(n1239), .ZN(n1235) );
NAND2_X1 U891 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
XOR2_X1 U892 ( .A(n1242), .B(KEYINPUT16), .Z(n1240) );
NOR2_X1 U893 ( .A1(n1186), .A2(n1243), .ZN(G51) );
XOR2_X1 U894 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND3_X1 U895 ( .A1(n1209), .A2(G210), .A3(KEYINPUT20), .ZN(n1244) );
INV_X1 U896 ( .A(n1221), .ZN(n1209) );
NAND2_X1 U897 ( .A1(G902), .A2(n1086), .ZN(n1221) );
NAND3_X1 U898 ( .A1(n1168), .A2(n1246), .A3(n1177), .ZN(n1086) );
AND4_X1 U899 ( .A1(n1247), .A2(n1214), .A3(n1248), .A4(n1249), .ZN(n1177) );
NOR4_X1 U900 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1081), .ZN(n1249) );
AND3_X1 U901 ( .A1(n1124), .A2(n1253), .A3(n1254), .ZN(n1081) );
INV_X1 U902 ( .A(n1255), .ZN(n1250) );
NOR2_X1 U903 ( .A1(n1256), .A2(n1257), .ZN(n1248) );
NOR2_X1 U904 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NOR2_X1 U905 ( .A1(n1260), .A2(n1261), .ZN(n1256) );
XNOR2_X1 U906 ( .A(n1109), .B(KEYINPUT46), .ZN(n1260) );
NAND3_X1 U907 ( .A1(n1254), .A2(n1253), .A3(n1125), .ZN(n1214) );
NAND3_X1 U908 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1247) );
NOR3_X1 U909 ( .A1(n1101), .A2(n1265), .A3(n1266), .ZN(n1264) );
INV_X1 U910 ( .A(n1253), .ZN(n1101) );
XNOR2_X1 U911 ( .A(n1103), .B(KEYINPUT60), .ZN(n1262) );
XOR2_X1 U912 ( .A(KEYINPUT5), .B(n1267), .Z(n1246) );
AND2_X1 U913 ( .A1(n1171), .A2(n1169), .ZN(n1267) );
AND3_X1 U914 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1169) );
NAND2_X1 U915 ( .A1(n1271), .A2(n1103), .ZN(n1270) );
XNOR2_X1 U916 ( .A(KEYINPUT25), .B(n1272), .ZN(n1271) );
NAND3_X1 U917 ( .A1(n1273), .A2(n1274), .A3(n1114), .ZN(n1268) );
AND4_X1 U918 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1168) );
NAND4_X1 U919 ( .A1(n1279), .A2(n1125), .A3(n1109), .A4(n1280), .ZN(n1275) );
XNOR2_X1 U920 ( .A(KEYINPUT32), .B(n1107), .ZN(n1280) );
INV_X1 U921 ( .A(n1114), .ZN(n1107) );
NOR2_X1 U922 ( .A1(n1165), .A2(G952), .ZN(n1186) );
NAND2_X1 U923 ( .A1(n1281), .A2(n1282), .ZN(G48) );
NAND2_X1 U924 ( .A1(G146), .A2(n1283), .ZN(n1282) );
XOR2_X1 U925 ( .A(n1284), .B(n1285), .Z(n1281) );
NOR2_X1 U926 ( .A1(n1286), .A2(n1272), .ZN(n1285) );
NAND2_X1 U927 ( .A1(n1273), .A2(n1125), .ZN(n1272) );
NOR2_X1 U928 ( .A1(G146), .A2(n1283), .ZN(n1284) );
INV_X1 U929 ( .A(KEYINPUT61), .ZN(n1283) );
XNOR2_X1 U930 ( .A(G143), .B(n1171), .ZN(G45) );
NAND3_X1 U931 ( .A1(n1279), .A2(n1109), .A3(n1287), .ZN(n1171) );
XNOR2_X1 U932 ( .A(G140), .B(n1269), .ZN(G42) );
NAND2_X1 U933 ( .A1(n1288), .A2(n1289), .ZN(n1269) );
XNOR2_X1 U934 ( .A(G137), .B(n1290), .ZN(G39) );
NAND4_X1 U935 ( .A1(KEYINPUT33), .A2(n1114), .A3(n1273), .A4(n1274), .ZN(n1290) );
XNOR2_X1 U936 ( .A(G134), .B(n1276), .ZN(G36) );
NAND3_X1 U937 ( .A1(n1109), .A2(n1124), .A3(n1288), .ZN(n1276) );
INV_X1 U938 ( .A(n1291), .ZN(n1288) );
XNOR2_X1 U939 ( .A(n1292), .B(n1293), .ZN(G33) );
NOR3_X1 U940 ( .A1(n1294), .A2(n1295), .A3(n1291), .ZN(n1293) );
NAND2_X1 U941 ( .A1(n1114), .A2(n1279), .ZN(n1291) );
NOR2_X1 U942 ( .A1(n1104), .A2(n1148), .ZN(n1114) );
INV_X1 U943 ( .A(n1105), .ZN(n1148) );
XNOR2_X1 U944 ( .A(KEYINPUT40), .B(n1258), .ZN(n1294) );
XNOR2_X1 U945 ( .A(G128), .B(n1277), .ZN(G30) );
NAND3_X1 U946 ( .A1(n1124), .A2(n1103), .A3(n1273), .ZN(n1277) );
AND3_X1 U947 ( .A1(n1132), .A2(n1111), .A3(n1279), .ZN(n1273) );
AND3_X1 U948 ( .A1(n1296), .A2(n1149), .A3(n1093), .ZN(n1279) );
XOR2_X1 U949 ( .A(G101), .B(n1252), .Z(G3) );
AND3_X1 U950 ( .A1(n1274), .A2(n1254), .A3(n1109), .ZN(n1252) );
XNOR2_X1 U951 ( .A(G125), .B(n1278), .ZN(G27) );
NAND4_X1 U952 ( .A1(n1296), .A2(n1149), .A3(n1121), .A4(n1297), .ZN(n1278) );
AND2_X1 U953 ( .A1(n1103), .A2(n1289), .ZN(n1297) );
NOR3_X1 U954 ( .A1(n1111), .A2(n1110), .A3(n1295), .ZN(n1289) );
NAND2_X1 U955 ( .A1(n1088), .A2(n1298), .ZN(n1296) );
NAND2_X1 U956 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U957 ( .A(G900), .ZN(n1300) );
XOR2_X1 U958 ( .A(n1301), .B(n1302), .Z(G24) );
NOR2_X1 U959 ( .A1(KEYINPUT12), .A2(n1303), .ZN(n1302) );
AND3_X1 U960 ( .A1(n1287), .A2(n1253), .A3(n1263), .ZN(n1301) );
NOR2_X1 U961 ( .A1(n1111), .A2(n1132), .ZN(n1253) );
NOR3_X1 U962 ( .A1(n1266), .A2(n1265), .A3(n1286), .ZN(n1287) );
XOR2_X1 U963 ( .A(n1251), .B(n1304), .Z(G21) );
NOR2_X1 U964 ( .A1(KEYINPUT27), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U965 ( .A(G119), .B(KEYINPUT49), .ZN(n1305) );
AND3_X1 U966 ( .A1(n1263), .A2(n1274), .A3(n1306), .ZN(n1251) );
NOR3_X1 U967 ( .A1(n1286), .A2(n1307), .A3(n1110), .ZN(n1306) );
INV_X1 U968 ( .A(n1132), .ZN(n1110) );
INV_X1 U969 ( .A(n1103), .ZN(n1286) );
XNOR2_X1 U970 ( .A(G116), .B(n1308), .ZN(G18) );
NAND3_X1 U971 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1308) );
XNOR2_X1 U972 ( .A(n1109), .B(KEYINPUT29), .ZN(n1311) );
XOR2_X1 U973 ( .A(KEYINPUT6), .B(KEYINPUT30), .Z(n1310) );
INV_X1 U974 ( .A(n1259), .ZN(n1309) );
NAND3_X1 U975 ( .A1(n1124), .A2(n1103), .A3(n1263), .ZN(n1259) );
XOR2_X1 U976 ( .A(n1312), .B(KEYINPUT58), .Z(n1103) );
NOR2_X1 U977 ( .A1(n1138), .A2(n1265), .ZN(n1124) );
XNOR2_X1 U978 ( .A(G113), .B(n1313), .ZN(G15) );
OR2_X1 U979 ( .A1(n1261), .A2(n1258), .ZN(n1313) );
INV_X1 U980 ( .A(n1109), .ZN(n1258) );
NOR2_X1 U981 ( .A1(n1132), .A2(n1307), .ZN(n1109) );
NAND3_X1 U982 ( .A1(n1263), .A2(n1312), .A3(n1125), .ZN(n1261) );
INV_X1 U983 ( .A(n1295), .ZN(n1125) );
NAND2_X1 U984 ( .A1(n1265), .A2(n1138), .ZN(n1295) );
AND3_X1 U985 ( .A1(n1314), .A2(n1149), .A3(n1121), .ZN(n1263) );
XNOR2_X1 U986 ( .A(G110), .B(n1255), .ZN(G12) );
NAND4_X1 U987 ( .A1(n1274), .A2(n1254), .A3(n1307), .A4(n1132), .ZN(n1255) );
NAND3_X1 U988 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1132) );
OR2_X1 U989 ( .A1(n1318), .A2(n1191), .ZN(n1317) );
NAND3_X1 U990 ( .A1(n1191), .A2(n1318), .A3(n1197), .ZN(n1316) );
NAND2_X1 U991 ( .A1(G217), .A2(n1198), .ZN(n1318) );
INV_X1 U992 ( .A(G234), .ZN(n1198) );
XOR2_X1 U993 ( .A(n1319), .B(n1320), .Z(n1191) );
XOR2_X1 U994 ( .A(n1321), .B(n1322), .Z(n1320) );
NAND2_X1 U995 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND2_X1 U996 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XNOR2_X1 U997 ( .A(KEYINPUT26), .B(n1327), .ZN(n1326) );
XNOR2_X1 U998 ( .A(G119), .B(G128), .ZN(n1325) );
NAND2_X1 U999 ( .A1(n1328), .A2(n1329), .ZN(n1323) );
XNOR2_X1 U1000 ( .A(KEYINPUT31), .B(n1327), .ZN(n1329) );
XOR2_X1 U1001 ( .A(G128), .B(G119), .Z(n1328) );
NAND3_X1 U1002 ( .A1(G234), .A2(n1165), .A3(G221), .ZN(n1321) );
XOR2_X1 U1003 ( .A(n1330), .B(n1331), .Z(n1319) );
NOR2_X1 U1004 ( .A1(KEYINPUT14), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1005 ( .A(G137), .B(G146), .ZN(n1330) );
NAND2_X1 U1006 ( .A1(G217), .A2(G902), .ZN(n1315) );
INV_X1 U1007 ( .A(n1111), .ZN(n1307) );
NAND2_X1 U1008 ( .A1(n1333), .A2(n1334), .ZN(n1111) );
NAND2_X1 U1009 ( .A1(n1335), .A2(n1134), .ZN(n1334) );
NAND2_X1 U1010 ( .A1(n1336), .A2(n1220), .ZN(n1335) );
INV_X1 U1011 ( .A(G472), .ZN(n1220) );
NAND2_X1 U1012 ( .A1(n1147), .A2(n1336), .ZN(n1333) );
INV_X1 U1013 ( .A(KEYINPUT45), .ZN(n1336) );
NOR2_X1 U1014 ( .A1(n1134), .A2(G472), .ZN(n1147) );
NAND2_X1 U1015 ( .A1(n1337), .A2(n1197), .ZN(n1134) );
XNOR2_X1 U1016 ( .A(n1229), .B(n1338), .ZN(n1337) );
XOR2_X1 U1017 ( .A(n1228), .B(n1339), .Z(n1338) );
OR2_X1 U1018 ( .A1(n1224), .A2(n1222), .ZN(n1339) );
AND3_X1 U1019 ( .A1(G101), .A2(G210), .A3(n1340), .ZN(n1222) );
NOR2_X1 U1020 ( .A1(G101), .A2(n1341), .ZN(n1224) );
AND2_X1 U1021 ( .A1(n1340), .A2(G210), .ZN(n1341) );
INV_X1 U1022 ( .A(n1342), .ZN(n1229) );
AND4_X1 U1023 ( .A1(n1093), .A2(n1312), .A3(n1314), .A4(n1149), .ZN(n1254) );
NAND2_X1 U1024 ( .A1(G221), .A2(n1343), .ZN(n1149) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1197), .ZN(n1343) );
NAND2_X1 U1026 ( .A1(n1088), .A2(n1344), .ZN(n1314) );
NAND2_X1 U1027 ( .A1(n1299), .A2(n1185), .ZN(n1344) );
INV_X1 U1028 ( .A(G898), .ZN(n1185) );
AND3_X1 U1029 ( .A1(n1345), .A2(n1346), .A3(G953), .ZN(n1299) );
XNOR2_X1 U1030 ( .A(KEYINPUT63), .B(n1197), .ZN(n1345) );
NAND3_X1 U1031 ( .A1(n1346), .A2(n1165), .A3(G952), .ZN(n1088) );
NAND2_X1 U1032 ( .A1(G234), .A2(G237), .ZN(n1346) );
AND2_X1 U1033 ( .A1(n1105), .A2(n1104), .ZN(n1312) );
NAND3_X1 U1034 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1104) );
OR2_X1 U1035 ( .A1(n1350), .A2(n1245), .ZN(n1349) );
NAND3_X1 U1036 ( .A1(n1245), .A2(n1350), .A3(n1197), .ZN(n1348) );
NAND2_X1 U1037 ( .A1(G237), .A2(G210), .ZN(n1350) );
XOR2_X1 U1038 ( .A(n1351), .B(n1352), .Z(n1245) );
XOR2_X1 U1039 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1040 ( .A(KEYINPUT23), .B(n1355), .Z(n1354) );
NOR2_X1 U1041 ( .A1(G953), .A2(n1184), .ZN(n1355) );
INV_X1 U1042 ( .A(G224), .ZN(n1184) );
XNOR2_X1 U1043 ( .A(n1342), .B(n1180), .ZN(n1351) );
XNOR2_X1 U1044 ( .A(n1356), .B(n1357), .ZN(n1180) );
XNOR2_X1 U1045 ( .A(KEYINPUT37), .B(n1303), .ZN(n1357) );
XNOR2_X1 U1046 ( .A(G110), .B(n1241), .ZN(n1356) );
XNOR2_X1 U1047 ( .A(n1358), .B(n1182), .ZN(n1342) );
XNOR2_X1 U1048 ( .A(n1359), .B(n1360), .ZN(n1182) );
XOR2_X1 U1049 ( .A(G119), .B(G116), .Z(n1360) );
INV_X1 U1050 ( .A(G113), .ZN(n1359) );
NAND3_X1 U1051 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1358) );
OR2_X1 U1052 ( .A1(n1364), .A2(G128), .ZN(n1363) );
NAND3_X1 U1053 ( .A1(G128), .A2(n1364), .A3(KEYINPUT22), .ZN(n1362) );
NOR2_X1 U1054 ( .A1(KEYINPUT53), .A2(n1365), .ZN(n1364) );
NAND2_X1 U1055 ( .A1(n1365), .A2(n1366), .ZN(n1361) );
INV_X1 U1056 ( .A(KEYINPUT22), .ZN(n1366) );
XOR2_X1 U1057 ( .A(n1367), .B(n1368), .Z(n1365) );
XOR2_X1 U1058 ( .A(KEYINPUT7), .B(G143), .Z(n1368) );
NAND2_X1 U1059 ( .A1(KEYINPUT42), .A2(G146), .ZN(n1367) );
NAND2_X1 U1060 ( .A1(G902), .A2(G210), .ZN(n1347) );
NAND2_X1 U1061 ( .A1(G214), .A2(n1369), .ZN(n1105) );
OR2_X1 U1062 ( .A1(G237), .A2(G902), .ZN(n1369) );
INV_X1 U1063 ( .A(n1121), .ZN(n1093) );
XNOR2_X1 U1064 ( .A(n1152), .B(n1370), .ZN(n1121) );
XOR2_X1 U1065 ( .A(KEYINPUT28), .B(G469), .Z(n1370) );
NAND2_X1 U1066 ( .A1(n1371), .A2(n1197), .ZN(n1152) );
XOR2_X1 U1067 ( .A(n1372), .B(n1373), .Z(n1371) );
XOR2_X1 U1068 ( .A(n1374), .B(n1233), .Z(n1373) );
AND2_X1 U1069 ( .A1(G227), .A2(n1165), .ZN(n1233) );
NOR2_X1 U1070 ( .A1(KEYINPUT24), .A2(n1375), .ZN(n1374) );
NOR3_X1 U1071 ( .A1(n1376), .A2(n1377), .A3(n1378), .ZN(n1375) );
NOR2_X1 U1072 ( .A1(KEYINPUT52), .A2(n1327), .ZN(n1378) );
INV_X1 U1073 ( .A(G110), .ZN(n1327) );
AND3_X1 U1074 ( .A1(KEYINPUT52), .A2(n1379), .A3(n1380), .ZN(n1377) );
NOR2_X1 U1075 ( .A1(n1380), .A2(n1379), .ZN(n1376) );
INV_X1 U1076 ( .A(G140), .ZN(n1379) );
NOR2_X1 U1077 ( .A1(G110), .A2(KEYINPUT3), .ZN(n1380) );
NAND2_X1 U1078 ( .A1(n1239), .A2(n1381), .ZN(n1372) );
NAND2_X1 U1079 ( .A1(n1242), .A2(n1241), .ZN(n1381) );
OR2_X1 U1080 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
XNOR2_X1 U1081 ( .A(n1382), .B(n1383), .ZN(n1242) );
INV_X1 U1082 ( .A(n1162), .ZN(n1383) );
XNOR2_X1 U1083 ( .A(n1384), .B(n1385), .ZN(n1162) );
XNOR2_X1 U1084 ( .A(KEYINPUT7), .B(G146), .ZN(n1384) );
XOR2_X1 U1085 ( .A(n1228), .B(KEYINPUT1), .Z(n1382) );
NAND2_X1 U1086 ( .A1(n1386), .A2(n1387), .ZN(n1228) );
NAND2_X1 U1087 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1088 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
NAND2_X1 U1089 ( .A1(n1292), .A2(n1392), .ZN(n1391) );
INV_X1 U1090 ( .A(KEYINPUT11), .ZN(n1390) );
NAND2_X1 U1091 ( .A1(G131), .A2(n1393), .ZN(n1386) );
NAND2_X1 U1092 ( .A1(n1392), .A2(n1394), .ZN(n1393) );
OR2_X1 U1093 ( .A1(n1388), .A2(KEYINPUT11), .ZN(n1394) );
XNOR2_X1 U1094 ( .A(G134), .B(n1164), .ZN(n1388) );
INV_X1 U1095 ( .A(G137), .ZN(n1164) );
INV_X1 U1096 ( .A(KEYINPUT15), .ZN(n1392) );
XNOR2_X1 U1097 ( .A(n1395), .B(n1396), .ZN(n1241) );
XOR2_X1 U1098 ( .A(G104), .B(G101), .Z(n1396) );
XNOR2_X1 U1099 ( .A(G107), .B(KEYINPUT8), .ZN(n1395) );
INV_X1 U1100 ( .A(n1091), .ZN(n1274) );
NAND2_X1 U1101 ( .A1(n1265), .A2(n1266), .ZN(n1091) );
INV_X1 U1102 ( .A(n1138), .ZN(n1266) );
XNOR2_X1 U1103 ( .A(n1397), .B(G475), .ZN(n1138) );
NAND2_X1 U1104 ( .A1(n1398), .A2(n1212), .ZN(n1397) );
XNOR2_X1 U1105 ( .A(n1399), .B(n1400), .ZN(n1212) );
XOR2_X1 U1106 ( .A(n1401), .B(n1402), .Z(n1400) );
XOR2_X1 U1107 ( .A(n1403), .B(G143), .Z(n1402) );
NAND2_X1 U1108 ( .A1(KEYINPUT10), .A2(G146), .ZN(n1403) );
NAND2_X1 U1109 ( .A1(n1404), .A2(n1405), .ZN(n1401) );
OR2_X1 U1110 ( .A1(n1406), .A2(G104), .ZN(n1405) );
XOR2_X1 U1111 ( .A(n1407), .B(KEYINPUT19), .Z(n1404) );
NAND2_X1 U1112 ( .A1(G104), .A2(n1406), .ZN(n1407) );
XNOR2_X1 U1113 ( .A(G113), .B(n1303), .ZN(n1406) );
XOR2_X1 U1114 ( .A(n1161), .B(n1408), .Z(n1399) );
AND2_X1 U1115 ( .A1(G214), .A2(n1340), .ZN(n1408) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1340) );
XNOR2_X1 U1117 ( .A(n1332), .B(n1292), .ZN(n1161) );
INV_X1 U1118 ( .A(G131), .ZN(n1292) );
XNOR2_X1 U1119 ( .A(G140), .B(n1353), .ZN(n1332) );
XOR2_X1 U1120 ( .A(G125), .B(KEYINPUT21), .Z(n1353) );
XNOR2_X1 U1121 ( .A(G902), .B(KEYINPUT48), .ZN(n1398) );
XOR2_X1 U1122 ( .A(n1143), .B(G478), .Z(n1265) );
NAND2_X1 U1123 ( .A1(n1208), .A2(n1197), .ZN(n1143) );
INV_X1 U1124 ( .A(G902), .ZN(n1197) );
XOR2_X1 U1125 ( .A(n1409), .B(n1410), .Z(n1208) );
XNOR2_X1 U1126 ( .A(n1385), .B(n1411), .ZN(n1410) );
XOR2_X1 U1127 ( .A(n1412), .B(n1413), .Z(n1411) );
AND3_X1 U1128 ( .A1(G217), .A2(n1165), .A3(G234), .ZN(n1413) );
INV_X1 U1129 ( .A(G953), .ZN(n1165) );
NAND2_X1 U1130 ( .A1(KEYINPUT38), .A2(n1303), .ZN(n1412) );
INV_X1 U1131 ( .A(G122), .ZN(n1303) );
XOR2_X1 U1132 ( .A(G143), .B(G128), .Z(n1385) );
XNOR2_X1 U1133 ( .A(G107), .B(n1414), .ZN(n1409) );
XOR2_X1 U1134 ( .A(G134), .B(G116), .Z(n1414) );
endmodule


