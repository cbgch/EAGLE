//Key = 0101111111010101000100001100101100101000110000100000110110000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349;

XOR2_X1 U738 ( .A(n1023), .B(n1024), .Z(G9) );
NAND2_X1 U739 ( .A1(KEYINPUT8), .A2(G107), .ZN(n1024) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
XOR2_X1 U741 ( .A(KEYINPUT57), .B(n1027), .Z(n1026) );
NOR2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U743 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U746 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
INV_X1 U747 ( .A(n1039), .ZN(n1038) );
NOR2_X1 U748 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR4_X1 U750 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1046) );
XOR2_X1 U753 ( .A(KEYINPUT52), .B(n1052), .Z(n1051) );
NOR3_X1 U754 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1045) );
NOR3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1044) );
XOR2_X1 U756 ( .A(n1049), .B(KEYINPUT43), .Z(n1057) );
NOR3_X1 U757 ( .A1(n1054), .A2(n1059), .A3(n1060), .ZN(n1040) );
NOR3_X1 U758 ( .A1(n1049), .A2(n1061), .A3(n1062), .ZN(n1060) );
AND2_X1 U759 ( .A1(n1063), .A2(KEYINPUT56), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1059) );
NOR2_X1 U761 ( .A1(KEYINPUT56), .A2(n1066), .ZN(n1065) );
NOR4_X1 U762 ( .A1(n1067), .A2(n1049), .A3(n1054), .A4(n1043), .ZN(n1035) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U764 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U765 ( .A1(n1052), .A2(n1064), .A3(n1070), .A4(n1071), .ZN(n1030) );
NOR4_X1 U766 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
XOR2_X1 U767 ( .A(n1076), .B(n1077), .Z(n1074) );
NOR2_X1 U768 ( .A1(n1078), .A2(KEYINPUT12), .ZN(n1077) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1073) );
NOR2_X1 U770 ( .A1(G902), .A2(n1081), .ZN(n1079) );
XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(n1070) );
XOR2_X1 U772 ( .A(KEYINPUT58), .B(KEYINPUT54), .Z(n1083) );
XOR2_X1 U773 ( .A(n1084), .B(n1085), .Z(G72) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
AND2_X1 U775 ( .A1(G227), .A2(G900), .ZN(n1086) );
NAND2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1087), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND3_X1 U779 ( .A1(G900), .A2(n1092), .A3(G953), .ZN(n1088) );
XOR2_X1 U780 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U781 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U782 ( .A1(KEYINPUT55), .A2(n1097), .ZN(n1095) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1093) );
XOR2_X1 U784 ( .A(KEYINPUT48), .B(G140), .Z(n1099) );
NAND2_X1 U785 ( .A1(KEYINPUT1), .A2(n1100), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1101), .B(n1102), .Z(G69) );
NOR2_X1 U787 ( .A1(n1103), .A2(n1087), .ZN(n1102) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U789 ( .A(KEYINPUT53), .B(G898), .Z(n1105) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1087), .ZN(n1107) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND3_X1 U793 ( .A1(G898), .A2(n1110), .A3(G953), .ZN(n1106) );
XOR2_X1 U794 ( .A(n1111), .B(KEYINPUT63), .Z(n1110) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(G66) );
NOR3_X1 U796 ( .A1(n1078), .A2(n1114), .A3(n1115), .ZN(n1113) );
NOR3_X1 U797 ( .A1(n1116), .A2(n1076), .A3(n1117), .ZN(n1115) );
NOR2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1120), .A2(n1076), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1121), .ZN(G63) );
XOR2_X1 U801 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U802 ( .A1(n1124), .A2(n1117), .ZN(n1122) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1125), .ZN(G60) );
XOR2_X1 U804 ( .A(n1081), .B(n1126), .Z(n1125) );
NOR2_X1 U805 ( .A1(n1080), .A2(n1117), .ZN(n1126) );
XNOR2_X1 U806 ( .A(G104), .B(n1127), .ZN(G6) );
NOR2_X1 U807 ( .A1(n1112), .A2(n1128), .ZN(G57) );
XOR2_X1 U808 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U809 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U810 ( .A(n1133), .B(n1100), .Z(n1132) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1129) );
NOR2_X1 U812 ( .A1(n1136), .A2(n1117), .ZN(n1135) );
INV_X1 U813 ( .A(G472), .ZN(n1136) );
XOR2_X1 U814 ( .A(n1137), .B(KEYINPUT15), .Z(n1134) );
NAND2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U817 ( .A(KEYINPUT25), .B(n1142), .Z(n1138) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1112), .A2(n1143), .ZN(G54) );
XOR2_X1 U820 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U821 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U822 ( .A1(KEYINPUT45), .A2(n1148), .ZN(n1147) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1117), .ZN(n1146) );
INV_X1 U824 ( .A(G469), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1112), .A2(n1150), .ZN(G51) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1117), .ZN(n1154) );
NAND2_X1 U829 ( .A1(G902), .A2(n1032), .ZN(n1117) );
INV_X1 U830 ( .A(n1120), .ZN(n1032) );
NOR2_X1 U831 ( .A1(n1109), .A2(n1091), .ZN(n1120) );
NAND4_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1091) );
AND4_X1 U833 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NOR2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U836 ( .A1(n1168), .A2(n1068), .ZN(n1166) );
AND2_X1 U837 ( .A1(n1069), .A2(KEYINPUT28), .ZN(n1168) );
NOR4_X1 U838 ( .A1(n1169), .A2(n1050), .A3(n1066), .A4(n1170), .ZN(n1164) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
NOR2_X1 U840 ( .A1(KEYINPUT6), .A2(n1173), .ZN(n1172) );
NOR3_X1 U841 ( .A1(n1054), .A2(KEYINPUT28), .A3(n1174), .ZN(n1171) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1157) );
XOR2_X1 U843 ( .A(n1177), .B(KEYINPUT34), .Z(n1175) );
NAND2_X1 U844 ( .A1(KEYINPUT6), .A2(n1178), .ZN(n1156) );
NAND4_X1 U845 ( .A1(n1127), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1109) );
NOR4_X1 U846 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
INV_X1 U847 ( .A(n1186), .ZN(n1183) );
NAND2_X1 U848 ( .A1(n1027), .A2(n1187), .ZN(n1180) );
NAND2_X1 U849 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U850 ( .A1(n1068), .A2(n1190), .A3(n1063), .ZN(n1189) );
XNOR2_X1 U851 ( .A(n1025), .B(KEYINPUT50), .ZN(n1188) );
AND4_X1 U852 ( .A1(n1039), .A2(n1061), .A3(n1191), .A4(n1192), .ZN(n1025) );
NAND3_X1 U853 ( .A1(n1193), .A2(n1039), .A3(n1063), .ZN(n1127) );
INV_X1 U854 ( .A(G210), .ZN(n1155) );
NOR2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1153) );
XOR2_X1 U856 ( .A(KEYINPUT38), .B(n1196), .Z(n1195) );
AND2_X1 U857 ( .A1(G953), .A2(n1197), .ZN(n1112) );
XOR2_X1 U858 ( .A(KEYINPUT41), .B(G952), .Z(n1197) );
XNOR2_X1 U859 ( .A(n1178), .B(n1198), .ZN(G48) );
NAND2_X1 U860 ( .A1(KEYINPUT46), .A2(G146), .ZN(n1198) );
AND4_X1 U861 ( .A1(n1063), .A2(n1199), .A3(n1200), .A4(n1170), .ZN(n1178) );
XNOR2_X1 U862 ( .A(G143), .B(n1163), .ZN(G45) );
NAND4_X1 U863 ( .A1(n1170), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1163) );
NOR3_X1 U864 ( .A1(n1204), .A2(n1048), .A3(n1050), .ZN(n1203) );
INV_X1 U865 ( .A(n1082), .ZN(n1202) );
XOR2_X1 U866 ( .A(n1205), .B(n1206), .Z(G42) );
OR2_X1 U867 ( .A1(n1167), .A2(n1174), .ZN(n1206) );
INV_X1 U868 ( .A(n1069), .ZN(n1174) );
XNOR2_X1 U869 ( .A(G137), .B(n1162), .ZN(G39) );
NAND4_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1075), .ZN(n1162) );
XOR2_X1 U871 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U872 ( .A(n1161), .B(n1212), .Z(G36) );
NOR2_X1 U873 ( .A1(G134), .A2(KEYINPUT10), .ZN(n1212) );
NAND3_X1 U874 ( .A1(n1068), .A2(n1061), .A3(n1207), .ZN(n1161) );
XOR2_X1 U875 ( .A(G131), .B(n1213), .Z(G33) );
NOR3_X1 U876 ( .A1(n1167), .A2(KEYINPUT42), .A3(n1204), .ZN(n1213) );
NAND2_X1 U877 ( .A1(n1207), .A2(n1063), .ZN(n1167) );
AND3_X1 U878 ( .A1(n1200), .A2(n1170), .A3(n1052), .ZN(n1207) );
INV_X1 U879 ( .A(n1054), .ZN(n1052) );
NAND2_X1 U880 ( .A1(n1214), .A2(n1056), .ZN(n1054) );
INV_X1 U881 ( .A(n1058), .ZN(n1214) );
INV_X1 U882 ( .A(n1050), .ZN(n1200) );
XNOR2_X1 U883 ( .A(G128), .B(n1160), .ZN(G30) );
NAND4_X1 U884 ( .A1(n1199), .A2(n1061), .A3(n1191), .A4(n1170), .ZN(n1160) );
INV_X1 U885 ( .A(n1173), .ZN(n1199) );
XOR2_X1 U886 ( .A(n1140), .B(n1179), .Z(G3) );
NAND3_X1 U887 ( .A1(n1208), .A2(n1193), .A3(n1068), .ZN(n1179) );
XOR2_X1 U888 ( .A(G125), .B(n1215), .Z(G27) );
NOR2_X1 U889 ( .A1(n1048), .A2(n1177), .ZN(n1215) );
NAND4_X1 U890 ( .A1(n1063), .A2(n1064), .A3(n1069), .A4(n1170), .ZN(n1177) );
NAND2_X1 U891 ( .A1(n1034), .A2(n1216), .ZN(n1170) );
NAND4_X1 U892 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1218), .ZN(n1216) );
INV_X1 U893 ( .A(G900), .ZN(n1218) );
XOR2_X1 U894 ( .A(n1182), .B(n1219), .Z(G24) );
NOR2_X1 U895 ( .A1(KEYINPUT21), .A2(n1220), .ZN(n1219) );
INV_X1 U896 ( .A(G122), .ZN(n1220) );
AND3_X1 U897 ( .A1(n1190), .A2(n1039), .A3(n1221), .ZN(n1182) );
NOR3_X1 U898 ( .A1(n1048), .A2(n1222), .A3(n1082), .ZN(n1221) );
XOR2_X1 U899 ( .A(G119), .B(n1185), .Z(G21) );
NOR3_X1 U900 ( .A1(n1043), .A2(n1223), .A3(n1173), .ZN(n1185) );
NAND3_X1 U901 ( .A1(n1224), .A2(n1225), .A3(n1176), .ZN(n1173) );
NAND2_X1 U902 ( .A1(n1204), .A2(n1210), .ZN(n1225) );
NAND2_X1 U903 ( .A1(KEYINPUT11), .A2(n1226), .ZN(n1224) );
NAND2_X1 U904 ( .A1(n1211), .A2(n1075), .ZN(n1226) );
NAND3_X1 U905 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(G18) );
NAND2_X1 U906 ( .A1(KEYINPUT37), .A2(n1184), .ZN(n1229) );
INV_X1 U907 ( .A(n1230), .ZN(n1184) );
NAND3_X1 U908 ( .A1(n1230), .A2(n1231), .A3(G116), .ZN(n1228) );
NAND2_X1 U909 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
NAND2_X1 U910 ( .A1(n1234), .A2(n1231), .ZN(n1232) );
INV_X1 U911 ( .A(KEYINPUT37), .ZN(n1231) );
XOR2_X1 U912 ( .A(n1230), .B(KEYINPUT16), .Z(n1234) );
NAND4_X1 U913 ( .A1(n1068), .A2(n1190), .A3(n1061), .A4(n1176), .ZN(n1230) );
INV_X1 U914 ( .A(n1048), .ZN(n1176) );
XOR2_X1 U915 ( .A(n1235), .B(KEYINPUT23), .Z(n1048) );
NOR2_X1 U916 ( .A1(n1201), .A2(n1082), .ZN(n1061) );
INV_X1 U917 ( .A(n1223), .ZN(n1190) );
XNOR2_X1 U918 ( .A(G113), .B(n1236), .ZN(G15) );
NAND3_X1 U919 ( .A1(n1237), .A2(n1063), .A3(n1238), .ZN(n1236) );
NOR3_X1 U920 ( .A1(n1204), .A2(KEYINPUT14), .A3(n1223), .ZN(n1238) );
NAND2_X1 U921 ( .A1(n1064), .A2(n1192), .ZN(n1223) );
INV_X1 U922 ( .A(n1049), .ZN(n1064) );
NAND2_X1 U923 ( .A1(n1239), .A2(n1053), .ZN(n1049) );
INV_X1 U924 ( .A(n1055), .ZN(n1239) );
INV_X1 U925 ( .A(n1068), .ZN(n1204) );
NOR2_X1 U926 ( .A1(n1240), .A2(n1211), .ZN(n1068) );
INV_X1 U927 ( .A(n1066), .ZN(n1063) );
NAND2_X1 U928 ( .A1(n1082), .A2(n1201), .ZN(n1066) );
INV_X1 U929 ( .A(n1222), .ZN(n1201) );
XOR2_X1 U930 ( .A(n1235), .B(KEYINPUT40), .Z(n1237) );
NAND2_X1 U931 ( .A1(n1241), .A2(n1242), .ZN(G12) );
OR2_X1 U932 ( .A1(n1186), .A2(G110), .ZN(n1242) );
XOR2_X1 U933 ( .A(n1243), .B(KEYINPUT35), .Z(n1241) );
NAND2_X1 U934 ( .A1(G110), .A2(n1186), .ZN(n1243) );
NAND3_X1 U935 ( .A1(n1193), .A2(n1069), .A3(n1208), .ZN(n1186) );
INV_X1 U936 ( .A(n1043), .ZN(n1208) );
NAND2_X1 U937 ( .A1(n1082), .A2(n1222), .ZN(n1043) );
NOR2_X1 U938 ( .A1(n1244), .A2(n1072), .ZN(n1222) );
NOR3_X1 U939 ( .A1(G475), .A2(G902), .A3(n1081), .ZN(n1072) );
AND2_X1 U940 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U941 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
INV_X1 U942 ( .A(n1081), .ZN(n1247) );
XOR2_X1 U943 ( .A(n1249), .B(n1250), .Z(n1081) );
XOR2_X1 U944 ( .A(G104), .B(n1251), .Z(n1250) );
XOR2_X1 U945 ( .A(G143), .B(G131), .Z(n1251) );
XOR2_X1 U946 ( .A(n1252), .B(n1253), .Z(n1249) );
XOR2_X1 U947 ( .A(n1254), .B(n1255), .Z(n1252) );
AND3_X1 U948 ( .A1(G214), .A2(n1087), .A3(n1256), .ZN(n1255) );
NAND2_X1 U949 ( .A1(n1257), .A2(n1258), .ZN(n1254) );
OR2_X1 U950 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U951 ( .A(n1261), .B(KEYINPUT39), .Z(n1257) );
NAND2_X1 U952 ( .A1(n1259), .A2(n1260), .ZN(n1261) );
XNOR2_X1 U953 ( .A(n1262), .B(G140), .ZN(n1259) );
NAND2_X1 U954 ( .A1(KEYINPUT5), .A2(n1097), .ZN(n1262) );
INV_X1 U955 ( .A(G125), .ZN(n1097) );
XOR2_X1 U956 ( .A(n1080), .B(KEYINPUT19), .Z(n1245) );
INV_X1 U957 ( .A(G475), .ZN(n1080) );
XOR2_X1 U958 ( .A(n1124), .B(n1263), .Z(n1082) );
NOR2_X1 U959 ( .A1(G902), .A2(n1123), .ZN(n1263) );
XNOR2_X1 U960 ( .A(n1264), .B(n1265), .ZN(n1123) );
AND4_X1 U961 ( .A1(n1266), .A2(n1087), .A3(G234), .A4(G217), .ZN(n1265) );
INV_X1 U962 ( .A(KEYINPUT29), .ZN(n1266) );
NAND2_X1 U963 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
NAND2_X1 U964 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U965 ( .A(KEYINPUT7), .B(n1271), .Z(n1267) );
NOR2_X1 U966 ( .A1(n1270), .A2(n1269), .ZN(n1271) );
XOR2_X1 U967 ( .A(n1272), .B(n1273), .Z(n1269) );
XOR2_X1 U968 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U969 ( .A(G143), .B(KEYINPUT3), .ZN(n1274) );
NOR2_X1 U970 ( .A1(G134), .A2(KEYINPUT61), .ZN(n1272) );
XOR2_X1 U971 ( .A(G107), .B(n1276), .Z(n1270) );
XOR2_X1 U972 ( .A(G122), .B(G116), .Z(n1276) );
INV_X1 U973 ( .A(G478), .ZN(n1124) );
NAND2_X1 U974 ( .A1(n1277), .A2(n1278), .ZN(n1069) );
NAND2_X1 U975 ( .A1(n1039), .A2(n1210), .ZN(n1278) );
INV_X1 U976 ( .A(KEYINPUT11), .ZN(n1210) );
NOR2_X1 U977 ( .A1(n1075), .A2(n1211), .ZN(n1039) );
INV_X1 U978 ( .A(n1240), .ZN(n1075) );
NAND3_X1 U979 ( .A1(n1240), .A2(n1211), .A3(KEYINPUT11), .ZN(n1277) );
XNOR2_X1 U980 ( .A(n1078), .B(n1279), .ZN(n1211) );
NOR2_X1 U981 ( .A1(KEYINPUT20), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U982 ( .A(KEYINPUT17), .B(n1076), .ZN(n1280) );
NAND2_X1 U983 ( .A1(G217), .A2(n1281), .ZN(n1076) );
NOR2_X1 U984 ( .A1(n1119), .A2(G902), .ZN(n1078) );
INV_X1 U985 ( .A(n1116), .ZN(n1119) );
XOR2_X1 U986 ( .A(n1282), .B(n1283), .Z(n1116) );
XOR2_X1 U987 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U988 ( .A(G110), .B(n1286), .Z(n1285) );
AND3_X1 U989 ( .A1(G234), .A2(n1087), .A3(G221), .ZN(n1286) );
XOR2_X1 U990 ( .A(G137), .B(G125), .Z(n1284) );
XOR2_X1 U991 ( .A(n1287), .B(n1288), .Z(n1282) );
XOR2_X1 U992 ( .A(n1289), .B(n1260), .Z(n1288) );
INV_X1 U993 ( .A(n1275), .ZN(n1289) );
XOR2_X1 U994 ( .A(n1290), .B(n1291), .Z(n1287) );
NOR2_X1 U995 ( .A1(KEYINPUT26), .A2(n1205), .ZN(n1291) );
INV_X1 U996 ( .A(G140), .ZN(n1205) );
NAND2_X1 U997 ( .A1(KEYINPUT13), .A2(n1292), .ZN(n1290) );
XOR2_X1 U998 ( .A(n1293), .B(G472), .Z(n1240) );
NAND2_X1 U999 ( .A1(n1294), .A2(n1248), .ZN(n1293) );
XOR2_X1 U1000 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1001 ( .A(n1140), .B(n1297), .Z(n1296) );
XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(KEYINPUT31), .ZN(n1297) );
XNOR2_X1 U1003 ( .A(n1298), .B(n1141), .ZN(n1295) );
NAND3_X1 U1004 ( .A1(n1256), .A2(n1087), .A3(G210), .ZN(n1141) );
NAND2_X1 U1005 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U1006 ( .A1(n1301), .A2(n1131), .ZN(n1300) );
XOR2_X1 U1007 ( .A(KEYINPUT4), .B(n1302), .Z(n1299) );
NOR2_X1 U1008 ( .A1(n1301), .A2(n1131), .ZN(n1302) );
XNOR2_X1 U1009 ( .A(n1303), .B(n1304), .ZN(n1131) );
XOR2_X1 U1010 ( .A(n1305), .B(n1306), .Z(n1304) );
NOR2_X1 U1011 ( .A1(KEYINPUT27), .A2(n1292), .ZN(n1305) );
INV_X1 U1012 ( .A(G119), .ZN(n1292) );
XOR2_X1 U1013 ( .A(n1233), .B(KEYINPUT51), .Z(n1303) );
XOR2_X1 U1014 ( .A(n1133), .B(n1307), .Z(n1301) );
NOR2_X1 U1015 ( .A1(KEYINPUT22), .A2(n1100), .ZN(n1307) );
AND3_X1 U1016 ( .A1(n1191), .A2(n1192), .A3(n1027), .ZN(n1193) );
INV_X1 U1017 ( .A(n1235), .ZN(n1027) );
NAND2_X1 U1018 ( .A1(n1058), .A2(n1056), .ZN(n1235) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1308), .ZN(n1056) );
NAND2_X1 U1020 ( .A1(n1248), .A2(n1256), .ZN(n1308) );
NAND2_X1 U1021 ( .A1(n1309), .A2(n1310), .ZN(n1058) );
NAND2_X1 U1022 ( .A1(G210), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1023 ( .A1(n1248), .A2(n1312), .ZN(n1311) );
OR2_X1 U1024 ( .A1(n1313), .A2(n1256), .ZN(n1312) );
INV_X1 U1025 ( .A(G237), .ZN(n1256) );
NAND3_X1 U1026 ( .A1(n1314), .A2(n1248), .A3(n1313), .ZN(n1309) );
XNOR2_X1 U1027 ( .A(n1315), .B(n1151), .ZN(n1313) );
XNOR2_X1 U1028 ( .A(n1111), .B(KEYINPUT60), .ZN(n1151) );
XOR2_X1 U1029 ( .A(n1316), .B(n1317), .Z(n1111) );
XOR2_X1 U1030 ( .A(n1253), .B(n1318), .Z(n1317) );
XOR2_X1 U1031 ( .A(G110), .B(n1319), .Z(n1318) );
NOR2_X1 U1032 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XOR2_X1 U1033 ( .A(n1322), .B(KEYINPUT36), .Z(n1321) );
NAND2_X1 U1034 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1035 ( .A(KEYINPUT18), .B(n1325), .Z(n1323) );
XOR2_X1 U1036 ( .A(G122), .B(n1306), .Z(n1253) );
XOR2_X1 U1037 ( .A(G113), .B(KEYINPUT47), .Z(n1306) );
XOR2_X1 U1038 ( .A(n1233), .B(n1326), .Z(n1316) );
XOR2_X1 U1039 ( .A(KEYINPUT2), .B(G119), .Z(n1326) );
INV_X1 U1040 ( .A(G116), .ZN(n1233) );
XOR2_X1 U1041 ( .A(n1327), .B(KEYINPUT9), .Z(n1315) );
OR2_X1 U1042 ( .A1(n1196), .A2(n1194), .ZN(n1327) );
AND3_X1 U1043 ( .A1(n1328), .A2(n1087), .A3(G224), .ZN(n1194) );
NOR2_X1 U1044 ( .A1(n1328), .A2(n1329), .ZN(n1196) );
NOR2_X1 U1045 ( .A1(n1104), .A2(G953), .ZN(n1329) );
INV_X1 U1046 ( .A(G224), .ZN(n1104) );
XNOR2_X1 U1047 ( .A(n1133), .B(n1330), .ZN(n1328) );
XOR2_X1 U1048 ( .A(KEYINPUT0), .B(G125), .Z(n1330) );
XOR2_X1 U1049 ( .A(n1275), .B(n1331), .Z(n1133) );
NOR2_X1 U1050 ( .A1(KEYINPUT33), .A2(n1332), .ZN(n1331) );
NAND2_X1 U1051 ( .A1(G237), .A2(G210), .ZN(n1314) );
NAND2_X1 U1052 ( .A1(n1034), .A2(n1333), .ZN(n1192) );
NAND4_X1 U1053 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1334), .ZN(n1333) );
INV_X1 U1054 ( .A(G898), .ZN(n1334) );
NAND3_X1 U1055 ( .A1(n1217), .A2(n1087), .A3(G952), .ZN(n1034) );
NAND2_X1 U1056 ( .A1(G237), .A2(G234), .ZN(n1217) );
XOR2_X1 U1057 ( .A(n1050), .B(KEYINPUT24), .Z(n1191) );
NAND2_X1 U1058 ( .A1(n1055), .A2(n1053), .ZN(n1050) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1281), .ZN(n1053) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1248), .ZN(n1281) );
XNOR2_X1 U1061 ( .A(n1335), .B(G469), .ZN(n1055) );
NAND2_X1 U1062 ( .A1(n1336), .A2(n1248), .ZN(n1335) );
INV_X1 U1063 ( .A(G902), .ZN(n1248) );
XOR2_X1 U1064 ( .A(n1148), .B(n1144), .Z(n1336) );
XNOR2_X1 U1065 ( .A(n1337), .B(n1338), .ZN(n1144) );
XOR2_X1 U1066 ( .A(G140), .B(G110), .Z(n1338) );
XOR2_X1 U1067 ( .A(n1339), .B(n1340), .Z(n1337) );
INV_X1 U1068 ( .A(n1100), .ZN(n1340) );
XOR2_X1 U1069 ( .A(n1341), .B(n1342), .Z(n1100) );
XOR2_X1 U1070 ( .A(KEYINPUT44), .B(G137), .Z(n1342) );
XNOR2_X1 U1071 ( .A(G131), .B(G134), .ZN(n1341) );
NAND2_X1 U1072 ( .A1(G227), .A2(n1087), .ZN(n1339) );
INV_X1 U1073 ( .A(G953), .ZN(n1087) );
NAND3_X1 U1074 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1148) );
NAND2_X1 U1075 ( .A1(n1320), .A2(n1346), .ZN(n1345) );
INV_X1 U1076 ( .A(n1096), .ZN(n1346) );
NOR2_X1 U1077 ( .A1(n1325), .A2(n1324), .ZN(n1320) );
NAND3_X1 U1078 ( .A1(n1324), .A2(n1096), .A3(n1347), .ZN(n1344) );
NAND2_X1 U1079 ( .A1(n1325), .A2(n1348), .ZN(n1343) );
XOR2_X1 U1080 ( .A(n1324), .B(n1096), .Z(n1348) );
XNOR2_X1 U1081 ( .A(n1332), .B(n1349), .ZN(n1096) );
NOR2_X1 U1082 ( .A1(KEYINPUT32), .A2(n1275), .ZN(n1349) );
XNOR2_X1 U1083 ( .A(G128), .B(KEYINPUT30), .ZN(n1275) );
XOR2_X1 U1084 ( .A(G143), .B(n1260), .Z(n1332) );
XOR2_X1 U1085 ( .A(G146), .B(KEYINPUT62), .Z(n1260) );
XNOR2_X1 U1086 ( .A(n1140), .B(KEYINPUT59), .ZN(n1324) );
INV_X1 U1087 ( .A(G101), .ZN(n1140) );
INV_X1 U1088 ( .A(n1347), .ZN(n1325) );
XNOR2_X1 U1089 ( .A(G104), .B(G107), .ZN(n1347) );
endmodule


