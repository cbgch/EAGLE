//Key = 1101110010011011100001100110001001100100110100110001110101111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363;

XNOR2_X1 U739 ( .A(n1033), .B(n1034), .ZN(G9) );
NAND4_X1 U740 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(G75) );
NAND4_X1 U741 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1037) );
NOR3_X1 U742 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NAND3_X1 U743 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1043) );
XNOR2_X1 U744 ( .A(n1049), .B(n1050), .ZN(n1048) );
XOR2_X1 U745 ( .A(KEYINPUT2), .B(G472), .Z(n1050) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NAND2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U748 ( .A1(KEYINPUT40), .A2(n1055), .ZN(n1054) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
INV_X1 U750 ( .A(KEYINPUT40), .ZN(n1057) );
OR2_X1 U751 ( .A1(n1052), .A2(n1055), .ZN(n1046) );
NAND2_X1 U752 ( .A1(KEYINPUT22), .A2(n1056), .ZN(n1055) );
XOR2_X1 U753 ( .A(n1058), .B(KEYINPUT37), .Z(n1056) );
NOR3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1041) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1040) );
NAND2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1036) );
NAND2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U758 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND3_X1 U759 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1069) );
NAND2_X1 U760 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U761 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U762 ( .A1(n1078), .A2(n1079), .ZN(n1072) );
NAND2_X1 U763 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U764 ( .A1(KEYINPUT52), .A2(n1082), .ZN(n1081) );
OR3_X1 U765 ( .A1(n1083), .A2(KEYINPUT52), .A3(n1078), .ZN(n1071) );
NAND3_X1 U766 ( .A1(n1074), .A2(n1084), .A3(n1078), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND3_X1 U768 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND3_X1 U769 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
NAND2_X1 U770 ( .A1(n1059), .A2(n1093), .ZN(n1090) );
NAND2_X1 U771 ( .A1(n1094), .A2(n1061), .ZN(n1087) );
XOR2_X1 U772 ( .A(KEYINPUT25), .B(n1070), .Z(n1094) );
NAND2_X1 U773 ( .A1(n1070), .A2(n1095), .ZN(n1085) );
INV_X1 U774 ( .A(n1096), .ZN(n1064) );
XOR2_X1 U775 ( .A(n1097), .B(n1098), .Z(G72) );
NAND2_X1 U776 ( .A1(G953), .A2(n1099), .ZN(n1098) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1099) );
NAND4_X1 U778 ( .A1(KEYINPUT57), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1097) );
NAND3_X1 U779 ( .A1(n1103), .A2(n1104), .A3(n1038), .ZN(n1102) );
NAND2_X1 U780 ( .A1(G953), .A2(n1105), .ZN(n1101) );
NAND2_X1 U781 ( .A1(G900), .A2(n1103), .ZN(n1105) );
OR2_X1 U782 ( .A1(n1104), .A2(n1103), .ZN(n1100) );
XNOR2_X1 U783 ( .A(n1106), .B(n1107), .ZN(n1103) );
XOR2_X1 U784 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U785 ( .A1(KEYINPUT55), .A2(n1110), .ZN(n1108) );
XOR2_X1 U786 ( .A(n1111), .B(KEYINPUT24), .Z(n1106) );
NAND2_X1 U787 ( .A1(n1112), .A2(n1113), .ZN(n1104) );
XNOR2_X1 U788 ( .A(n1114), .B(KEYINPUT0), .ZN(n1112) );
XOR2_X1 U789 ( .A(n1115), .B(n1116), .Z(G69) );
XOR2_X1 U790 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U791 ( .A1(n1119), .A2(n1038), .ZN(n1118) );
NOR2_X1 U792 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U793 ( .A1(n1122), .A2(n1123), .ZN(n1117) );
NAND2_X1 U794 ( .A1(G953), .A2(n1121), .ZN(n1123) );
XNOR2_X1 U795 ( .A(n1124), .B(n1125), .ZN(n1122) );
XOR2_X1 U796 ( .A(KEYINPUT39), .B(n1126), .Z(n1125) );
NAND2_X1 U797 ( .A1(n1038), .A2(n1127), .ZN(n1115) );
NOR2_X1 U798 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U799 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U800 ( .A(KEYINPUT53), .B(n1132), .Z(n1131) );
NOR2_X1 U801 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U802 ( .A1(n1135), .A2(n1136), .ZN(G63) );
XNOR2_X1 U803 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U804 ( .A1(n1139), .A2(n1134), .ZN(n1137) );
NOR2_X1 U805 ( .A1(n1038), .A2(n1140), .ZN(n1135) );
XOR2_X1 U806 ( .A(KEYINPUT62), .B(G952), .Z(n1140) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1141), .ZN(G60) );
XOR2_X1 U808 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U809 ( .A1(n1144), .A2(n1134), .ZN(n1142) );
XNOR2_X1 U810 ( .A(G104), .B(n1145), .ZN(G6) );
NAND2_X1 U811 ( .A1(KEYINPUT3), .A2(n1146), .ZN(n1145) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1147), .ZN(G57) );
XOR2_X1 U813 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U814 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U815 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U816 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND3_X1 U817 ( .A1(G472), .A2(G902), .A3(n1156), .ZN(n1155) );
XNOR2_X1 U818 ( .A(n1035), .B(KEYINPUT13), .ZN(n1156) );
NAND4_X1 U819 ( .A1(n1157), .A2(n1158), .A3(G472), .A4(n1159), .ZN(n1152) );
NAND2_X1 U820 ( .A1(n1134), .A2(n1160), .ZN(n1158) );
INV_X1 U821 ( .A(KEYINPUT13), .ZN(n1160) );
NAND2_X1 U822 ( .A1(KEYINPUT13), .A2(n1161), .ZN(n1157) );
NAND2_X1 U823 ( .A1(n1035), .A2(G902), .ZN(n1161) );
INV_X1 U824 ( .A(n1162), .ZN(n1035) );
XNOR2_X1 U825 ( .A(G101), .B(KEYINPUT63), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1128), .A2(n1163), .ZN(G54) );
XOR2_X1 U827 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U828 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U829 ( .A1(n1168), .A2(KEYINPUT1), .ZN(n1167) );
XOR2_X1 U830 ( .A(n1169), .B(KEYINPUT16), .Z(n1168) );
XOR2_X1 U831 ( .A(n1170), .B(n1171), .Z(n1164) );
NOR2_X1 U832 ( .A1(n1172), .A2(n1134), .ZN(n1171) );
INV_X1 U833 ( .A(G469), .ZN(n1172) );
NAND4_X1 U834 ( .A1(KEYINPUT12), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1170) );
NAND3_X1 U835 ( .A1(KEYINPUT51), .A2(n1176), .A3(n1177), .ZN(n1175) );
OR2_X1 U836 ( .A1(n1177), .A2(n1176), .ZN(n1174) );
NOR2_X1 U837 ( .A1(G110), .A2(KEYINPUT36), .ZN(n1176) );
NAND2_X1 U838 ( .A1(G110), .A2(n1178), .ZN(n1173) );
INV_X1 U839 ( .A(KEYINPUT51), .ZN(n1178) );
NOR2_X1 U840 ( .A1(n1128), .A2(n1179), .ZN(G51) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U842 ( .A(n1182), .B(n1183), .ZN(n1181) );
XNOR2_X1 U843 ( .A(n1184), .B(n1185), .ZN(n1180) );
NOR2_X1 U844 ( .A1(n1063), .A2(n1134), .ZN(n1185) );
NAND2_X1 U845 ( .A1(G902), .A2(n1162), .ZN(n1134) );
NAND3_X1 U846 ( .A1(n1113), .A2(n1114), .A3(n1186), .ZN(n1162) );
INV_X1 U847 ( .A(n1127), .ZN(n1186) );
NAND2_X1 U848 ( .A1(n1187), .A2(n1188), .ZN(n1127) );
NOR4_X1 U849 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NOR4_X1 U850 ( .A1(n1146), .A2(n1034), .A3(n1193), .A4(n1194), .ZN(n1187) );
NOR3_X1 U851 ( .A1(n1083), .A2(n1077), .A3(n1195), .ZN(n1194) );
NOR3_X1 U852 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
NAND3_X1 U853 ( .A1(n1199), .A2(n1200), .A3(n1074), .ZN(n1196) );
NAND2_X1 U854 ( .A1(KEYINPUT21), .A2(n1195), .ZN(n1200) );
NAND2_X1 U855 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
INV_X1 U856 ( .A(KEYINPUT21), .ZN(n1202) );
NAND3_X1 U857 ( .A1(n1203), .A2(n1091), .A3(n1068), .ZN(n1201) );
AND3_X1 U858 ( .A1(n1204), .A2(n1074), .A3(n1205), .ZN(n1034) );
AND3_X1 U859 ( .A1(n1205), .A2(n1074), .A3(n1206), .ZN(n1146) );
NOR3_X1 U860 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1114) );
AND3_X1 U861 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NAND2_X1 U862 ( .A1(n1213), .A2(n1214), .ZN(n1210) );
AND3_X1 U863 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1113) );
NAND2_X1 U864 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U865 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U866 ( .A1(n1222), .A2(n1078), .ZN(n1221) );
NAND2_X1 U867 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
XNOR2_X1 U868 ( .A(KEYINPUT42), .B(n1076), .ZN(n1224) );
NOR2_X1 U869 ( .A1(n1038), .A2(G952), .ZN(n1128) );
XNOR2_X1 U870 ( .A(G146), .B(n1215), .ZN(G48) );
NAND3_X1 U871 ( .A1(n1222), .A2(n1206), .A3(n1225), .ZN(n1215) );
XNOR2_X1 U872 ( .A(G143), .B(n1216), .ZN(G45) );
NAND4_X1 U873 ( .A1(n1225), .A2(n1082), .A3(n1226), .A4(n1045), .ZN(n1216) );
AND3_X1 U874 ( .A1(n1095), .A2(n1211), .A3(n1212), .ZN(n1225) );
XNOR2_X1 U875 ( .A(n1177), .B(n1227), .ZN(G42) );
NOR3_X1 U876 ( .A1(n1228), .A2(n1080), .A3(n1076), .ZN(n1227) );
XNOR2_X1 U877 ( .A(G137), .B(n1229), .ZN(G39) );
NAND4_X1 U878 ( .A1(KEYINPUT41), .A2(n1218), .A3(n1222), .A4(n1078), .ZN(n1229) );
INV_X1 U879 ( .A(n1228), .ZN(n1218) );
XOR2_X1 U880 ( .A(G134), .B(n1207), .Z(G36) );
NOR3_X1 U881 ( .A1(n1083), .A2(n1077), .A3(n1228), .ZN(n1207) );
XOR2_X1 U882 ( .A(n1230), .B(n1208), .Z(G33) );
NOR3_X1 U883 ( .A1(n1076), .A2(n1083), .A3(n1228), .ZN(n1208) );
NAND3_X1 U884 ( .A1(n1095), .A2(n1211), .A3(n1070), .ZN(n1228) );
AND2_X1 U885 ( .A1(n1093), .A2(n1231), .ZN(n1070) );
XNOR2_X1 U886 ( .A(G131), .B(KEYINPUT58), .ZN(n1230) );
XOR2_X1 U887 ( .A(G128), .B(n1232), .Z(G30) );
NOR3_X1 U888 ( .A1(n1214), .A2(n1233), .A3(n1234), .ZN(n1232) );
XNOR2_X1 U889 ( .A(n1212), .B(KEYINPUT6), .ZN(n1234) );
NAND3_X1 U890 ( .A1(n1204), .A2(n1235), .A3(n1222), .ZN(n1214) );
XOR2_X1 U891 ( .A(n1192), .B(n1236), .Z(G3) );
NOR2_X1 U892 ( .A1(KEYINPUT28), .A2(n1237), .ZN(n1236) );
AND3_X1 U893 ( .A1(n1078), .A2(n1205), .A3(n1082), .ZN(n1192) );
XOR2_X1 U894 ( .A(n1238), .B(n1239), .Z(G27) );
NOR2_X1 U895 ( .A1(KEYINPUT10), .A2(n1240), .ZN(n1239) );
INV_X1 U896 ( .A(G125), .ZN(n1240) );
NAND2_X1 U897 ( .A1(n1241), .A2(n1242), .ZN(n1238) );
OR4_X1 U898 ( .A1(n1091), .A2(n1233), .A3(n1213), .A4(KEYINPUT7), .ZN(n1242) );
INV_X1 U899 ( .A(n1212), .ZN(n1091) );
NAND3_X1 U900 ( .A1(n1212), .A2(n1243), .A3(KEYINPUT7), .ZN(n1241) );
OR2_X1 U901 ( .A1(n1213), .A2(n1233), .ZN(n1243) );
INV_X1 U902 ( .A(n1211), .ZN(n1233) );
NAND2_X1 U903 ( .A1(n1096), .A2(n1244), .ZN(n1211) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1246), .ZN(n1244) );
INV_X1 U905 ( .A(G900), .ZN(n1246) );
NAND3_X1 U906 ( .A1(n1068), .A2(n1223), .A3(n1206), .ZN(n1213) );
INV_X1 U907 ( .A(n1076), .ZN(n1206) );
XNOR2_X1 U908 ( .A(G122), .B(n1247), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1248), .A2(n1074), .A3(n1226), .A4(n1045), .ZN(n1247) );
INV_X1 U910 ( .A(n1198), .ZN(n1226) );
AND2_X1 U911 ( .A1(n1249), .A2(n1250), .ZN(n1074) );
XNOR2_X1 U912 ( .A(n1251), .B(n1191), .ZN(G21) );
AND3_X1 U913 ( .A1(n1248), .A2(n1078), .A3(n1222), .ZN(n1191) );
AND2_X1 U914 ( .A1(n1252), .A2(n1044), .ZN(n1222) );
INV_X1 U915 ( .A(n1195), .ZN(n1248) );
XNOR2_X1 U916 ( .A(n1253), .B(n1254), .ZN(G18) );
NOR3_X1 U917 ( .A1(n1195), .A2(n1255), .A3(n1077), .ZN(n1254) );
INV_X1 U918 ( .A(n1204), .ZN(n1077) );
NOR2_X1 U919 ( .A1(n1045), .A2(n1198), .ZN(n1204) );
XNOR2_X1 U920 ( .A(n1039), .B(KEYINPUT59), .ZN(n1198) );
XNOR2_X1 U921 ( .A(n1082), .B(KEYINPUT38), .ZN(n1255) );
INV_X1 U922 ( .A(n1083), .ZN(n1082) );
NAND2_X1 U923 ( .A1(n1256), .A2(n1257), .ZN(G15) );
OR2_X1 U924 ( .A1(n1258), .A2(n1190), .ZN(n1257) );
XOR2_X1 U925 ( .A(n1259), .B(KEYINPUT18), .Z(n1256) );
NAND2_X1 U926 ( .A1(n1190), .A2(n1258), .ZN(n1259) );
NOR3_X1 U927 ( .A1(n1083), .A2(n1195), .A3(n1076), .ZN(n1190) );
NAND2_X1 U928 ( .A1(n1260), .A2(n1045), .ZN(n1076) );
NAND3_X1 U929 ( .A1(n1212), .A2(n1203), .A3(n1068), .ZN(n1195) );
AND2_X1 U930 ( .A1(n1089), .A2(n1092), .ZN(n1068) );
NAND2_X1 U931 ( .A1(n1252), .A2(n1250), .ZN(n1083) );
XOR2_X1 U932 ( .A(n1044), .B(KEYINPUT14), .Z(n1250) );
INV_X1 U933 ( .A(n1249), .ZN(n1252) );
XOR2_X1 U934 ( .A(G110), .B(n1189), .Z(G12) );
AND3_X1 U935 ( .A1(n1223), .A2(n1205), .A3(n1078), .ZN(n1189) );
AND2_X1 U936 ( .A1(n1260), .A2(n1197), .ZN(n1078) );
INV_X1 U937 ( .A(n1045), .ZN(n1197) );
XNOR2_X1 U938 ( .A(n1261), .B(n1262), .ZN(n1045) );
XNOR2_X1 U939 ( .A(KEYINPUT20), .B(n1144), .ZN(n1262) );
INV_X1 U940 ( .A(G475), .ZN(n1144) );
OR2_X1 U941 ( .A1(n1143), .A2(G902), .ZN(n1261) );
XNOR2_X1 U942 ( .A(n1263), .B(n1264), .ZN(n1143) );
XOR2_X1 U943 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U944 ( .A(n1267), .B(n1268), .ZN(n1266) );
AND3_X1 U945 ( .A1(G214), .A2(n1038), .A3(n1269), .ZN(n1268) );
XNOR2_X1 U946 ( .A(G131), .B(n1270), .ZN(n1265) );
XOR2_X1 U947 ( .A(n1109), .B(n1271), .Z(n1263) );
XOR2_X1 U948 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U949 ( .A(G125), .B(G140), .ZN(n1109) );
XOR2_X1 U950 ( .A(n1039), .B(KEYINPUT50), .Z(n1260) );
XNOR2_X1 U951 ( .A(n1274), .B(n1139), .ZN(n1039) );
INV_X1 U952 ( .A(G478), .ZN(n1139) );
NAND2_X1 U953 ( .A1(n1138), .A2(n1275), .ZN(n1274) );
XNOR2_X1 U954 ( .A(KEYINPUT8), .B(n1276), .ZN(n1275) );
XOR2_X1 U955 ( .A(n1277), .B(n1278), .Z(n1138) );
XOR2_X1 U956 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U957 ( .A1(G217), .A2(n1281), .ZN(n1280) );
NAND2_X1 U958 ( .A1(n1282), .A2(n1283), .ZN(n1279) );
NAND2_X1 U959 ( .A1(G122), .A2(n1253), .ZN(n1283) );
INV_X1 U960 ( .A(G116), .ZN(n1253) );
XOR2_X1 U961 ( .A(n1284), .B(KEYINPUT35), .Z(n1282) );
NAND2_X1 U962 ( .A1(G116), .A2(n1270), .ZN(n1284) );
XOR2_X1 U963 ( .A(n1285), .B(n1286), .Z(n1277) );
XNOR2_X1 U964 ( .A(G134), .B(n1033), .ZN(n1286) );
NAND2_X1 U965 ( .A1(KEYINPUT26), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U966 ( .A(n1288), .B(G128), .ZN(n1287) );
AND3_X1 U967 ( .A1(n1235), .A2(n1203), .A3(n1212), .ZN(n1205) );
NOR2_X1 U968 ( .A1(n1059), .A2(n1093), .ZN(n1212) );
NOR2_X1 U969 ( .A1(n1289), .A2(n1060), .ZN(n1093) );
NOR2_X1 U970 ( .A1(n1063), .A2(n1062), .ZN(n1060) );
AND2_X1 U971 ( .A1(n1290), .A2(n1062), .ZN(n1289) );
AND2_X1 U972 ( .A1(n1291), .A2(n1292), .ZN(n1062) );
XNOR2_X1 U973 ( .A(KEYINPUT11), .B(n1276), .ZN(n1292) );
XOR2_X1 U974 ( .A(n1293), .B(n1183), .Z(n1291) );
XNOR2_X1 U975 ( .A(n1294), .B(n1126), .ZN(n1183) );
XNOR2_X1 U976 ( .A(n1270), .B(n1295), .ZN(n1126) );
NOR2_X1 U977 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1295) );
INV_X1 U978 ( .A(G122), .ZN(n1270) );
NAND2_X1 U979 ( .A1(KEYINPUT46), .A2(n1124), .ZN(n1294) );
XNOR2_X1 U980 ( .A(n1296), .B(n1297), .ZN(n1124) );
NOR2_X1 U981 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR3_X1 U982 ( .A1(n1033), .A2(G104), .A3(n1300), .ZN(n1299) );
NOR2_X1 U983 ( .A1(G107), .A2(n1301), .ZN(n1298) );
NOR2_X1 U984 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NOR2_X1 U985 ( .A1(n1304), .A2(n1267), .ZN(n1303) );
NOR2_X1 U986 ( .A1(G104), .A2(n1305), .ZN(n1302) );
NOR2_X1 U987 ( .A1(n1300), .A2(n1304), .ZN(n1305) );
XOR2_X1 U988 ( .A(KEYINPUT34), .B(KEYINPUT15), .Z(n1304) );
XOR2_X1 U989 ( .A(KEYINPUT54), .B(KEYINPUT49), .Z(n1300) );
XNOR2_X1 U990 ( .A(n1306), .B(n1237), .ZN(n1296) );
NAND2_X1 U991 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U992 ( .A1(n1309), .A2(n1251), .ZN(n1307) );
XOR2_X1 U993 ( .A(KEYINPUT61), .B(n1310), .Z(n1309) );
NAND2_X1 U994 ( .A1(n1311), .A2(n1312), .ZN(n1293) );
NAND2_X1 U995 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U996 ( .A1(n1315), .A2(n1184), .ZN(n1311) );
XNOR2_X1 U997 ( .A(KEYINPUT56), .B(n1313), .ZN(n1315) );
INV_X1 U998 ( .A(n1182), .ZN(n1313) );
XOR2_X1 U999 ( .A(G125), .B(n1316), .Z(n1182) );
NOR2_X1 U1000 ( .A1(G953), .A2(n1120), .ZN(n1316) );
INV_X1 U1001 ( .A(G224), .ZN(n1120) );
XOR2_X1 U1002 ( .A(n1063), .B(KEYINPUT44), .Z(n1290) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1317), .ZN(n1063) );
INV_X1 U1004 ( .A(n1231), .ZN(n1059) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1317), .ZN(n1231) );
NAND2_X1 U1006 ( .A1(n1269), .A2(n1276), .ZN(n1317) );
NAND2_X1 U1007 ( .A1(n1096), .A2(n1318), .ZN(n1203) );
NAND4_X1 U1008 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1121), .ZN(n1318) );
INV_X1 U1009 ( .A(G898), .ZN(n1121) );
NAND3_X1 U1010 ( .A1(n1245), .A2(n1038), .A3(G952), .ZN(n1096) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1245) );
XOR2_X1 U1012 ( .A(n1095), .B(KEYINPUT9), .Z(n1235) );
NOR2_X1 U1013 ( .A1(n1089), .A2(n1061), .ZN(n1095) );
INV_X1 U1014 ( .A(n1092), .ZN(n1061) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1319), .ZN(n1092) );
XOR2_X1 U1016 ( .A(n1052), .B(n1058), .Z(n1089) );
XNOR2_X1 U1017 ( .A(G469), .B(KEYINPUT4), .ZN(n1058) );
NAND2_X1 U1018 ( .A1(n1320), .A2(n1276), .ZN(n1052) );
XOR2_X1 U1019 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1020 ( .A(n1169), .B(n1166), .ZN(n1322) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1038), .ZN(n1166) );
XOR2_X1 U1022 ( .A(n1323), .B(n1324), .Z(n1169) );
XNOR2_X1 U1023 ( .A(n1267), .B(n1325), .ZN(n1324) );
XNOR2_X1 U1024 ( .A(KEYINPUT29), .B(n1033), .ZN(n1325) );
INV_X1 U1025 ( .A(G107), .ZN(n1033) );
INV_X1 U1026 ( .A(G104), .ZN(n1267) );
XNOR2_X1 U1027 ( .A(n1326), .B(n1110), .ZN(n1323) );
XNOR2_X1 U1028 ( .A(n1111), .B(n1237), .ZN(n1326) );
NAND2_X1 U1029 ( .A1(n1327), .A2(n1328), .ZN(n1111) );
NAND2_X1 U1030 ( .A1(G128), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1031 ( .A(KEYINPUT5), .B(n1330), .Z(n1327) );
NOR2_X1 U1032 ( .A1(G128), .A2(n1329), .ZN(n1330) );
XOR2_X1 U1033 ( .A(G146), .B(n1331), .Z(n1329) );
NOR2_X1 U1034 ( .A1(KEYINPUT45), .A2(n1288), .ZN(n1331) );
XNOR2_X1 U1035 ( .A(G110), .B(G140), .ZN(n1321) );
INV_X1 U1036 ( .A(n1080), .ZN(n1223) );
NAND2_X1 U1037 ( .A1(n1332), .A2(n1249), .ZN(n1080) );
XOR2_X1 U1038 ( .A(G472), .B(n1333), .Z(n1249) );
NOR2_X1 U1039 ( .A1(n1049), .A2(KEYINPUT17), .ZN(n1333) );
AND2_X1 U1040 ( .A1(n1334), .A2(n1276), .ZN(n1049) );
NAND2_X1 U1041 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1042 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XNOR2_X1 U1043 ( .A(n1237), .B(n1339), .ZN(n1338) );
INV_X1 U1044 ( .A(G101), .ZN(n1237) );
XNOR2_X1 U1045 ( .A(n1154), .B(KEYINPUT30), .ZN(n1337) );
INV_X1 U1046 ( .A(n1159), .ZN(n1154) );
XOR2_X1 U1047 ( .A(n1340), .B(KEYINPUT19), .Z(n1335) );
NAND2_X1 U1048 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1049 ( .A(KEYINPUT30), .B(n1159), .ZN(n1342) );
NAND3_X1 U1050 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1159) );
OR2_X1 U1051 ( .A1(n1308), .A2(n1346), .ZN(n1345) );
OR2_X1 U1052 ( .A1(n1251), .A2(n1310), .ZN(n1308) );
NAND3_X1 U1053 ( .A1(n1346), .A2(n1310), .A3(G119), .ZN(n1344) );
NAND2_X1 U1054 ( .A1(n1347), .A2(n1251), .ZN(n1343) );
XOR2_X1 U1055 ( .A(n1346), .B(n1310), .Z(n1347) );
XOR2_X1 U1056 ( .A(G116), .B(n1273), .Z(n1310) );
XNOR2_X1 U1057 ( .A(n1258), .B(KEYINPUT33), .ZN(n1273) );
INV_X1 U1058 ( .A(G113), .ZN(n1258) );
XOR2_X1 U1059 ( .A(n1110), .B(n1314), .Z(n1346) );
INV_X1 U1060 ( .A(n1184), .ZN(n1314) );
XNOR2_X1 U1061 ( .A(n1348), .B(n1272), .ZN(n1184) );
XNOR2_X1 U1062 ( .A(n1288), .B(G146), .ZN(n1272) );
INV_X1 U1063 ( .A(G143), .ZN(n1288) );
XNOR2_X1 U1064 ( .A(G128), .B(KEYINPUT43), .ZN(n1348) );
XNOR2_X1 U1065 ( .A(G131), .B(n1349), .ZN(n1110) );
XOR2_X1 U1066 ( .A(G137), .B(G134), .Z(n1349) );
XNOR2_X1 U1067 ( .A(G101), .B(n1339), .ZN(n1341) );
NOR2_X1 U1068 ( .A1(KEYINPUT27), .A2(n1150), .ZN(n1339) );
NAND3_X1 U1069 ( .A1(n1350), .A2(n1269), .A3(G210), .ZN(n1150) );
INV_X1 U1070 ( .A(G237), .ZN(n1269) );
XNOR2_X1 U1071 ( .A(KEYINPUT47), .B(n1038), .ZN(n1350) );
XOR2_X1 U1072 ( .A(KEYINPUT32), .B(n1044), .Z(n1332) );
XOR2_X1 U1073 ( .A(n1351), .B(n1133), .Z(n1044) );
NAND2_X1 U1074 ( .A1(G217), .A2(n1319), .ZN(n1133) );
NAND2_X1 U1075 ( .A1(G234), .A2(n1276), .ZN(n1319) );
NAND2_X1 U1076 ( .A1(n1130), .A2(n1276), .ZN(n1351) );
INV_X1 U1077 ( .A(G902), .ZN(n1276) );
XNOR2_X1 U1078 ( .A(n1352), .B(n1353), .ZN(n1130) );
XOR2_X1 U1079 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1080 ( .A(n1251), .B(G110), .ZN(n1355) );
INV_X1 U1081 ( .A(G119), .ZN(n1251) );
XOR2_X1 U1082 ( .A(G137), .B(G128), .Z(n1354) );
XOR2_X1 U1083 ( .A(n1356), .B(n1357), .Z(n1352) );
NOR2_X1 U1084 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NOR2_X1 U1085 ( .A1(n1177), .A2(n1360), .ZN(n1359) );
XNOR2_X1 U1086 ( .A(G125), .B(KEYINPUT60), .ZN(n1360) );
INV_X1 U1087 ( .A(G140), .ZN(n1177) );
NOR2_X1 U1088 ( .A1(G140), .A2(n1361), .ZN(n1358) );
XNOR2_X1 U1089 ( .A(G125), .B(KEYINPUT31), .ZN(n1361) );
XOR2_X1 U1090 ( .A(n1362), .B(n1363), .Z(n1356) );
NOR2_X1 U1091 ( .A1(G146), .A2(KEYINPUT48), .ZN(n1363) );
NAND2_X1 U1092 ( .A1(n1281), .A2(G221), .ZN(n1362) );
AND2_X1 U1093 ( .A1(G234), .A2(n1038), .ZN(n1281) );
INV_X1 U1094 ( .A(G953), .ZN(n1038) );
endmodule


