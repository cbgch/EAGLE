//Key = 0010000111101010100000000000010100001101110001001011000100100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360;

XOR2_X1 U751 ( .A(n1037), .B(G107), .Z(G9) );
NAND2_X1 U752 ( .A1(KEYINPUT37), .A2(n1038), .ZN(n1037) );
NOR2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1041), .A2(n1042), .A3(G953), .A4(n1043), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
XOR2_X1 U756 ( .A(n1046), .B(KEYINPUT30), .Z(n1044) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND4_X1 U759 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
OR2_X1 U760 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U761 ( .A1(n1057), .A2(n1058), .A3(n1055), .ZN(n1053) );
NAND2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1056), .A2(n1061), .ZN(n1049) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U765 ( .A1(n1055), .A2(n1064), .A3(n1051), .ZN(n1063) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1066) );
XOR2_X1 U768 ( .A(KEYINPUT24), .B(n1071), .Z(n1069) );
NAND2_X1 U769 ( .A1(n1052), .A2(n1072), .ZN(n1062) );
INV_X1 U770 ( .A(n1073), .ZN(n1047) );
NOR3_X1 U771 ( .A1(n1043), .A2(G953), .A3(G952), .ZN(n1039) );
AND4_X1 U772 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1043) );
NOR4_X1 U773 ( .A1(n1078), .A2(n1079), .A3(n1059), .A4(n1070), .ZN(n1077) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND3_X1 U775 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1078) );
NOR4_X1 U776 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1076) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1091), .B(KEYINPUT63), .ZN(n1090) );
NOR2_X1 U779 ( .A1(G475), .A2(n1092), .ZN(n1087) );
XNOR2_X1 U780 ( .A(n1091), .B(KEYINPUT28), .ZN(n1092) );
NOR3_X1 U781 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1086) );
AND2_X1 U782 ( .A1(n1093), .A2(n1095), .ZN(n1085) );
INV_X1 U783 ( .A(KEYINPUT50), .ZN(n1093) );
XOR2_X1 U784 ( .A(n1096), .B(KEYINPUT54), .Z(n1075) );
NAND2_X1 U785 ( .A1(n1081), .A2(n1080), .ZN(n1096) );
XOR2_X1 U786 ( .A(G469), .B(KEYINPUT18), .Z(n1081) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1074) );
XOR2_X1 U788 ( .A(n1099), .B(n1100), .Z(n1097) );
NOR2_X1 U789 ( .A1(KEYINPUT49), .A2(n1101), .ZN(n1100) );
XNOR2_X1 U790 ( .A(G472), .B(KEYINPUT47), .ZN(n1099) );
NAND2_X1 U791 ( .A1(n1102), .A2(n1103), .ZN(G72) );
NAND3_X1 U792 ( .A1(n1104), .A2(n1105), .A3(G953), .ZN(n1103) );
XOR2_X1 U793 ( .A(n1106), .B(KEYINPUT1), .Z(n1102) );
NAND2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U795 ( .A1(G953), .A2(n1104), .ZN(n1108) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1104) );
XNOR2_X1 U797 ( .A(n1105), .B(n1109), .ZN(n1107) );
NOR3_X1 U798 ( .A1(n1110), .A2(KEYINPUT56), .A3(G953), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1105) );
NAND2_X1 U800 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1111) );
XOR2_X1 U802 ( .A(G140), .B(n1116), .Z(n1115) );
NOR2_X1 U803 ( .A1(KEYINPUT42), .A2(n1117), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U805 ( .A(n1120), .B(n1121), .ZN(n1118) );
NAND2_X1 U806 ( .A1(KEYINPUT51), .A2(n1122), .ZN(n1120) );
NAND2_X1 U807 ( .A1(KEYINPUT29), .A2(n1123), .ZN(n1114) );
INV_X1 U808 ( .A(G125), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(G69) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U811 ( .A1(KEYINPUT12), .A2(n1128), .ZN(n1127) );
NAND2_X1 U812 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U813 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1126) );
NAND2_X1 U814 ( .A1(G953), .A2(n1134), .ZN(n1133) );
NAND2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
OR2_X1 U817 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
INV_X1 U818 ( .A(n1141), .ZN(n1135) );
NAND2_X1 U819 ( .A1(n1142), .A2(n1141), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1139), .B(n1140), .Z(n1142) );
NAND2_X1 U821 ( .A1(G953), .A2(n1143), .ZN(n1124) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1144), .A2(n1150), .ZN(G63) );
XOR2_X1 U827 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U828 ( .A1(n1148), .A2(G478), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1144), .A2(n1153), .ZN(G60) );
NOR3_X1 U830 ( .A1(n1091), .A2(n1154), .A3(n1155), .ZN(n1153) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1089), .ZN(n1156) );
NOR2_X1 U833 ( .A1(n1042), .A2(n1129), .ZN(n1158) );
AND3_X1 U834 ( .A1(n1157), .A2(G475), .A3(n1148), .ZN(n1154) );
XNOR2_X1 U835 ( .A(n1159), .B(n1160), .ZN(G6) );
NOR2_X1 U836 ( .A1(n1144), .A2(n1161), .ZN(G57) );
XOR2_X1 U837 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U838 ( .A1(n1148), .A2(G472), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1144), .A2(n1164), .ZN(G54) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U841 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U842 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
INV_X1 U844 ( .A(n1169), .ZN(n1172) );
XNOR2_X1 U845 ( .A(n1173), .B(n1174), .ZN(n1169) );
NOR2_X1 U846 ( .A1(KEYINPUT11), .A2(n1175), .ZN(n1174) );
XNOR2_X1 U847 ( .A(KEYINPUT20), .B(n1170), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1176), .B(n1177), .Z(n1170) );
NOR2_X1 U849 ( .A1(KEYINPUT25), .A2(n1178), .ZN(n1177) );
XNOR2_X1 U850 ( .A(n1179), .B(KEYINPUT27), .ZN(n1178) );
NAND2_X1 U851 ( .A1(n1148), .A2(G469), .ZN(n1165) );
INV_X1 U852 ( .A(n1180), .ZN(n1148) );
NOR2_X1 U853 ( .A1(n1144), .A2(n1181), .ZN(G51) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR3_X1 U855 ( .A1(n1180), .A2(KEYINPUT32), .A3(n1184), .ZN(n1183) );
INV_X1 U856 ( .A(G210), .ZN(n1184) );
NAND2_X1 U857 ( .A1(G902), .A2(n1185), .ZN(n1180) );
NAND2_X1 U858 ( .A1(n1045), .A2(n1110), .ZN(n1185) );
INV_X1 U859 ( .A(n1042), .ZN(n1110) );
NAND3_X1 U860 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1042) );
AND3_X1 U861 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1187) );
NAND2_X1 U863 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U864 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND3_X1 U866 ( .A1(n1200), .A2(n1201), .A3(n1056), .ZN(n1199) );
XOR2_X1 U867 ( .A(KEYINPUT53), .B(n1072), .Z(n1200) );
XNOR2_X1 U868 ( .A(n1202), .B(KEYINPUT46), .ZN(n1194) );
OR2_X1 U869 ( .A1(n1067), .A2(n1203), .ZN(n1186) );
NAND2_X1 U870 ( .A1(n1204), .A2(n1205), .ZN(n1067) );
NAND2_X1 U871 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
INV_X1 U872 ( .A(n1129), .ZN(n1045) );
NAND4_X1 U873 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1129) );
NOR4_X1 U874 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
INV_X1 U875 ( .A(n1038), .ZN(n1213) );
NAND2_X1 U876 ( .A1(n1216), .A2(n1217), .ZN(n1038) );
NOR3_X1 U877 ( .A1(n1160), .A2(n1218), .A3(n1219), .ZN(n1210) );
AND2_X1 U878 ( .A1(KEYINPUT39), .A2(n1220), .ZN(n1219) );
NOR4_X1 U879 ( .A1(KEYINPUT39), .A2(n1221), .A3(n1222), .A4(n1098), .ZN(n1218) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
AND2_X1 U881 ( .A1(n1196), .A2(n1217), .ZN(n1160) );
NOR3_X1 U882 ( .A1(n1225), .A2(n1226), .A3(n1058), .ZN(n1217) );
NOR2_X1 U883 ( .A1(n1130), .A2(G952), .ZN(n1144) );
XNOR2_X1 U884 ( .A(G146), .B(n1227), .ZN(G48) );
NAND4_X1 U885 ( .A1(KEYINPUT14), .A2(n1228), .A3(n1196), .A4(n1192), .ZN(n1227) );
XOR2_X1 U886 ( .A(n1229), .B(n1230), .Z(G45) );
XOR2_X1 U887 ( .A(KEYINPUT8), .B(G143), .Z(n1230) );
NAND2_X1 U888 ( .A1(n1202), .A2(n1192), .ZN(n1229) );
AND3_X1 U889 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1202) );
XOR2_X1 U890 ( .A(G140), .B(n1234), .Z(G42) );
NOR2_X1 U891 ( .A1(KEYINPUT3), .A2(n1189), .ZN(n1234) );
NAND4_X1 U892 ( .A1(n1204), .A2(n1235), .A3(n1196), .A4(n1072), .ZN(n1189) );
XOR2_X1 U893 ( .A(n1191), .B(n1236), .Z(G39) );
NAND2_X1 U894 ( .A1(KEYINPUT31), .A2(G137), .ZN(n1236) );
NAND2_X1 U895 ( .A1(n1052), .A2(n1228), .ZN(n1191) );
AND2_X1 U896 ( .A1(n1204), .A2(n1071), .ZN(n1052) );
XOR2_X1 U897 ( .A(G134), .B(n1237), .Z(G36) );
NOR4_X1 U898 ( .A1(KEYINPUT13), .A2(n1207), .A3(n1238), .A4(n1203), .ZN(n1237) );
INV_X1 U899 ( .A(n1216), .ZN(n1207) );
XOR2_X1 U900 ( .A(n1239), .B(n1240), .Z(G33) );
NOR2_X1 U901 ( .A1(KEYINPUT21), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U902 ( .A(G131), .B(KEYINPUT19), .ZN(n1241) );
NOR4_X1 U903 ( .A1(n1242), .A2(n1243), .A3(n1206), .A4(n1238), .ZN(n1239) );
INV_X1 U904 ( .A(n1204), .ZN(n1238) );
NOR2_X1 U905 ( .A1(n1244), .A2(n1070), .ZN(n1204) );
NOR2_X1 U906 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
INV_X1 U907 ( .A(KEYINPUT5), .ZN(n1246) );
NOR4_X1 U908 ( .A1(n1058), .A2(n1098), .A3(n1201), .A4(n1055), .ZN(n1245) );
NOR2_X1 U909 ( .A1(KEYINPUT5), .A2(n1233), .ZN(n1242) );
INV_X1 U910 ( .A(n1203), .ZN(n1233) );
NAND3_X1 U911 ( .A1(n1051), .A2(n1226), .A3(n1235), .ZN(n1203) );
XNOR2_X1 U912 ( .A(G128), .B(n1190), .ZN(G30) );
NAND3_X1 U913 ( .A1(n1216), .A2(n1192), .A3(n1228), .ZN(n1190) );
INV_X1 U914 ( .A(n1198), .ZN(n1228) );
NAND2_X1 U915 ( .A1(n1235), .A2(n1247), .ZN(n1198) );
NOR2_X1 U916 ( .A1(n1058), .A2(n1248), .ZN(n1235) );
INV_X1 U917 ( .A(n1249), .ZN(n1058) );
XNOR2_X1 U918 ( .A(G101), .B(n1250), .ZN(G3) );
NOR2_X1 U919 ( .A1(n1212), .A2(KEYINPUT38), .ZN(n1250) );
AND4_X1 U920 ( .A1(n1226), .A2(n1071), .A3(n1249), .A4(n1251), .ZN(n1212) );
XNOR2_X1 U921 ( .A(G125), .B(n1252), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1253), .A2(n1056), .A3(n1254), .A4(n1072), .ZN(n1252) );
NOR2_X1 U923 ( .A1(n1248), .A2(n1223), .ZN(n1254) );
INV_X1 U924 ( .A(n1192), .ZN(n1223) );
INV_X1 U925 ( .A(n1201), .ZN(n1248) );
NAND2_X1 U926 ( .A1(n1073), .A2(n1255), .ZN(n1201) );
NAND2_X1 U927 ( .A1(n1256), .A2(n1113), .ZN(n1255) );
XOR2_X1 U928 ( .A(KEYINPUT58), .B(G900), .Z(n1113) );
XNOR2_X1 U929 ( .A(n1196), .B(KEYINPUT7), .ZN(n1253) );
XOR2_X1 U930 ( .A(n1220), .B(n1257), .Z(G24) );
NOR2_X1 U931 ( .A1(KEYINPUT17), .A2(n1258), .ZN(n1257) );
NOR2_X1 U932 ( .A1(n1222), .A2(n1225), .ZN(n1220) );
NAND4_X1 U933 ( .A1(n1056), .A2(n1055), .A3(n1231), .A4(n1232), .ZN(n1222) );
XNOR2_X1 U934 ( .A(G119), .B(n1208), .ZN(G21) );
NAND4_X1 U935 ( .A1(n1247), .A2(n1056), .A3(n1259), .A4(n1224), .ZN(n1208) );
AND2_X1 U936 ( .A1(n1226), .A2(n1260), .ZN(n1247) );
XNOR2_X1 U937 ( .A(KEYINPUT23), .B(n1051), .ZN(n1260) );
XNOR2_X1 U938 ( .A(G116), .B(n1209), .ZN(G18) );
NAND2_X1 U939 ( .A1(n1261), .A2(n1216), .ZN(n1209) );
NOR2_X1 U940 ( .A1(n1231), .A2(n1262), .ZN(n1216) );
XOR2_X1 U941 ( .A(G113), .B(n1215), .Z(G15) );
AND2_X1 U942 ( .A1(n1196), .A2(n1261), .ZN(n1215) );
AND3_X1 U943 ( .A1(n1226), .A2(n1251), .A3(n1056), .ZN(n1261) );
NOR2_X1 U944 ( .A1(n1263), .A2(n1059), .ZN(n1056) );
INV_X1 U945 ( .A(n1225), .ZN(n1251) );
NAND3_X1 U946 ( .A1(n1051), .A2(n1224), .A3(n1192), .ZN(n1225) );
INV_X1 U947 ( .A(n1206), .ZN(n1196) );
NAND2_X1 U948 ( .A1(n1262), .A2(n1231), .ZN(n1206) );
INV_X1 U949 ( .A(n1232), .ZN(n1262) );
XOR2_X1 U950 ( .A(G110), .B(n1214), .Z(G12) );
AND4_X1 U951 ( .A1(n1259), .A2(n1072), .A3(n1249), .A4(n1224), .ZN(n1214) );
NAND2_X1 U952 ( .A1(n1264), .A2(n1073), .ZN(n1224) );
NAND3_X1 U953 ( .A1(n1265), .A2(n1130), .A3(G952), .ZN(n1073) );
NAND2_X1 U954 ( .A1(n1256), .A2(n1134), .ZN(n1264) );
INV_X1 U955 ( .A(G898), .ZN(n1134) );
AND3_X1 U956 ( .A1(G902), .A2(n1265), .A3(G953), .ZN(n1256) );
NAND2_X1 U957 ( .A1(G237), .A2(G234), .ZN(n1265) );
NOR2_X1 U958 ( .A1(n1060), .A2(n1059), .ZN(n1249) );
AND2_X1 U959 ( .A1(G221), .A2(n1266), .ZN(n1059) );
INV_X1 U960 ( .A(n1263), .ZN(n1060) );
XNOR2_X1 U961 ( .A(n1080), .B(G469), .ZN(n1263) );
NAND2_X1 U962 ( .A1(n1267), .A2(n1268), .ZN(n1080) );
XOR2_X1 U963 ( .A(n1269), .B(n1270), .Z(n1267) );
XNOR2_X1 U964 ( .A(n1175), .B(n1271), .ZN(n1270) );
INV_X1 U965 ( .A(n1179), .ZN(n1271) );
XOR2_X1 U966 ( .A(n1122), .B(n1272), .Z(n1179) );
XNOR2_X1 U967 ( .A(G101), .B(n1273), .ZN(n1272) );
NAND2_X1 U968 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
OR2_X1 U969 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U970 ( .A(n1278), .B(KEYINPUT57), .Z(n1274) );
NAND2_X1 U971 ( .A1(n1277), .A2(n1276), .ZN(n1278) );
XOR2_X1 U972 ( .A(G107), .B(KEYINPUT2), .Z(n1276) );
XOR2_X1 U973 ( .A(n1279), .B(n1280), .Z(n1122) );
XNOR2_X1 U974 ( .A(G110), .B(G140), .ZN(n1175) );
XNOR2_X1 U975 ( .A(n1176), .B(n1173), .ZN(n1269) );
NAND2_X1 U976 ( .A1(G227), .A2(n1130), .ZN(n1173) );
NOR2_X1 U977 ( .A1(n1051), .A2(n1226), .ZN(n1072) );
INV_X1 U978 ( .A(n1055), .ZN(n1226) );
XOR2_X1 U979 ( .A(G472), .B(n1281), .Z(n1055) );
NOR2_X1 U980 ( .A1(n1101), .A2(KEYINPUT43), .ZN(n1281) );
AND2_X1 U981 ( .A1(n1282), .A2(n1268), .ZN(n1101) );
XOR2_X1 U982 ( .A(n1163), .B(KEYINPUT52), .Z(n1282) );
XOR2_X1 U983 ( .A(n1283), .B(n1284), .Z(n1163) );
XOR2_X1 U984 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U985 ( .A(G101), .B(G113), .ZN(n1286) );
NAND2_X1 U986 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
OR2_X1 U987 ( .A1(n1289), .A2(G116), .ZN(n1288) );
XOR2_X1 U988 ( .A(n1290), .B(KEYINPUT33), .Z(n1287) );
NAND2_X1 U989 ( .A1(G116), .A2(n1289), .ZN(n1290) );
XOR2_X1 U990 ( .A(n1176), .B(n1291), .Z(n1283) );
XOR2_X1 U991 ( .A(n1292), .B(n1293), .Z(n1291) );
NAND3_X1 U992 ( .A1(n1294), .A2(n1130), .A3(G210), .ZN(n1292) );
NAND3_X1 U993 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1176) );
NAND2_X1 U994 ( .A1(KEYINPUT4), .A2(n1119), .ZN(n1297) );
NAND3_X1 U995 ( .A1(n1298), .A2(n1299), .A3(n1121), .ZN(n1296) );
INV_X1 U996 ( .A(KEYINPUT4), .ZN(n1299) );
OR2_X1 U997 ( .A1(n1121), .A2(n1298), .ZN(n1295) );
NOR2_X1 U998 ( .A1(KEYINPUT34), .A2(n1119), .ZN(n1298) );
XOR2_X1 U999 ( .A(G137), .B(n1300), .Z(n1119) );
INV_X1 U1000 ( .A(n1098), .ZN(n1051) );
XNOR2_X1 U1001 ( .A(n1301), .B(n1149), .ZN(n1098) );
AND2_X1 U1002 ( .A1(G217), .A2(n1266), .ZN(n1149) );
NAND2_X1 U1003 ( .A1(G234), .A2(n1268), .ZN(n1266) );
NAND2_X1 U1004 ( .A1(n1147), .A2(n1268), .ZN(n1301) );
XOR2_X1 U1005 ( .A(n1302), .B(n1303), .Z(n1147) );
XOR2_X1 U1006 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1007 ( .A(n1306), .B(G119), .ZN(n1305) );
INV_X1 U1008 ( .A(G128), .ZN(n1306) );
XOR2_X1 U1009 ( .A(G140), .B(G137), .Z(n1304) );
XOR2_X1 U1010 ( .A(n1307), .B(n1308), .Z(n1302) );
XNOR2_X1 U1011 ( .A(n1309), .B(n1310), .ZN(n1308) );
NOR2_X1 U1012 ( .A1(G125), .A2(KEYINPUT22), .ZN(n1310) );
NAND2_X1 U1013 ( .A1(KEYINPUT41), .A2(n1280), .ZN(n1309) );
XNOR2_X1 U1014 ( .A(G110), .B(n1311), .ZN(n1307) );
AND3_X1 U1015 ( .A1(G221), .A2(n1130), .A3(G234), .ZN(n1311) );
INV_X1 U1016 ( .A(n1065), .ZN(n1259) );
NAND2_X1 U1017 ( .A1(n1071), .A2(n1192), .ZN(n1065) );
NOR2_X1 U1018 ( .A1(n1070), .A2(n1068), .ZN(n1192) );
INV_X1 U1019 ( .A(n1244), .ZN(n1068) );
NAND3_X1 U1020 ( .A1(n1312), .A2(n1313), .A3(n1082), .ZN(n1244) );
NAND2_X1 U1021 ( .A1(n1094), .A2(n1095), .ZN(n1082) );
NAND2_X1 U1022 ( .A1(n1095), .A2(n1314), .ZN(n1313) );
OR3_X1 U1023 ( .A1(n1095), .A2(n1094), .A3(n1314), .ZN(n1312) );
INV_X1 U1024 ( .A(KEYINPUT36), .ZN(n1314) );
NOR2_X1 U1025 ( .A1(n1182), .A2(G902), .ZN(n1094) );
XOR2_X1 U1026 ( .A(n1315), .B(n1316), .Z(n1182) );
XOR2_X1 U1027 ( .A(n1293), .B(n1317), .Z(n1316) );
XNOR2_X1 U1028 ( .A(G125), .B(KEYINPUT45), .ZN(n1317) );
NAND3_X1 U1029 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1293) );
NAND2_X1 U1030 ( .A1(KEYINPUT15), .A2(n1321), .ZN(n1320) );
INV_X1 U1031 ( .A(n1322), .ZN(n1321) );
OR3_X1 U1032 ( .A1(n1323), .A2(KEYINPUT15), .A3(G128), .ZN(n1319) );
NAND2_X1 U1033 ( .A1(G128), .A2(n1323), .ZN(n1318) );
NAND2_X1 U1034 ( .A1(KEYINPUT55), .A2(n1322), .ZN(n1323) );
XOR2_X1 U1035 ( .A(G143), .B(n1280), .Z(n1322) );
XNOR2_X1 U1036 ( .A(n1324), .B(n1141), .ZN(n1315) );
XOR2_X1 U1037 ( .A(G110), .B(n1258), .Z(n1141) );
XOR2_X1 U1038 ( .A(n1325), .B(n1326), .Z(n1324) );
AND2_X1 U1039 ( .A1(n1130), .A2(G224), .ZN(n1326) );
NAND2_X1 U1040 ( .A1(n1327), .A2(n1137), .ZN(n1325) );
NAND2_X1 U1041 ( .A1(n1140), .A2(n1139), .ZN(n1137) );
XOR2_X1 U1042 ( .A(KEYINPUT9), .B(n1328), .Z(n1327) );
NOR2_X1 U1043 ( .A1(n1140), .A2(n1139), .ZN(n1328) );
XNOR2_X1 U1044 ( .A(n1329), .B(n1330), .ZN(n1139) );
NOR2_X1 U1045 ( .A1(KEYINPUT61), .A2(n1289), .ZN(n1330) );
INV_X1 U1046 ( .A(G119), .ZN(n1289) );
XNOR2_X1 U1047 ( .A(G113), .B(G116), .ZN(n1329) );
XNOR2_X1 U1048 ( .A(n1331), .B(n1277), .ZN(n1140) );
XOR2_X1 U1049 ( .A(n1159), .B(KEYINPUT16), .Z(n1277) );
XNOR2_X1 U1050 ( .A(G101), .B(G107), .ZN(n1331) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1332), .ZN(n1095) );
AND2_X1 U1052 ( .A1(G214), .A2(n1332), .ZN(n1070) );
NAND2_X1 U1053 ( .A1(n1294), .A2(n1268), .ZN(n1332) );
NOR2_X1 U1054 ( .A1(n1232), .A2(n1231), .ZN(n1071) );
XNOR2_X1 U1055 ( .A(n1091), .B(n1089), .ZN(n1231) );
INV_X1 U1056 ( .A(G475), .ZN(n1089) );
NOR2_X1 U1057 ( .A1(n1157), .A2(G902), .ZN(n1091) );
XOR2_X1 U1058 ( .A(n1333), .B(n1334), .Z(n1157) );
NOR2_X1 U1059 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NOR2_X1 U1060 ( .A1(G104), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1061 ( .A(n1338), .B(n1339), .ZN(n1337) );
XOR2_X1 U1062 ( .A(KEYINPUT35), .B(KEYINPUT26), .Z(n1339) );
NOR2_X1 U1063 ( .A1(n1338), .A2(n1159), .ZN(n1335) );
INV_X1 U1064 ( .A(G104), .ZN(n1159) );
XNOR2_X1 U1065 ( .A(n1340), .B(n1341), .ZN(n1338) );
XNOR2_X1 U1066 ( .A(G113), .B(n1342), .ZN(n1341) );
NAND2_X1 U1067 ( .A1(KEYINPUT40), .A2(n1258), .ZN(n1342) );
XNOR2_X1 U1068 ( .A(G125), .B(n1343), .ZN(n1340) );
XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G140), .Z(n1343) );
XOR2_X1 U1070 ( .A(n1344), .B(n1345), .Z(n1333) );
NOR2_X1 U1071 ( .A1(KEYINPUT62), .A2(n1280), .ZN(n1345) );
XOR2_X1 U1072 ( .A(G146), .B(KEYINPUT60), .Z(n1280) );
NAND2_X1 U1073 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
OR2_X1 U1074 ( .A1(n1121), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1075 ( .A(n1349), .B(KEYINPUT44), .Z(n1346) );
NAND2_X1 U1076 ( .A1(n1348), .A2(n1121), .ZN(n1349) );
INV_X1 U1077 ( .A(G131), .ZN(n1121) );
XOR2_X1 U1078 ( .A(G143), .B(n1350), .Z(n1348) );
AND3_X1 U1079 ( .A1(G214), .A2(n1130), .A3(n1294), .ZN(n1350) );
INV_X1 U1080 ( .A(G237), .ZN(n1294) );
NAND2_X1 U1081 ( .A1(n1351), .A2(n1083), .ZN(n1232) );
NAND3_X1 U1082 ( .A1(n1352), .A2(n1268), .A3(n1152), .ZN(n1083) );
INV_X1 U1083 ( .A(G478), .ZN(n1352) );
XOR2_X1 U1084 ( .A(n1084), .B(KEYINPUT0), .Z(n1351) );
NAND2_X1 U1085 ( .A1(G478), .A2(n1353), .ZN(n1084) );
NAND2_X1 U1086 ( .A1(n1152), .A2(n1268), .ZN(n1353) );
INV_X1 U1087 ( .A(G902), .ZN(n1268) );
XNOR2_X1 U1088 ( .A(n1354), .B(n1355), .ZN(n1152) );
XOR2_X1 U1089 ( .A(n1300), .B(n1279), .Z(n1355) );
XOR2_X1 U1090 ( .A(G128), .B(G143), .Z(n1279) );
XOR2_X1 U1091 ( .A(G134), .B(KEYINPUT10), .Z(n1300) );
XOR2_X1 U1092 ( .A(n1356), .B(n1357), .Z(n1354) );
NOR2_X1 U1093 ( .A1(KEYINPUT6), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1094 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1095 ( .A(KEYINPUT48), .B(n1258), .ZN(n1360) );
INV_X1 U1096 ( .A(G122), .ZN(n1258) );
XNOR2_X1 U1097 ( .A(G107), .B(G116), .ZN(n1359) );
NAND3_X1 U1098 ( .A1(G217), .A2(n1130), .A3(G234), .ZN(n1356) );
INV_X1 U1099 ( .A(G953), .ZN(n1130) );
endmodule


