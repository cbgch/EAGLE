//Key = 1101100101011110000111101010001111011110000000010000010000010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352;

XOR2_X1 U742 ( .A(n1027), .B(n1028), .Z(G9) );
NOR2_X1 U743 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U744 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
XOR2_X1 U745 ( .A(KEYINPUT54), .B(n1034), .Z(n1033) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1052), .A2(n1057), .A3(n1048), .ZN(n1041) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
AND2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR4_X1 U760 ( .A1(n1062), .A2(n1048), .A3(n1044), .A4(n1052), .ZN(n1037) );
INV_X1 U761 ( .A(n1063), .ZN(n1044) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U764 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND3_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1031) );
NOR3_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
XNOR2_X1 U767 ( .A(n1074), .B(KEYINPUT37), .ZN(n1071) );
XOR2_X1 U768 ( .A(n1075), .B(KEYINPUT61), .Z(n1068) );
NAND4_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
XOR2_X1 U771 ( .A(n1082), .B(KEYINPUT20), .Z(n1081) );
NAND2_X1 U772 ( .A1(G478), .A2(n1083), .ZN(n1082) );
NOR2_X1 U773 ( .A1(G478), .A2(n1083), .ZN(n1080) );
XNOR2_X1 U774 ( .A(n1084), .B(n1085), .ZN(n1077) );
XOR2_X1 U775 ( .A(n1086), .B(G472), .Z(n1076) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(G72) );
NAND2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U778 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
XOR2_X1 U779 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1091) );
NAND3_X1 U781 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1089) );
XNOR2_X1 U782 ( .A(n1095), .B(n1094), .ZN(n1098) );
XNOR2_X1 U783 ( .A(n1099), .B(n1100), .ZN(n1094) );
NOR2_X1 U784 ( .A1(KEYINPUT25), .A2(n1101), .ZN(n1100) );
NAND2_X1 U785 ( .A1(KEYINPUT19), .A2(n1102), .ZN(n1099) );
XNOR2_X1 U786 ( .A(n1103), .B(n1104), .ZN(n1095) );
XOR2_X1 U787 ( .A(KEYINPUT2), .B(G131), .Z(n1104) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NAND2_X1 U789 ( .A1(G125), .A2(n1107), .ZN(n1106) );
XOR2_X1 U790 ( .A(n1108), .B(KEYINPUT17), .Z(n1105) );
NAND2_X1 U791 ( .A1(G140), .A2(n1109), .ZN(n1108) );
INV_X1 U792 ( .A(G125), .ZN(n1109) );
NAND2_X1 U793 ( .A1(n1110), .A2(n1111), .ZN(n1096) );
XOR2_X1 U794 ( .A(KEYINPUT48), .B(n1112), .Z(n1111) );
NAND2_X1 U795 ( .A1(n1092), .A2(n1113), .ZN(n1087) );
NAND2_X1 U796 ( .A1(G953), .A2(n1114), .ZN(n1113) );
INV_X1 U797 ( .A(n1115), .ZN(n1092) );
XOR2_X1 U798 ( .A(n1116), .B(n1117), .Z(G69) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U800 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U801 ( .A1(G224), .A2(G898), .ZN(n1120) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1121) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
INV_X1 U806 ( .A(KEYINPUT60), .ZN(n1128) );
NAND3_X1 U807 ( .A1(n1129), .A2(n1130), .A3(KEYINPUT60), .ZN(n1125) );
NOR2_X1 U808 ( .A1(n1131), .A2(G953), .ZN(n1116) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1084), .A2(n1136), .ZN(n1135) );
NOR3_X1 U812 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G63) );
AND2_X1 U813 ( .A1(KEYINPUT13), .A2(n1132), .ZN(n1139) );
NOR3_X1 U814 ( .A1(KEYINPUT13), .A2(n1097), .A3(n1140), .ZN(n1138) );
INV_X1 U815 ( .A(G952), .ZN(n1140) );
NOR3_X1 U816 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1137) );
NOR3_X1 U817 ( .A1(n1144), .A2(n1145), .A3(n1136), .ZN(n1143) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1145), .ZN(n1147) );
XNOR2_X1 U820 ( .A(G478), .B(KEYINPUT23), .ZN(n1145) );
INV_X1 U821 ( .A(n1032), .ZN(n1148) );
INV_X1 U822 ( .A(n1144), .ZN(n1146) );
INV_X1 U823 ( .A(n1083), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1132), .A2(n1149), .ZN(G60) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U826 ( .A1(n1152), .A2(n1136), .ZN(n1150) );
INV_X1 U827 ( .A(G475), .ZN(n1152) );
XNOR2_X1 U828 ( .A(G104), .B(n1153), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1132), .A2(n1154), .ZN(G57) );
XNOR2_X1 U830 ( .A(n1155), .B(n1156), .ZN(n1154) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1155) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1136), .ZN(n1158) );
INV_X1 U833 ( .A(G472), .ZN(n1159) );
NAND2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
INV_X1 U835 ( .A(n1162), .ZN(n1161) );
XOR2_X1 U836 ( .A(KEYINPUT59), .B(n1163), .Z(n1160) );
NOR2_X1 U837 ( .A1(n1132), .A2(n1164), .ZN(G54) );
XOR2_X1 U838 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U839 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U840 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U841 ( .A1(KEYINPUT32), .A2(n1171), .ZN(n1170) );
NAND3_X1 U842 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1169) );
OR2_X1 U843 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND3_X1 U844 ( .A1(n1175), .A2(n1176), .A3(KEYINPUT1), .ZN(n1173) );
NOR2_X1 U845 ( .A1(KEYINPUT16), .A2(n1177), .ZN(n1175) );
INV_X1 U846 ( .A(n1178), .ZN(n1177) );
OR2_X1 U847 ( .A1(n1178), .A2(KEYINPUT1), .ZN(n1172) );
XOR2_X1 U848 ( .A(n1179), .B(n1180), .Z(n1165) );
XNOR2_X1 U849 ( .A(KEYINPUT27), .B(n1101), .ZN(n1180) );
NOR2_X1 U850 ( .A1(n1181), .A2(n1136), .ZN(n1179) );
INV_X1 U851 ( .A(G469), .ZN(n1181) );
NOR2_X1 U852 ( .A1(n1132), .A2(n1182), .ZN(G51) );
XOR2_X1 U853 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U854 ( .A(G125), .B(n1185), .Z(n1184) );
NOR2_X1 U855 ( .A1(KEYINPUT50), .A2(n1186), .ZN(n1185) );
XOR2_X1 U856 ( .A(n1187), .B(n1188), .Z(n1183) );
NOR2_X1 U857 ( .A1(n1189), .A2(KEYINPUT8), .ZN(n1188) );
NOR2_X1 U858 ( .A1(n1190), .A2(n1136), .ZN(n1189) );
NAND2_X1 U859 ( .A1(G902), .A2(n1032), .ZN(n1136) );
NAND3_X1 U860 ( .A1(n1112), .A2(n1110), .A3(n1131), .ZN(n1032) );
AND4_X1 U861 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1131) );
AND4_X1 U862 ( .A1(n1153), .A2(n1028), .A3(n1195), .A4(n1196), .ZN(n1194) );
OR3_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1195) );
INV_X1 U864 ( .A(n1200), .ZN(n1198) );
XOR2_X1 U865 ( .A(n1054), .B(KEYINPUT21), .Z(n1197) );
NAND3_X1 U866 ( .A1(n1063), .A2(n1201), .A3(n1049), .ZN(n1028) );
NAND3_X1 U867 ( .A1(n1063), .A2(n1201), .A3(n1050), .ZN(n1153) );
NOR2_X1 U868 ( .A1(n1202), .A2(n1203), .ZN(n1193) );
AND4_X1 U869 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1110) );
NAND2_X1 U870 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
AND4_X1 U871 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1112) );
NOR2_X1 U872 ( .A1(n1097), .A2(G952), .ZN(n1132) );
XNOR2_X1 U873 ( .A(G146), .B(n1210), .ZN(G48) );
NAND3_X1 U874 ( .A1(n1050), .A2(n1054), .A3(n1214), .ZN(n1210) );
XOR2_X1 U875 ( .A(n1215), .B(n1211), .Z(G45) );
NAND4_X1 U876 ( .A1(n1216), .A2(n1065), .A3(n1059), .A4(n1217), .ZN(n1211) );
AND3_X1 U877 ( .A1(n1054), .A2(n1209), .A3(n1218), .ZN(n1217) );
XOR2_X1 U878 ( .A(n1107), .B(n1212), .Z(G42) );
NAND2_X1 U879 ( .A1(n1219), .A2(n1220), .ZN(n1212) );
XOR2_X1 U880 ( .A(G137), .B(n1221), .Z(G39) );
NOR2_X1 U881 ( .A1(KEYINPUT55), .A2(n1213), .ZN(n1221) );
NAND3_X1 U882 ( .A1(n1222), .A2(n1223), .A3(n1214), .ZN(n1213) );
NAND3_X1 U883 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(G36) );
NAND2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U885 ( .A1(n1229), .A2(KEYINPUT53), .ZN(n1228) );
XNOR2_X1 U886 ( .A(G134), .B(KEYINPUT35), .ZN(n1229) );
INV_X1 U887 ( .A(n1205), .ZN(n1227) );
NAND3_X1 U888 ( .A1(KEYINPUT53), .A2(n1205), .A3(G134), .ZN(n1225) );
NAND3_X1 U889 ( .A1(n1059), .A2(n1049), .A3(n1219), .ZN(n1205) );
OR2_X1 U890 ( .A1(G134), .A2(KEYINPUT53), .ZN(n1224) );
XNOR2_X1 U891 ( .A(G131), .B(n1206), .ZN(G33) );
NAND3_X1 U892 ( .A1(n1050), .A2(n1059), .A3(n1219), .ZN(n1206) );
AND3_X1 U893 ( .A1(n1223), .A2(n1209), .A3(n1065), .ZN(n1219) );
XNOR2_X1 U894 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U895 ( .A1(n1049), .A2(n1054), .A3(n1214), .ZN(n1207) );
AND4_X1 U896 ( .A1(n1230), .A2(n1065), .A3(n1060), .A4(n1209), .ZN(n1214) );
XOR2_X1 U897 ( .A(n1231), .B(n1232), .Z(G3) );
NAND2_X1 U898 ( .A1(KEYINPUT14), .A2(n1203), .ZN(n1232) );
AND3_X1 U899 ( .A1(n1222), .A2(n1201), .A3(n1059), .ZN(n1203) );
NAND2_X1 U900 ( .A1(n1233), .A2(n1234), .ZN(G27) );
NAND2_X1 U901 ( .A1(G125), .A2(n1235), .ZN(n1234) );
XOR2_X1 U902 ( .A(n1236), .B(KEYINPUT45), .Z(n1233) );
OR2_X1 U903 ( .A1(n1235), .A2(G125), .ZN(n1236) );
NAND2_X1 U904 ( .A1(n1208), .A2(n1237), .ZN(n1235) );
XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n1209), .ZN(n1237) );
NAND2_X1 U906 ( .A1(n1036), .A2(n1238), .ZN(n1209) );
NAND3_X1 U907 ( .A1(G902), .A2(n1239), .A3(n1115), .ZN(n1238) );
NOR2_X1 U908 ( .A1(G900), .A2(n1097), .ZN(n1115) );
AND3_X1 U909 ( .A1(n1069), .A2(n1054), .A3(n1220), .ZN(n1208) );
AND3_X1 U910 ( .A1(n1061), .A2(n1060), .A3(n1050), .ZN(n1220) );
XOR2_X1 U911 ( .A(G122), .B(n1240), .Z(G24) );
NOR3_X1 U912 ( .A1(n1199), .A2(KEYINPUT34), .A3(n1241), .ZN(n1240) );
NAND4_X1 U913 ( .A1(n1069), .A2(n1063), .A3(n1216), .A4(n1218), .ZN(n1199) );
NOR2_X1 U914 ( .A1(n1060), .A2(n1230), .ZN(n1063) );
XOR2_X1 U915 ( .A(n1242), .B(n1196), .Z(G21) );
NAND4_X1 U916 ( .A1(n1243), .A2(n1060), .A3(n1069), .A4(n1244), .ZN(n1196) );
NOR2_X1 U917 ( .A1(n1052), .A2(n1061), .ZN(n1244) );
INV_X1 U918 ( .A(n1222), .ZN(n1052) );
XOR2_X1 U919 ( .A(G116), .B(n1202), .Z(G18) );
AND2_X1 U920 ( .A1(n1245), .A2(n1049), .ZN(n1202) );
AND2_X1 U921 ( .A1(n1079), .A2(n1216), .ZN(n1049) );
XNOR2_X1 U922 ( .A(n1191), .B(n1246), .ZN(G15) );
NOR2_X1 U923 ( .A1(KEYINPUT57), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U924 ( .A(G113), .B(KEYINPUT15), .ZN(n1247) );
NAND2_X1 U925 ( .A1(n1050), .A2(n1245), .ZN(n1191) );
AND3_X1 U926 ( .A1(n1069), .A2(n1243), .A3(n1059), .ZN(n1245) );
NOR2_X1 U927 ( .A1(n1061), .A2(n1060), .ZN(n1059) );
INV_X1 U928 ( .A(n1040), .ZN(n1069) );
NAND2_X1 U929 ( .A1(n1248), .A2(n1067), .ZN(n1040) );
INV_X1 U930 ( .A(n1066), .ZN(n1248) );
NOR2_X1 U931 ( .A1(n1216), .A2(n1079), .ZN(n1050) );
NAND2_X1 U932 ( .A1(n1249), .A2(n1250), .ZN(G12) );
NAND2_X1 U933 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U934 ( .A(KEYINPUT9), .B(n1253), .Z(n1249) );
NOR2_X1 U935 ( .A1(n1251), .A2(n1252), .ZN(n1253) );
INV_X1 U936 ( .A(n1192), .ZN(n1251) );
NAND4_X1 U937 ( .A1(n1222), .A2(n1201), .A3(n1061), .A4(n1060), .ZN(n1192) );
XNOR2_X1 U938 ( .A(n1084), .B(n1254), .ZN(n1060) );
NOR2_X1 U939 ( .A1(KEYINPUT29), .A2(n1085), .ZN(n1254) );
NAND2_X1 U940 ( .A1(n1134), .A2(n1255), .ZN(n1085) );
XNOR2_X1 U941 ( .A(n1256), .B(n1257), .ZN(n1134) );
XNOR2_X1 U942 ( .A(n1258), .B(n1259), .ZN(n1257) );
XOR2_X1 U943 ( .A(n1260), .B(n1261), .Z(n1259) );
NAND2_X1 U944 ( .A1(KEYINPUT0), .A2(n1262), .ZN(n1260) );
NAND2_X1 U945 ( .A1(G221), .A2(n1263), .ZN(n1262) );
XOR2_X1 U946 ( .A(n1264), .B(n1265), .Z(n1256) );
NOR2_X1 U947 ( .A1(KEYINPUT39), .A2(n1266), .ZN(n1265) );
XOR2_X1 U948 ( .A(n1252), .B(n1267), .Z(n1266) );
XOR2_X1 U949 ( .A(G128), .B(G119), .Z(n1267) );
XOR2_X1 U950 ( .A(n1107), .B(G125), .Z(n1264) );
INV_X1 U951 ( .A(G140), .ZN(n1107) );
NAND2_X1 U952 ( .A1(G217), .A2(n1268), .ZN(n1084) );
INV_X1 U953 ( .A(n1230), .ZN(n1061) );
XOR2_X1 U954 ( .A(n1086), .B(n1269), .Z(n1230) );
NOR2_X1 U955 ( .A1(G472), .A2(KEYINPUT63), .ZN(n1269) );
NAND2_X1 U956 ( .A1(n1270), .A2(n1255), .ZN(n1086) );
XOR2_X1 U957 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U958 ( .A1(n1163), .A2(n1162), .ZN(n1272) );
NOR2_X1 U959 ( .A1(n1231), .A2(n1273), .ZN(n1162) );
AND2_X1 U960 ( .A1(n1231), .A2(n1273), .ZN(n1163) );
NAND3_X1 U961 ( .A1(n1274), .A2(n1275), .A3(G210), .ZN(n1273) );
XOR2_X1 U962 ( .A(KEYINPUT12), .B(G953), .Z(n1274) );
NOR2_X1 U963 ( .A1(KEYINPUT51), .A2(n1156), .ZN(n1271) );
XOR2_X1 U964 ( .A(n1276), .B(n1277), .Z(n1156) );
XOR2_X1 U965 ( .A(n1167), .B(n1278), .Z(n1277) );
XOR2_X1 U966 ( .A(G113), .B(n1279), .Z(n1278) );
INV_X1 U967 ( .A(n1280), .ZN(n1167) );
XNOR2_X1 U968 ( .A(G116), .B(n1281), .ZN(n1276) );
XOR2_X1 U969 ( .A(KEYINPUT5), .B(G119), .Z(n1281) );
AND2_X1 U970 ( .A1(n1065), .A2(n1243), .ZN(n1201) );
INV_X1 U971 ( .A(n1241), .ZN(n1243) );
NAND2_X1 U972 ( .A1(n1054), .A2(n1200), .ZN(n1241) );
NAND2_X1 U973 ( .A1(n1036), .A2(n1282), .ZN(n1200) );
NAND3_X1 U974 ( .A1(n1283), .A2(n1239), .A3(G902), .ZN(n1282) );
INV_X1 U975 ( .A(n1122), .ZN(n1283) );
NAND2_X1 U976 ( .A1(G953), .A2(n1284), .ZN(n1122) );
XOR2_X1 U977 ( .A(KEYINPUT11), .B(G898), .Z(n1284) );
NAND3_X1 U978 ( .A1(n1239), .A2(n1097), .A3(G952), .ZN(n1036) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1239) );
NAND2_X1 U980 ( .A1(n1285), .A2(n1286), .ZN(n1054) );
OR2_X1 U981 ( .A1(n1048), .A2(KEYINPUT4), .ZN(n1286) );
INV_X1 U982 ( .A(n1223), .ZN(n1048) );
NOR2_X1 U983 ( .A1(n1055), .A2(n1073), .ZN(n1223) );
INV_X1 U984 ( .A(n1056), .ZN(n1073) );
NAND3_X1 U985 ( .A1(n1056), .A2(n1055), .A3(KEYINPUT4), .ZN(n1285) );
OR2_X1 U986 ( .A1(n1072), .A2(n1074), .ZN(n1055) );
AND3_X1 U987 ( .A1(n1190), .A2(n1255), .A3(n1287), .ZN(n1074) );
NOR2_X1 U988 ( .A1(n1190), .A2(n1288), .ZN(n1072) );
AND2_X1 U989 ( .A1(n1287), .A2(n1255), .ZN(n1288) );
XOR2_X1 U990 ( .A(n1289), .B(n1290), .Z(n1287) );
XOR2_X1 U991 ( .A(n1291), .B(n1187), .Z(n1290) );
XOR2_X1 U992 ( .A(n1292), .B(n1279), .Z(n1187) );
XNOR2_X1 U993 ( .A(n1293), .B(n1294), .ZN(n1279) );
NOR3_X1 U994 ( .A1(KEYINPUT56), .A2(n1295), .A3(n1296), .ZN(n1294) );
NOR2_X1 U995 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
INV_X1 U996 ( .A(KEYINPUT10), .ZN(n1297) );
NOR2_X1 U997 ( .A1(KEYINPUT10), .A2(n1299), .ZN(n1295) );
XNOR2_X1 U998 ( .A(G128), .B(KEYINPUT47), .ZN(n1293) );
NAND2_X1 U999 ( .A1(G224), .A2(n1097), .ZN(n1292) );
NAND2_X1 U1000 ( .A1(KEYINPUT3), .A2(G125), .ZN(n1291) );
XNOR2_X1 U1001 ( .A(KEYINPUT58), .B(n1300), .ZN(n1289) );
NOR2_X1 U1002 ( .A1(KEYINPUT52), .A2(n1186), .ZN(n1300) );
XNOR2_X1 U1003 ( .A(n1301), .B(n1127), .ZN(n1186) );
XOR2_X1 U1004 ( .A(n1129), .B(n1130), .Z(n1127) );
AND2_X1 U1005 ( .A1(n1302), .A2(n1303), .ZN(n1130) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1242), .ZN(n1303) );
INV_X1 U1007 ( .A(G119), .ZN(n1242) );
XOR2_X1 U1008 ( .A(KEYINPUT30), .B(n1305), .Z(n1304) );
NAND2_X1 U1009 ( .A1(n1305), .A2(G119), .ZN(n1302) );
XOR2_X1 U1010 ( .A(G113), .B(G116), .Z(n1305) );
XNOR2_X1 U1011 ( .A(n1306), .B(n1307), .ZN(n1129) );
NOR2_X1 U1012 ( .A1(KEYINPUT42), .A2(n1027), .ZN(n1307) );
XOR2_X1 U1013 ( .A(n1124), .B(KEYINPUT24), .Z(n1301) );
XOR2_X1 U1014 ( .A(n1252), .B(G122), .Z(n1124) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1308), .ZN(n1190) );
NAND2_X1 U1016 ( .A1(G214), .A2(n1308), .ZN(n1056) );
NAND2_X1 U1017 ( .A1(n1275), .A2(n1255), .ZN(n1308) );
AND2_X1 U1018 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1268), .ZN(n1067) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1255), .ZN(n1268) );
XNOR2_X1 U1021 ( .A(n1309), .B(G469), .ZN(n1066) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1255), .ZN(n1309) );
XOR2_X1 U1023 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U1024 ( .A(n1313), .B(n1171), .ZN(n1312) );
XNOR2_X1 U1025 ( .A(n1314), .B(n1306), .ZN(n1171) );
XOR2_X1 U1026 ( .A(n1231), .B(n1315), .Z(n1306) );
XOR2_X1 U1027 ( .A(KEYINPUT49), .B(G104), .Z(n1315) );
INV_X1 U1028 ( .A(G101), .ZN(n1231) );
NAND2_X1 U1029 ( .A1(KEYINPUT7), .A2(n1027), .ZN(n1314) );
XOR2_X1 U1030 ( .A(n1280), .B(n1178), .Z(n1313) );
XNOR2_X1 U1031 ( .A(n1252), .B(G140), .ZN(n1178) );
INV_X1 U1032 ( .A(G110), .ZN(n1252) );
XNOR2_X1 U1033 ( .A(n1102), .B(n1316), .ZN(n1280) );
XOR2_X1 U1034 ( .A(KEYINPUT38), .B(G131), .Z(n1316) );
XOR2_X1 U1035 ( .A(G134), .B(n1258), .Z(n1102) );
XOR2_X1 U1036 ( .A(G137), .B(KEYINPUT62), .Z(n1258) );
XNOR2_X1 U1037 ( .A(n1317), .B(n1101), .ZN(n1311) );
NAND2_X1 U1038 ( .A1(n1318), .A2(n1319), .ZN(n1101) );
NAND2_X1 U1039 ( .A1(G128), .A2(n1320), .ZN(n1319) );
XOR2_X1 U1040 ( .A(n1321), .B(KEYINPUT43), .Z(n1318) );
OR2_X1 U1041 ( .A1(n1320), .A2(G128), .ZN(n1321) );
NAND3_X1 U1042 ( .A1(n1322), .A2(n1323), .A3(n1298), .ZN(n1320) );
OR3_X1 U1043 ( .A1(n1215), .A2(n1324), .A3(KEYINPUT46), .ZN(n1323) );
NAND2_X1 U1044 ( .A1(KEYINPUT46), .A2(n1215), .ZN(n1322) );
XNOR2_X1 U1045 ( .A(n1176), .B(KEYINPUT6), .ZN(n1317) );
NOR2_X1 U1046 ( .A1(n1114), .A2(G953), .ZN(n1176) );
INV_X1 U1047 ( .A(G227), .ZN(n1114) );
NOR2_X1 U1048 ( .A1(n1218), .A2(n1216), .ZN(n1222) );
XOR2_X1 U1049 ( .A(n1083), .B(n1325), .Z(n1216) );
NOR2_X1 U1050 ( .A1(G478), .A2(KEYINPUT28), .ZN(n1325) );
NAND2_X1 U1051 ( .A1(n1144), .A2(n1255), .ZN(n1083) );
INV_X1 U1052 ( .A(G902), .ZN(n1255) );
NAND2_X1 U1053 ( .A1(n1326), .A2(n1327), .ZN(n1144) );
NAND3_X1 U1054 ( .A1(G217), .A2(n1263), .A3(n1328), .ZN(n1327) );
XOR2_X1 U1055 ( .A(n1329), .B(KEYINPUT31), .Z(n1328) );
XOR2_X1 U1056 ( .A(n1330), .B(KEYINPUT18), .Z(n1326) );
NAND2_X1 U1057 ( .A1(n1329), .A2(n1331), .ZN(n1330) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1263), .ZN(n1331) );
AND2_X1 U1059 ( .A1(G234), .A2(n1097), .ZN(n1263) );
XOR2_X1 U1060 ( .A(n1332), .B(n1333), .Z(n1329) );
XOR2_X1 U1061 ( .A(n1334), .B(n1335), .Z(n1333) );
NAND2_X1 U1062 ( .A1(KEYINPUT22), .A2(n1336), .ZN(n1335) );
INV_X1 U1063 ( .A(G122), .ZN(n1336) );
NAND2_X1 U1064 ( .A1(n1337), .A2(n1338), .ZN(n1334) );
NAND2_X1 U1065 ( .A1(n1339), .A2(G134), .ZN(n1338) );
XOR2_X1 U1066 ( .A(KEYINPUT26), .B(n1340), .Z(n1337) );
NOR2_X1 U1067 ( .A1(G134), .A2(n1339), .ZN(n1340) );
XNOR2_X1 U1068 ( .A(G128), .B(n1341), .ZN(n1339) );
NOR2_X1 U1069 ( .A1(KEYINPUT41), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1070 ( .A(KEYINPUT40), .B(G143), .Z(n1342) );
XOR2_X1 U1071 ( .A(n1027), .B(G116), .Z(n1332) );
INV_X1 U1072 ( .A(G107), .ZN(n1027) );
INV_X1 U1073 ( .A(n1079), .ZN(n1218) );
XOR2_X1 U1074 ( .A(n1343), .B(G475), .Z(n1079) );
OR2_X1 U1075 ( .A1(n1151), .A2(G902), .ZN(n1343) );
XNOR2_X1 U1076 ( .A(n1299), .B(n1344), .ZN(n1151) );
XOR2_X1 U1077 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1078 ( .A(n1347), .B(n1348), .Z(n1346) );
XOR2_X1 U1079 ( .A(G104), .B(n1349), .Z(n1348) );
AND3_X1 U1080 ( .A1(G214), .A2(n1097), .A3(n1275), .ZN(n1349) );
INV_X1 U1081 ( .A(G237), .ZN(n1275) );
INV_X1 U1082 ( .A(G953), .ZN(n1097) );
XOR2_X1 U1083 ( .A(G122), .B(G113), .Z(n1347) );
XOR2_X1 U1084 ( .A(n1350), .B(n1351), .Z(n1345) );
XOR2_X1 U1085 ( .A(G131), .B(G125), .Z(n1351) );
XOR2_X1 U1086 ( .A(KEYINPUT44), .B(G140), .Z(n1350) );
NAND2_X1 U1087 ( .A1(n1298), .A2(n1352), .ZN(n1299) );
NAND2_X1 U1088 ( .A1(G143), .A2(n1261), .ZN(n1352) );
INV_X1 U1089 ( .A(n1324), .ZN(n1261) );
NAND2_X1 U1090 ( .A1(n1324), .A2(n1215), .ZN(n1298) );
INV_X1 U1091 ( .A(G143), .ZN(n1215) );
XNOR2_X1 U1092 ( .A(G146), .B(KEYINPUT33), .ZN(n1324) );
endmodule


