//Key = 0110010100110011010110000000010100001100000111000111111011010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;

XOR2_X1 U749 ( .A(n1036), .B(n1037), .Z(G9) );
NAND2_X1 U750 ( .A1(KEYINPUT11), .A2(G107), .ZN(n1037) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR4_X1 U752 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
XOR2_X1 U753 ( .A(n1044), .B(KEYINPUT51), .Z(n1042) );
NAND4_X1 U754 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044) );
NAND4_X1 U755 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1040) );
NAND4_X1 U756 ( .A1(n1045), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1046), .A2(n1058), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1063), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U769 ( .A(n1078), .ZN(n1045) );
NAND2_X1 U770 ( .A1(n1047), .A2(n1079), .ZN(n1049) );
XOR2_X1 U771 ( .A(KEYINPUT30), .B(n1080), .Z(n1079) );
NOR3_X1 U772 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
INV_X1 U773 ( .A(n1084), .ZN(n1082) );
XNOR2_X1 U774 ( .A(KEYINPUT37), .B(n1078), .ZN(n1081) );
NOR3_X1 U775 ( .A1(n1085), .A2(G953), .A3(G952), .ZN(n1038) );
INV_X1 U776 ( .A(n1051), .ZN(n1085) );
NAND4_X1 U777 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1051) );
NOR4_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
XNOR2_X1 U779 ( .A(G472), .B(n1094), .ZN(n1093) );
XOR2_X1 U780 ( .A(n1095), .B(n1096), .Z(n1091) );
NOR2_X1 U781 ( .A1(KEYINPUT18), .A2(n1097), .ZN(n1096) );
XOR2_X1 U782 ( .A(n1098), .B(KEYINPUT2), .Z(n1097) );
XOR2_X1 U783 ( .A(n1099), .B(n1100), .Z(n1090) );
NAND2_X1 U784 ( .A1(KEYINPUT53), .A2(n1101), .ZN(n1099) );
NOR3_X1 U785 ( .A1(n1061), .A2(n1102), .A3(n1103), .ZN(n1088) );
INV_X1 U786 ( .A(n1104), .ZN(n1103) );
OR2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1086) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(G72) );
NOR2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U790 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U791 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U792 ( .A(n1115), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1115), .ZN(n1109) );
NAND3_X1 U794 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
XOR2_X1 U795 ( .A(KEYINPUT62), .B(n1119), .Z(n1118) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XNOR2_X1 U798 ( .A(n1122), .B(G140), .ZN(n1121) );
NAND2_X1 U799 ( .A1(KEYINPUT54), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U800 ( .A(n1124), .B(n1125), .ZN(n1120) );
XNOR2_X1 U801 ( .A(n1126), .B(n1127), .ZN(n1125) );
XNOR2_X1 U802 ( .A(KEYINPUT16), .B(n1128), .ZN(n1127) );
XNOR2_X1 U803 ( .A(n1129), .B(G131), .ZN(n1124) );
INV_X1 U804 ( .A(n1114), .ZN(n1116) );
NOR2_X1 U805 ( .A1(G227), .A2(n1052), .ZN(n1113) );
NAND2_X1 U806 ( .A1(n1052), .A2(n1041), .ZN(n1107) );
NAND2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(G69) );
NAND2_X1 U808 ( .A1(n1132), .A2(n1052), .ZN(n1131) );
XNOR2_X1 U809 ( .A(n1133), .B(n1043), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1134), .A2(G953), .ZN(n1130) );
NAND2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1133), .A2(n1137), .ZN(n1136) );
INV_X1 U813 ( .A(G224), .ZN(n1137) );
NAND2_X1 U814 ( .A1(G224), .A2(n1138), .ZN(n1135) );
NAND2_X1 U815 ( .A1(G898), .A2(n1133), .ZN(n1138) );
NAND2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1133) );
NAND2_X1 U817 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1139) );
XNOR2_X1 U819 ( .A(KEYINPUT58), .B(n1144), .ZN(n1143) );
NOR2_X1 U820 ( .A1(KEYINPUT47), .A2(n1145), .ZN(n1144) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U823 ( .A1(n1105), .A2(n1150), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1146), .A2(n1151), .ZN(G63) );
XNOR2_X1 U825 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR3_X1 U826 ( .A1(n1150), .A2(KEYINPUT6), .A3(n1154), .ZN(n1153) );
INV_X1 U827 ( .A(G478), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1146), .A2(n1155), .ZN(G60) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U830 ( .A1(KEYINPUT21), .A2(n1158), .ZN(n1157) );
OR2_X1 U831 ( .A1(n1150), .A2(n1101), .ZN(n1156) );
XOR2_X1 U832 ( .A(G104), .B(n1159), .Z(G6) );
NOR2_X1 U833 ( .A1(n1160), .A2(n1059), .ZN(n1159) );
XOR2_X1 U834 ( .A(n1161), .B(KEYINPUT23), .Z(n1160) );
NOR2_X1 U835 ( .A1(n1146), .A2(n1162), .ZN(G57) );
XOR2_X1 U836 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U838 ( .A1(n1167), .A2(n1150), .ZN(n1166) );
INV_X1 U839 ( .A(G472), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1168), .A2(KEYINPUT14), .ZN(n1165) );
XNOR2_X1 U841 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U842 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U843 ( .A1(n1173), .A2(KEYINPUT38), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1146), .A2(n1174), .ZN(G54) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U846 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U847 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1150), .ZN(n1180) );
NOR3_X1 U849 ( .A1(n1182), .A2(KEYINPUT13), .A3(n1183), .ZN(n1177) );
INV_X1 U850 ( .A(G227), .ZN(n1182) );
XOR2_X1 U851 ( .A(n1184), .B(n1185), .Z(n1175) );
NOR2_X1 U852 ( .A1(n1146), .A2(n1186), .ZN(G51) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U854 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NAND2_X1 U856 ( .A1(G125), .A2(n1193), .ZN(n1192) );
XOR2_X1 U857 ( .A(KEYINPUT1), .B(n1194), .Z(n1191) );
NOR2_X1 U858 ( .A1(G125), .A2(n1193), .ZN(n1194) );
XOR2_X1 U859 ( .A(n1195), .B(n1196), .Z(n1187) );
NOR2_X1 U860 ( .A1(n1095), .A2(n1150), .ZN(n1196) );
NAND2_X1 U861 ( .A1(G902), .A2(n1197), .ZN(n1150) );
OR2_X1 U862 ( .A1(n1041), .A2(n1043), .ZN(n1197) );
NAND4_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1043) );
AND4_X1 U864 ( .A1(n1202), .A2(n1036), .A3(n1203), .A4(n1204), .ZN(n1201) );
NAND3_X1 U865 ( .A1(n1048), .A2(n1205), .A3(n1206), .ZN(n1036) );
NOR3_X1 U866 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
AND4_X1 U868 ( .A1(n1210), .A2(n1212), .A3(n1068), .A4(n1213), .ZN(n1208) );
INV_X1 U869 ( .A(n1214), .ZN(n1068) );
INV_X1 U870 ( .A(KEYINPUT10), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1059), .A2(n1161), .ZN(n1207) );
NAND2_X1 U872 ( .A1(n1084), .A2(n1205), .ZN(n1161) );
AND3_X1 U873 ( .A1(n1066), .A2(n1215), .A3(n1214), .ZN(n1205) );
NAND4_X1 U874 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1041) );
NOR4_X1 U875 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
INV_X1 U876 ( .A(n1224), .ZN(n1223) );
NOR2_X1 U877 ( .A1(n1225), .A2(n1226), .ZN(n1218) );
AND3_X1 U878 ( .A1(n1047), .A2(n1214), .A3(n1227), .ZN(n1226) );
NOR2_X1 U879 ( .A1(n1052), .A2(G952), .ZN(n1146) );
XOR2_X1 U880 ( .A(n1225), .B(n1228), .Z(G48) );
NOR2_X1 U881 ( .A1(KEYINPUT33), .A2(n1229), .ZN(n1228) );
AND3_X1 U882 ( .A1(n1230), .A2(n1206), .A3(n1084), .ZN(n1225) );
XNOR2_X1 U883 ( .A(G143), .B(n1216), .ZN(G45) );
NAND4_X1 U884 ( .A1(n1231), .A2(n1206), .A3(n1232), .A4(n1233), .ZN(n1216) );
XNOR2_X1 U885 ( .A(G140), .B(n1234), .ZN(G42) );
NAND4_X1 U886 ( .A1(KEYINPUT5), .A2(n1047), .A3(n1227), .A4(n1214), .ZN(n1234) );
INV_X1 U887 ( .A(n1235), .ZN(n1227) );
XNOR2_X1 U888 ( .A(G137), .B(n1217), .ZN(G39) );
NAND4_X1 U889 ( .A1(n1047), .A2(n1053), .A3(n1054), .A4(n1230), .ZN(n1217) );
XNOR2_X1 U890 ( .A(G134), .B(n1224), .ZN(G36) );
NAND3_X1 U891 ( .A1(n1231), .A2(n1048), .A3(n1047), .ZN(n1224) );
XOR2_X1 U892 ( .A(G131), .B(n1222), .Z(G33) );
AND3_X1 U893 ( .A1(n1231), .A2(n1084), .A3(n1047), .ZN(n1222) );
NOR2_X1 U894 ( .A1(n1236), .A2(n1061), .ZN(n1047) );
AND3_X1 U895 ( .A1(n1214), .A2(n1237), .A3(n1213), .ZN(n1231) );
XNOR2_X1 U896 ( .A(n1238), .B(n1220), .ZN(G30) );
AND3_X1 U897 ( .A1(n1206), .A2(n1048), .A3(n1230), .ZN(n1220) );
AND4_X1 U898 ( .A1(n1239), .A2(n1214), .A3(n1237), .A4(n1077), .ZN(n1230) );
XNOR2_X1 U899 ( .A(n1240), .B(n1211), .ZN(G3) );
NAND3_X1 U900 ( .A1(n1213), .A2(n1214), .A3(n1212), .ZN(n1211) );
NAND2_X1 U901 ( .A1(KEYINPUT50), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U902 ( .A(n1123), .B(n1221), .ZN(G27) );
NOR3_X1 U903 ( .A1(n1092), .A2(n1059), .A3(n1235), .ZN(n1221) );
NAND4_X1 U904 ( .A1(n1084), .A2(n1076), .A3(n1237), .A4(n1077), .ZN(n1235) );
NAND2_X1 U905 ( .A1(n1078), .A2(n1242), .ZN(n1237) );
NAND3_X1 U906 ( .A1(G902), .A2(n1243), .A3(n1114), .ZN(n1242) );
NOR2_X1 U907 ( .A1(G900), .A2(n1052), .ZN(n1114) );
INV_X1 U908 ( .A(G125), .ZN(n1123) );
XNOR2_X1 U909 ( .A(G122), .B(n1202), .ZN(G24) );
NAND3_X1 U910 ( .A1(n1046), .A2(n1206), .A3(n1244), .ZN(n1202) );
NOR3_X1 U911 ( .A1(n1054), .A2(n1053), .A3(n1245), .ZN(n1244) );
INV_X1 U912 ( .A(n1083), .ZN(n1046) );
NAND2_X1 U913 ( .A1(n1072), .A2(n1066), .ZN(n1083) );
NOR2_X1 U914 ( .A1(n1077), .A2(n1239), .ZN(n1066) );
XNOR2_X1 U915 ( .A(G119), .B(n1198), .ZN(G21) );
NAND4_X1 U916 ( .A1(n1239), .A2(n1212), .A3(n1072), .A4(n1077), .ZN(n1198) );
INV_X1 U917 ( .A(n1092), .ZN(n1072) );
INV_X1 U918 ( .A(n1076), .ZN(n1239) );
XNOR2_X1 U919 ( .A(G116), .B(n1199), .ZN(G18) );
NAND2_X1 U920 ( .A1(n1246), .A2(n1048), .ZN(n1199) );
NOR2_X1 U921 ( .A1(n1232), .A2(n1053), .ZN(n1048) );
INV_X1 U922 ( .A(n1233), .ZN(n1053) );
XNOR2_X1 U923 ( .A(G113), .B(n1204), .ZN(G15) );
NAND2_X1 U924 ( .A1(n1246), .A2(n1084), .ZN(n1204) );
NOR2_X1 U925 ( .A1(n1233), .A2(n1054), .ZN(n1084) );
NOR4_X1 U926 ( .A1(n1074), .A2(n1092), .A3(n1059), .A4(n1245), .ZN(n1246) );
NAND2_X1 U927 ( .A1(n1071), .A2(n1247), .ZN(n1092) );
INV_X1 U928 ( .A(n1213), .ZN(n1074) );
NOR2_X1 U929 ( .A1(n1076), .A2(n1077), .ZN(n1213) );
XNOR2_X1 U930 ( .A(n1248), .B(n1249), .ZN(G12) );
NOR2_X1 U931 ( .A1(KEYINPUT25), .A2(n1203), .ZN(n1249) );
NAND4_X1 U932 ( .A1(n1212), .A2(n1214), .A3(n1076), .A4(n1077), .ZN(n1203) );
NAND3_X1 U933 ( .A1(n1250), .A2(n1251), .A3(n1104), .ZN(n1077) );
NAND2_X1 U934 ( .A1(n1106), .A2(n1105), .ZN(n1104) );
OR3_X1 U935 ( .A1(n1105), .A2(n1106), .A3(KEYINPUT28), .ZN(n1251) );
NOR2_X1 U936 ( .A1(n1252), .A2(n1149), .ZN(n1106) );
XNOR2_X1 U937 ( .A(n1253), .B(n1254), .ZN(n1149) );
NOR2_X1 U938 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NOR2_X1 U939 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U940 ( .A(G137), .B(KEYINPUT40), .ZN(n1258) );
AND2_X1 U941 ( .A1(n1128), .A2(n1257), .ZN(n1255) );
NAND3_X1 U942 ( .A1(n1259), .A2(G234), .A3(G221), .ZN(n1257) );
NAND2_X1 U943 ( .A1(n1260), .A2(n1261), .ZN(n1253) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U945 ( .A(KEYINPUT20), .B(n1264), .ZN(n1263) );
XOR2_X1 U946 ( .A(KEYINPUT59), .B(n1265), .Z(n1260) );
NOR2_X1 U947 ( .A1(n1262), .A2(n1264), .ZN(n1265) );
XOR2_X1 U948 ( .A(n1266), .B(n1267), .Z(n1264) );
XNOR2_X1 U949 ( .A(KEYINPUT39), .B(n1268), .ZN(n1267) );
XNOR2_X1 U950 ( .A(n1269), .B(n1248), .ZN(n1266) );
NAND2_X1 U951 ( .A1(KEYINPUT49), .A2(G128), .ZN(n1269) );
XOR2_X1 U952 ( .A(n1270), .B(n1271), .Z(n1262) );
NOR2_X1 U953 ( .A1(G146), .A2(KEYINPUT22), .ZN(n1271) );
XNOR2_X1 U954 ( .A(G125), .B(n1272), .ZN(n1270) );
NOR2_X1 U955 ( .A1(KEYINPUT9), .A2(n1273), .ZN(n1272) );
INV_X1 U956 ( .A(G140), .ZN(n1273) );
NAND2_X1 U957 ( .A1(KEYINPUT28), .A2(n1105), .ZN(n1250) );
NAND2_X1 U958 ( .A1(G217), .A2(n1274), .ZN(n1105) );
XOR2_X1 U959 ( .A(G472), .B(n1275), .Z(n1076) );
NOR2_X1 U960 ( .A1(KEYINPUT3), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U961 ( .A(KEYINPUT63), .B(n1094), .ZN(n1276) );
NAND2_X1 U962 ( .A1(n1277), .A2(n1278), .ZN(n1094) );
XOR2_X1 U963 ( .A(n1279), .B(n1280), .Z(n1277) );
XNOR2_X1 U964 ( .A(n1173), .B(n1281), .ZN(n1280) );
NAND2_X1 U965 ( .A1(KEYINPUT15), .A2(n1172), .ZN(n1281) );
XNOR2_X1 U966 ( .A(n1163), .B(n1282), .ZN(n1279) );
INV_X1 U967 ( .A(n1169), .ZN(n1282) );
XNOR2_X1 U968 ( .A(n1283), .B(G113), .ZN(n1169) );
NAND2_X1 U969 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U970 ( .A1(G116), .A2(n1268), .ZN(n1285) );
XOR2_X1 U971 ( .A(n1286), .B(KEYINPUT34), .Z(n1284) );
NAND2_X1 U972 ( .A1(G119), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U973 ( .A(n1288), .B(n1241), .ZN(n1163) );
INV_X1 U974 ( .A(G101), .ZN(n1241) );
NAND3_X1 U975 ( .A1(n1289), .A2(n1290), .A3(G210), .ZN(n1288) );
XNOR2_X1 U976 ( .A(KEYINPUT17), .B(n1259), .ZN(n1289) );
NOR2_X1 U977 ( .A1(n1071), .A2(n1070), .ZN(n1214) );
INV_X1 U978 ( .A(n1247), .ZN(n1070) );
NAND2_X1 U979 ( .A1(n1291), .A2(n1274), .ZN(n1247) );
NAND2_X1 U980 ( .A1(G234), .A2(n1292), .ZN(n1274) );
XNOR2_X1 U981 ( .A(G221), .B(KEYINPUT57), .ZN(n1291) );
XNOR2_X1 U982 ( .A(n1293), .B(n1181), .ZN(n1071) );
INV_X1 U983 ( .A(G469), .ZN(n1181) );
NAND3_X1 U984 ( .A1(n1294), .A2(n1295), .A3(n1278), .ZN(n1293) );
NAND2_X1 U985 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U986 ( .A1(G227), .A2(n1259), .ZN(n1297) );
XOR2_X1 U987 ( .A(n1298), .B(n1299), .Z(n1296) );
NOR2_X1 U988 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND3_X1 U989 ( .A1(n1259), .A2(G227), .A3(n1302), .ZN(n1294) );
XOR2_X1 U990 ( .A(n1298), .B(n1303), .Z(n1302) );
NOR2_X1 U991 ( .A1(n1304), .A2(n1301), .ZN(n1303) );
INV_X1 U992 ( .A(KEYINPUT45), .ZN(n1301) );
XNOR2_X1 U993 ( .A(n1300), .B(KEYINPUT24), .ZN(n1304) );
XNOR2_X1 U994 ( .A(n1184), .B(KEYINPUT29), .ZN(n1300) );
XNOR2_X1 U995 ( .A(G110), .B(G140), .ZN(n1184) );
XNOR2_X1 U996 ( .A(n1185), .B(n1305), .ZN(n1298) );
XNOR2_X1 U997 ( .A(n1306), .B(KEYINPUT48), .ZN(n1305) );
NAND2_X1 U998 ( .A1(KEYINPUT56), .A2(n1129), .ZN(n1306) );
INV_X1 U999 ( .A(n1179), .ZN(n1129) );
NAND3_X1 U1000 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1179) );
NAND2_X1 U1001 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
INV_X1 U1002 ( .A(KEYINPUT52), .ZN(n1311) );
NAND2_X1 U1003 ( .A1(G128), .A2(n1312), .ZN(n1310) );
XNOR2_X1 U1004 ( .A(KEYINPUT41), .B(n1313), .ZN(n1312) );
NAND2_X1 U1005 ( .A1(KEYINPUT52), .A2(n1314), .ZN(n1307) );
NAND2_X1 U1006 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
OR3_X1 U1007 ( .A1(n1238), .A2(n1313), .A3(KEYINPUT41), .ZN(n1316) );
NAND2_X1 U1008 ( .A1(KEYINPUT41), .A2(n1313), .ZN(n1315) );
XNOR2_X1 U1009 ( .A(n1317), .B(n1172), .ZN(n1185) );
XNOR2_X1 U1010 ( .A(n1318), .B(G131), .ZN(n1172) );
NAND2_X1 U1011 ( .A1(n1319), .A2(KEYINPUT31), .ZN(n1318) );
XOR2_X1 U1012 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1013 ( .A(KEYINPUT4), .B(n1128), .ZN(n1321) );
INV_X1 U1014 ( .A(G137), .ZN(n1128) );
NAND2_X1 U1015 ( .A1(KEYINPUT19), .A2(n1126), .ZN(n1320) );
NOR4_X1 U1016 ( .A1(n1233), .A2(n1059), .A3(n1232), .A4(n1245), .ZN(n1212) );
INV_X1 U1017 ( .A(n1215), .ZN(n1245) );
NAND2_X1 U1018 ( .A1(n1078), .A2(n1322), .ZN(n1215) );
NAND4_X1 U1019 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1141), .ZN(n1322) );
INV_X1 U1020 ( .A(G898), .ZN(n1141) );
NAND3_X1 U1021 ( .A1(n1243), .A2(n1052), .A3(G952), .ZN(n1078) );
INV_X1 U1022 ( .A(G953), .ZN(n1052) );
NAND2_X1 U1023 ( .A1(G237), .A2(G234), .ZN(n1243) );
INV_X1 U1024 ( .A(n1054), .ZN(n1232) );
XOR2_X1 U1025 ( .A(n1100), .B(n1101), .Z(n1054) );
INV_X1 U1026 ( .A(G475), .ZN(n1101) );
NOR2_X1 U1027 ( .A1(n1158), .A2(n1252), .ZN(n1100) );
XNOR2_X1 U1028 ( .A(n1323), .B(n1324), .ZN(n1158) );
XOR2_X1 U1029 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1030 ( .A(n1327), .B(n1328), .ZN(n1326) );
NAND2_X1 U1031 ( .A1(KEYINPUT43), .A2(n1329), .ZN(n1328) );
INV_X1 U1032 ( .A(G143), .ZN(n1329) );
NAND2_X1 U1033 ( .A1(KEYINPUT36), .A2(n1330), .ZN(n1327) );
XOR2_X1 U1034 ( .A(G113), .B(n1331), .Z(n1330) );
XOR2_X1 U1035 ( .A(KEYINPUT26), .B(G122), .Z(n1331) );
XNOR2_X1 U1036 ( .A(G104), .B(n1332), .ZN(n1325) );
AND3_X1 U1037 ( .A1(n1259), .A2(n1290), .A3(G214), .ZN(n1332) );
XOR2_X1 U1038 ( .A(n1333), .B(n1334), .Z(n1323) );
XNOR2_X1 U1039 ( .A(n1229), .B(G140), .ZN(n1334) );
XNOR2_X1 U1040 ( .A(G131), .B(G125), .ZN(n1333) );
INV_X1 U1041 ( .A(n1206), .ZN(n1059) );
NOR2_X1 U1042 ( .A1(n1062), .A2(n1061), .ZN(n1206) );
AND2_X1 U1043 ( .A1(G214), .A2(n1335), .ZN(n1061) );
INV_X1 U1044 ( .A(n1236), .ZN(n1062) );
XOR2_X1 U1045 ( .A(n1098), .B(n1095), .Z(n1236) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1335), .ZN(n1095) );
NAND2_X1 U1047 ( .A1(n1290), .A2(n1292), .ZN(n1335) );
INV_X1 U1048 ( .A(G902), .ZN(n1292) );
INV_X1 U1049 ( .A(G237), .ZN(n1290) );
NAND2_X1 U1050 ( .A1(n1336), .A2(n1278), .ZN(n1098) );
XNOR2_X1 U1051 ( .A(n1337), .B(n1338), .ZN(n1336) );
INV_X1 U1052 ( .A(n1190), .ZN(n1338) );
XNOR2_X1 U1053 ( .A(n1142), .B(n1145), .ZN(n1190) );
XNOR2_X1 U1054 ( .A(n1248), .B(G122), .ZN(n1145) );
XOR2_X1 U1055 ( .A(n1339), .B(n1340), .Z(n1142) );
XNOR2_X1 U1056 ( .A(n1287), .B(n1341), .ZN(n1340) );
XNOR2_X1 U1057 ( .A(KEYINPUT32), .B(n1268), .ZN(n1341) );
INV_X1 U1058 ( .A(G119), .ZN(n1268) );
XOR2_X1 U1059 ( .A(n1317), .B(G113), .Z(n1339) );
XNOR2_X1 U1060 ( .A(G101), .B(n1342), .ZN(n1317) );
XOR2_X1 U1061 ( .A(G107), .B(G104), .Z(n1342) );
XNOR2_X1 U1062 ( .A(KEYINPUT35), .B(n1343), .ZN(n1337) );
NOR2_X1 U1063 ( .A1(KEYINPUT61), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1064 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1065 ( .A(n1173), .B(G125), .ZN(n1346) );
INV_X1 U1066 ( .A(n1193), .ZN(n1173) );
NAND2_X1 U1067 ( .A1(n1347), .A2(n1348), .ZN(n1193) );
NAND2_X1 U1068 ( .A1(G128), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1069 ( .A(n1309), .B(KEYINPUT12), .Z(n1347) );
NAND2_X1 U1070 ( .A1(n1313), .A2(n1238), .ZN(n1309) );
INV_X1 U1071 ( .A(G128), .ZN(n1238) );
INV_X1 U1072 ( .A(n1349), .ZN(n1313) );
XNOR2_X1 U1073 ( .A(G143), .B(n1229), .ZN(n1349) );
INV_X1 U1074 ( .A(G146), .ZN(n1229) );
NAND2_X1 U1075 ( .A1(KEYINPUT44), .A2(n1195), .ZN(n1345) );
AND2_X1 U1076 ( .A1(n1350), .A2(G224), .ZN(n1195) );
XNOR2_X1 U1077 ( .A(n1183), .B(KEYINPUT55), .ZN(n1350) );
NAND2_X1 U1078 ( .A1(n1351), .A2(n1087), .ZN(n1233) );
NAND2_X1 U1079 ( .A1(G478), .A2(n1352), .ZN(n1087) );
XOR2_X1 U1080 ( .A(KEYINPUT7), .B(n1102), .Z(n1351) );
NOR2_X1 U1081 ( .A1(n1352), .A2(G478), .ZN(n1102) );
NAND2_X1 U1082 ( .A1(n1278), .A2(n1152), .ZN(n1352) );
NAND2_X1 U1083 ( .A1(n1353), .A2(n1354), .ZN(n1152) );
NAND2_X1 U1084 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
XOR2_X1 U1085 ( .A(n1357), .B(KEYINPUT27), .Z(n1353) );
OR2_X1 U1086 ( .A1(n1356), .A2(n1355), .ZN(n1357) );
XOR2_X1 U1087 ( .A(n1358), .B(n1359), .Z(n1355) );
XOR2_X1 U1088 ( .A(G107), .B(n1360), .Z(n1359) );
XNOR2_X1 U1089 ( .A(n1126), .B(G128), .ZN(n1360) );
INV_X1 U1090 ( .A(G134), .ZN(n1126) );
XNOR2_X1 U1091 ( .A(n1361), .B(n1362), .ZN(n1358) );
NOR2_X1 U1092 ( .A1(G143), .A2(KEYINPUT46), .ZN(n1362) );
NOR2_X1 U1093 ( .A1(KEYINPUT42), .A2(n1363), .ZN(n1361) );
XNOR2_X1 U1094 ( .A(n1287), .B(n1364), .ZN(n1363) );
NOR2_X1 U1095 ( .A1(G122), .A2(KEYINPUT60), .ZN(n1364) );
INV_X1 U1096 ( .A(G116), .ZN(n1287) );
NAND3_X1 U1097 ( .A1(n1259), .A2(G217), .A3(G234), .ZN(n1356) );
INV_X1 U1098 ( .A(n1183), .ZN(n1259) );
XOR2_X1 U1099 ( .A(G953), .B(KEYINPUT0), .Z(n1183) );
INV_X1 U1100 ( .A(n1252), .ZN(n1278) );
XOR2_X1 U1101 ( .A(G902), .B(KEYINPUT8), .Z(n1252) );
INV_X1 U1102 ( .A(G110), .ZN(n1248) );
endmodule


