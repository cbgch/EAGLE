//Key = 0100111011100111110000001111000101001010111100011001111010110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U742 ( .A(G107), .B(n1023), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n1025) );
NOR4_X1 U745 ( .A1(n1027), .A2(n1028), .A3(n1026), .A4(n1029), .ZN(n1024) );
NOR2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
AND4_X1 U747 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1030) );
AND4_X1 U748 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1026) );
NOR3_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1034), .ZN(n1039) );
XOR2_X1 U750 ( .A(n1042), .B(G469), .Z(n1038) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1037) );
XOR2_X1 U752 ( .A(KEYINPUT50), .B(n1045), .Z(n1036) );
NOR3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
XOR2_X1 U754 ( .A(KEYINPUT18), .B(n1049), .Z(n1048) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
XOR2_X1 U756 ( .A(KEYINPUT7), .B(n1052), .Z(n1047) );
NAND3_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(n1054) );
XOR2_X1 U759 ( .A(KEYINPUT6), .B(G472), .Z(n1051) );
INV_X1 U760 ( .A(n1056), .ZN(n1050) );
XOR2_X1 U761 ( .A(KEYINPUT12), .B(n1057), .Z(n1053) );
NOR2_X1 U762 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
XOR2_X1 U763 ( .A(n1060), .B(KEYINPUT27), .Z(n1059) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
INV_X1 U765 ( .A(n1063), .ZN(n1028) );
NAND3_X1 U766 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1027) );
NAND4_X1 U767 ( .A1(n1033), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1066) );
NAND3_X1 U768 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U770 ( .A(n1075), .B(KEYINPUT58), .ZN(n1073) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
OR2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
AND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1068) );
NAND2_X1 U774 ( .A1(n1035), .A2(n1082), .ZN(n1064) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U776 ( .A1(n1085), .A2(n1086), .A3(n1032), .ZN(n1084) );
INV_X1 U777 ( .A(n1087), .ZN(n1032) );
NAND2_X1 U778 ( .A1(n1034), .A2(n1088), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1033), .A2(n1031), .ZN(n1088) );
INV_X1 U780 ( .A(KEYINPUT3), .ZN(n1031) );
NAND3_X1 U781 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1085) );
NAND2_X1 U782 ( .A1(n1040), .A2(n1092), .ZN(n1089) );
AND4_X1 U783 ( .A1(n1075), .A2(n1076), .A3(n1081), .A4(n1080), .ZN(n1035) );
INV_X1 U784 ( .A(KEYINPUT34), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(G72) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
INV_X1 U787 ( .A(n1097), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
NAND2_X1 U789 ( .A1(n1099), .A2(n1096), .ZN(n1098) );
NAND2_X1 U790 ( .A1(G953), .A2(n1100), .ZN(n1096) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(n1097) );
AND2_X1 U792 ( .A1(n1103), .A2(n1065), .ZN(n1102) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1099), .ZN(n1101) );
INV_X1 U794 ( .A(n1105), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1104) );
NAND2_X1 U796 ( .A1(n1108), .A2(KEYINPUT4), .ZN(n1106) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U798 ( .A(n1111), .B(G131), .Z(n1109) );
NAND2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U801 ( .A(KEYINPUT61), .B(n1116), .Z(n1112) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1114), .ZN(n1116) );
XOR2_X1 U803 ( .A(KEYINPUT23), .B(G134), .Z(n1114) );
XOR2_X1 U804 ( .A(n1117), .B(n1118), .Z(G69) );
NOR3_X1 U805 ( .A1(KEYINPUT44), .A2(n1119), .A3(n1120), .ZN(n1118) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U807 ( .A(KEYINPUT53), .B(n1123), .Z(n1122) );
INV_X1 U808 ( .A(n1124), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
NAND2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U811 ( .A1(G953), .A2(n1127), .ZN(n1126) );
XOR2_X1 U812 ( .A(n1128), .B(KEYINPUT55), .Z(n1125) );
AND2_X1 U813 ( .A1(n1065), .A2(n1129), .ZN(n1123) );
NAND2_X1 U814 ( .A1(G953), .A2(n1130), .ZN(n1117) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U818 ( .A(n1135), .B(KEYINPUT40), .Z(n1133) );
NAND3_X1 U819 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
OR2_X1 U820 ( .A1(n1139), .A2(KEYINPUT21), .ZN(n1137) );
NAND2_X1 U821 ( .A1(KEYINPUT21), .A2(n1140), .ZN(n1136) );
NAND2_X1 U822 ( .A1(n1063), .A2(G902), .ZN(n1140) );
NOR2_X1 U823 ( .A1(n1131), .A2(n1141), .ZN(G63) );
XOR2_X1 U824 ( .A(n1142), .B(n1143), .Z(n1141) );
AND2_X1 U825 ( .A1(G478), .A2(n1139), .ZN(n1143) );
AND3_X1 U826 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1142) );
INV_X1 U827 ( .A(KEYINPUT60), .ZN(n1145) );
NOR2_X1 U828 ( .A1(n1131), .A2(n1147), .ZN(G60) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U830 ( .A1(n1139), .A2(G475), .ZN(n1148) );
XOR2_X1 U831 ( .A(G104), .B(n1150), .Z(G6) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(G57) );
XOR2_X1 U833 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U834 ( .A(n1155), .B(KEYINPUT0), .ZN(n1154) );
NAND3_X1 U835 ( .A1(n1139), .A2(G472), .A3(KEYINPUT36), .ZN(n1155) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1153) );
NOR2_X1 U837 ( .A1(n1158), .A2(n1065), .ZN(n1151) );
XNOR2_X1 U838 ( .A(G952), .B(KEYINPUT26), .ZN(n1158) );
NOR2_X1 U839 ( .A1(n1131), .A2(n1159), .ZN(G54) );
XOR2_X1 U840 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U841 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NAND2_X1 U843 ( .A1(KEYINPUT38), .A2(n1166), .ZN(n1165) );
NAND2_X1 U844 ( .A1(KEYINPUT39), .A2(n1167), .ZN(n1164) );
INV_X1 U845 ( .A(n1166), .ZN(n1167) );
XOR2_X1 U846 ( .A(n1168), .B(n1169), .Z(n1166) );
XOR2_X1 U847 ( .A(n1170), .B(n1171), .Z(n1160) );
NOR2_X1 U848 ( .A1(KEYINPUT45), .A2(n1172), .ZN(n1171) );
XNOR2_X1 U849 ( .A(G110), .B(n1173), .ZN(n1172) );
NAND2_X1 U850 ( .A1(n1139), .A2(G469), .ZN(n1170) );
NOR2_X1 U851 ( .A1(n1131), .A2(n1174), .ZN(G51) );
XOR2_X1 U852 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U853 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U854 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
INV_X1 U855 ( .A(n1181), .ZN(n1180) );
NOR2_X1 U856 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
NOR2_X1 U857 ( .A1(KEYINPUT20), .A2(n1184), .ZN(n1182) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(n1177) );
NOR2_X1 U859 ( .A1(n1187), .A2(KEYINPUT20), .ZN(n1185) );
NOR2_X1 U860 ( .A1(n1181), .A2(n1183), .ZN(n1187) );
INV_X1 U861 ( .A(KEYINPUT13), .ZN(n1183) );
NAND2_X1 U862 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
NAND2_X1 U863 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U864 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
XNOR2_X1 U865 ( .A(KEYINPUT29), .B(n1191), .ZN(n1192) );
NAND2_X1 U866 ( .A1(n1139), .A2(n1043), .ZN(n1175) );
NOR2_X1 U867 ( .A1(n1194), .A2(n1063), .ZN(n1139) );
NOR2_X1 U868 ( .A1(n1129), .A2(n1103), .ZN(n1063) );
NAND4_X1 U869 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1103) );
AND4_X1 U870 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NOR2_X1 U871 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
NOR3_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1204) );
XOR2_X1 U873 ( .A(n1208), .B(KEYINPUT32), .Z(n1206) );
INV_X1 U874 ( .A(n1209), .ZN(n1203) );
NAND4_X1 U875 ( .A1(n1023), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1129) );
NOR4_X1 U876 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1150), .ZN(n1212) );
AND3_X1 U877 ( .A1(n1216), .A2(n1076), .A3(n1078), .ZN(n1150) );
NOR2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1214) );
NOR2_X1 U879 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U880 ( .A1(KEYINPUT43), .A2(n1221), .ZN(n1220) );
NOR3_X1 U881 ( .A1(n1222), .A2(KEYINPUT14), .A3(n1223), .ZN(n1219) );
NOR2_X1 U882 ( .A1(n1224), .A2(n1090), .ZN(n1213) );
NOR3_X1 U883 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1224) );
NOR2_X1 U884 ( .A1(n1221), .A2(n1228), .ZN(n1227) );
INV_X1 U885 ( .A(KEYINPUT43), .ZN(n1228) );
AND3_X1 U886 ( .A1(KEYINPUT14), .A2(n1229), .A3(n1230), .ZN(n1226) );
XOR2_X1 U887 ( .A(n1231), .B(KEYINPUT52), .Z(n1225) );
NAND3_X1 U888 ( .A1(n1079), .A2(n1076), .A3(n1216), .ZN(n1023) );
NOR2_X1 U889 ( .A1(n1065), .A2(G952), .ZN(n1131) );
XNOR2_X1 U890 ( .A(G146), .B(n1202), .ZN(G48) );
NAND3_X1 U891 ( .A1(n1078), .A2(n1217), .A3(n1232), .ZN(n1202) );
XOR2_X1 U892 ( .A(n1233), .B(n1209), .Z(G45) );
NAND4_X1 U893 ( .A1(n1234), .A2(n1217), .A3(n1074), .A4(n1235), .ZN(n1209) );
AND3_X1 U894 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
XOR2_X1 U895 ( .A(n1239), .B(n1240), .Z(G42) );
NAND2_X1 U896 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U897 ( .A(n1201), .B(n1243), .Z(G39) );
NAND2_X1 U898 ( .A1(KEYINPUT48), .A2(G137), .ZN(n1243) );
NAND3_X1 U899 ( .A1(n1033), .A2(n1075), .A3(n1232), .ZN(n1201) );
XNOR2_X1 U900 ( .A(n1244), .B(n1200), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1230), .A2(n1238), .A3(n1241), .ZN(n1200) );
INV_X1 U902 ( .A(n1222), .ZN(n1230) );
NAND2_X1 U903 ( .A1(KEYINPUT24), .A2(n1245), .ZN(n1244) );
INV_X1 U904 ( .A(G134), .ZN(n1245) );
NAND2_X1 U905 ( .A1(n1246), .A2(n1247), .ZN(G33) );
NAND2_X1 U906 ( .A1(G131), .A2(n1195), .ZN(n1247) );
XOR2_X1 U907 ( .A(KEYINPUT63), .B(n1248), .Z(n1246) );
NOR2_X1 U908 ( .A1(G131), .A2(n1195), .ZN(n1248) );
NAND4_X1 U909 ( .A1(n1241), .A2(n1078), .A3(n1074), .A4(n1238), .ZN(n1195) );
INV_X1 U910 ( .A(n1083), .ZN(n1241) );
NAND2_X1 U911 ( .A1(n1033), .A2(n1234), .ZN(n1083) );
INV_X1 U912 ( .A(n1205), .ZN(n1033) );
NAND2_X1 U913 ( .A1(n1092), .A2(n1249), .ZN(n1205) );
XOR2_X1 U914 ( .A(G128), .B(n1250), .Z(G30) );
NOR2_X1 U915 ( .A1(KEYINPUT11), .A2(n1196), .ZN(n1250) );
NAND3_X1 U916 ( .A1(n1079), .A2(n1217), .A3(n1232), .ZN(n1196) );
AND4_X1 U917 ( .A1(n1251), .A2(n1234), .A3(n1052), .A4(n1238), .ZN(n1232) );
XNOR2_X1 U918 ( .A(n1215), .B(n1252), .ZN(G3) );
NAND2_X1 U919 ( .A1(KEYINPUT42), .A2(G101), .ZN(n1252) );
AND3_X1 U920 ( .A1(n1075), .A2(n1216), .A3(n1074), .ZN(n1215) );
XNOR2_X1 U921 ( .A(G125), .B(n1199), .ZN(G27) );
NAND3_X1 U922 ( .A1(n1067), .A2(n1217), .A3(n1242), .ZN(n1199) );
INV_X1 U923 ( .A(n1207), .ZN(n1242) );
NAND4_X1 U924 ( .A1(n1253), .A2(n1078), .A3(n1052), .A4(n1238), .ZN(n1207) );
NAND2_X1 U925 ( .A1(n1254), .A2(n1255), .ZN(n1238) );
NAND3_X1 U926 ( .A1(G902), .A2(n1081), .A3(n1105), .ZN(n1255) );
NOR2_X1 U927 ( .A1(G900), .A2(n1065), .ZN(n1105) );
XOR2_X1 U928 ( .A(G122), .B(n1256), .Z(G24) );
NOR2_X1 U929 ( .A1(n1090), .A2(n1221), .ZN(n1256) );
NAND4_X1 U930 ( .A1(n1229), .A2(n1076), .A3(n1236), .A4(n1237), .ZN(n1221) );
NOR2_X1 U931 ( .A1(n1257), .A2(n1052), .ZN(n1076) );
XOR2_X1 U932 ( .A(G119), .B(n1258), .Z(G21) );
NOR2_X1 U933 ( .A1(n1090), .A2(n1231), .ZN(n1258) );
NAND4_X1 U934 ( .A1(n1251), .A2(n1229), .A3(n1075), .A4(n1052), .ZN(n1231) );
XOR2_X1 U935 ( .A(n1253), .B(KEYINPUT51), .Z(n1251) );
XOR2_X1 U936 ( .A(G116), .B(n1259), .Z(G18) );
NOR3_X1 U937 ( .A1(n1222), .A2(n1090), .A3(n1223), .ZN(n1259) );
NAND2_X1 U938 ( .A1(n1074), .A2(n1079), .ZN(n1222) );
NOR2_X1 U939 ( .A1(n1237), .A2(n1055), .ZN(n1079) );
XOR2_X1 U940 ( .A(n1260), .B(n1211), .Z(G15) );
NAND4_X1 U941 ( .A1(n1078), .A2(n1229), .A3(n1261), .A4(n1074), .ZN(n1211) );
NOR2_X1 U942 ( .A1(n1052), .A2(n1253), .ZN(n1074) );
INV_X1 U943 ( .A(n1223), .ZN(n1229) );
NAND2_X1 U944 ( .A1(n1067), .A2(n1262), .ZN(n1223) );
NOR2_X1 U945 ( .A1(n1087), .A2(n1034), .ZN(n1067) );
INV_X1 U946 ( .A(n1091), .ZN(n1034) );
AND2_X1 U947 ( .A1(n1055), .A2(n1237), .ZN(n1078) );
XNOR2_X1 U948 ( .A(G110), .B(n1210), .ZN(G12) );
NAND2_X1 U949 ( .A1(n1263), .A2(n1216), .ZN(n1210) );
AND3_X1 U950 ( .A1(n1261), .A2(n1262), .A3(n1234), .ZN(n1216) );
INV_X1 U951 ( .A(n1208), .ZN(n1234) );
NAND2_X1 U952 ( .A1(n1087), .A2(n1091), .ZN(n1208) );
NAND2_X1 U953 ( .A1(G221), .A2(n1264), .ZN(n1091) );
NAND3_X1 U954 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1087) );
NAND2_X1 U955 ( .A1(G469), .A2(n1268), .ZN(n1267) );
OR3_X1 U956 ( .A1(n1268), .A2(G469), .A3(KEYINPUT19), .ZN(n1266) );
AND2_X1 U957 ( .A1(KEYINPUT54), .A2(n1042), .ZN(n1268) );
NAND2_X1 U958 ( .A1(KEYINPUT19), .A2(n1269), .ZN(n1265) );
OR2_X1 U959 ( .A1(n1042), .A2(G469), .ZN(n1269) );
NAND2_X1 U960 ( .A1(n1270), .A2(n1194), .ZN(n1042) );
XOR2_X1 U961 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U962 ( .A(n1163), .B(n1273), .Z(n1272) );
XOR2_X1 U963 ( .A(KEYINPUT35), .B(KEYINPUT2), .Z(n1273) );
XNOR2_X1 U964 ( .A(n1169), .B(n1274), .ZN(n1271) );
XOR2_X1 U965 ( .A(n1275), .B(n1173), .Z(n1274) );
XOR2_X1 U966 ( .A(G140), .B(n1276), .Z(n1173) );
NOR2_X1 U967 ( .A1(G953), .A2(n1100), .ZN(n1276) );
INV_X1 U968 ( .A(G227), .ZN(n1100) );
XOR2_X1 U969 ( .A(G104), .B(n1110), .Z(n1169) );
XOR2_X1 U970 ( .A(n1190), .B(KEYINPUT16), .Z(n1110) );
NAND2_X1 U971 ( .A1(n1254), .A2(n1277), .ZN(n1262) );
NAND4_X1 U972 ( .A1(G953), .A2(G902), .A3(n1081), .A4(n1127), .ZN(n1277) );
INV_X1 U973 ( .A(G898), .ZN(n1127) );
NAND3_X1 U974 ( .A1(n1081), .A2(n1065), .A3(G952), .ZN(n1254) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1081) );
XOR2_X1 U976 ( .A(n1090), .B(KEYINPUT25), .Z(n1261) );
INV_X1 U977 ( .A(n1217), .ZN(n1090) );
NOR2_X1 U978 ( .A1(n1040), .A2(n1092), .ZN(n1217) );
NOR2_X1 U979 ( .A1(n1278), .A2(n1041), .ZN(n1092) );
NOR2_X1 U980 ( .A1(n1044), .A2(n1043), .ZN(n1041) );
AND2_X1 U981 ( .A1(n1043), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U982 ( .A(KEYINPUT15), .B(n1044), .ZN(n1279) );
NAND2_X1 U983 ( .A1(n1280), .A2(n1194), .ZN(n1044) );
XOR2_X1 U984 ( .A(n1281), .B(n1186), .Z(n1280) );
INV_X1 U985 ( .A(n1184), .ZN(n1186) );
XOR2_X1 U986 ( .A(n1128), .B(KEYINPUT30), .Z(n1184) );
XOR2_X1 U987 ( .A(n1282), .B(n1283), .Z(n1128) );
XOR2_X1 U988 ( .A(G113), .B(n1284), .Z(n1283) );
XOR2_X1 U989 ( .A(G119), .B(G116), .Z(n1284) );
XNOR2_X1 U990 ( .A(n1275), .B(n1285), .ZN(n1282) );
XOR2_X1 U991 ( .A(G110), .B(n1286), .Z(n1275) );
INV_X1 U992 ( .A(n1168), .ZN(n1286) );
XNOR2_X1 U993 ( .A(G101), .B(G107), .ZN(n1168) );
NAND2_X1 U994 ( .A1(n1287), .A2(KEYINPUT47), .ZN(n1281) );
XOR2_X1 U995 ( .A(n1190), .B(n1191), .Z(n1287) );
XNOR2_X1 U996 ( .A(G125), .B(n1288), .ZN(n1191) );
AND2_X1 U997 ( .A1(n1065), .A2(G224), .ZN(n1288) );
AND2_X1 U998 ( .A1(G210), .A2(n1289), .ZN(n1043) );
INV_X1 U999 ( .A(n1249), .ZN(n1040) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1289), .ZN(n1249) );
NAND2_X1 U1001 ( .A1(n1290), .A2(n1194), .ZN(n1289) );
XOR2_X1 U1002 ( .A(KEYINPUT8), .B(G237), .Z(n1290) );
INV_X1 U1003 ( .A(n1071), .ZN(n1263) );
NAND3_X1 U1004 ( .A1(n1253), .A2(n1052), .A3(n1075), .ZN(n1071) );
NOR2_X1 U1005 ( .A1(n1236), .A2(n1237), .ZN(n1075) );
NAND2_X1 U1006 ( .A1(n1060), .A2(n1291), .ZN(n1237) );
NAND2_X1 U1007 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U1008 ( .A(n1062), .B(KEYINPUT17), .Z(n1292) );
NAND2_X1 U1009 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U1010 ( .A(G475), .ZN(n1062) );
INV_X1 U1011 ( .A(n1293), .ZN(n1061) );
NAND2_X1 U1012 ( .A1(n1149), .A2(n1194), .ZN(n1293) );
XNOR2_X1 U1013 ( .A(n1285), .B(n1294), .ZN(n1149) );
XOR2_X1 U1014 ( .A(n1260), .B(n1295), .Z(n1294) );
NAND2_X1 U1015 ( .A1(n1296), .A2(KEYINPUT9), .ZN(n1295) );
XOR2_X1 U1016 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1017 ( .A(n1299), .B(n1300), .Z(n1298) );
NOR2_X1 U1018 ( .A1(KEYINPUT46), .A2(n1239), .ZN(n1299) );
XOR2_X1 U1019 ( .A(n1301), .B(n1302), .Z(n1297) );
XOR2_X1 U1020 ( .A(G131), .B(G125), .Z(n1302) );
NAND4_X1 U1021 ( .A1(KEYINPUT33), .A2(G214), .A3(n1303), .A4(n1065), .ZN(n1301) );
XOR2_X1 U1022 ( .A(G104), .B(G122), .Z(n1285) );
INV_X1 U1023 ( .A(n1055), .ZN(n1236) );
XOR2_X1 U1024 ( .A(n1304), .B(G478), .Z(n1055) );
NAND2_X1 U1025 ( .A1(n1194), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1026 ( .A1(n1144), .A2(n1146), .ZN(n1305) );
NAND4_X1 U1027 ( .A1(G217), .A2(G234), .A3(n1306), .A4(n1065), .ZN(n1146) );
XOR2_X1 U1028 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1029 ( .A(KEYINPUT59), .B(KEYINPUT37), .Z(n1308) );
NAND2_X1 U1030 ( .A1(n1307), .A2(n1309), .ZN(n1144) );
NAND3_X1 U1031 ( .A1(G234), .A2(n1065), .A3(G217), .ZN(n1309) );
XNOR2_X1 U1032 ( .A(n1310), .B(n1311), .ZN(n1307) );
XOR2_X1 U1033 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1034 ( .A(n1314), .B(G107), .Z(n1313) );
NAND2_X1 U1035 ( .A1(KEYINPUT56), .A2(n1233), .ZN(n1314) );
INV_X1 U1036 ( .A(G143), .ZN(n1233) );
NAND2_X1 U1037 ( .A1(KEYINPUT5), .A2(n1315), .ZN(n1312) );
INV_X1 U1038 ( .A(G122), .ZN(n1315) );
XOR2_X1 U1039 ( .A(n1316), .B(n1317), .Z(n1310) );
XOR2_X1 U1040 ( .A(KEYINPUT22), .B(G134), .Z(n1317) );
XNOR2_X1 U1041 ( .A(G116), .B(G128), .ZN(n1316) );
XNOR2_X1 U1042 ( .A(n1318), .B(n1138), .ZN(n1052) );
AND2_X1 U1043 ( .A1(G217), .A2(n1264), .ZN(n1138) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1194), .ZN(n1264) );
OR2_X1 U1045 ( .A1(n1134), .A2(G902), .ZN(n1318) );
XNOR2_X1 U1046 ( .A(n1319), .B(n1320), .ZN(n1134) );
XOR2_X1 U1047 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1048 ( .A(G146), .B(n1323), .ZN(n1322) );
NAND2_X1 U1049 ( .A1(KEYINPUT31), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1050 ( .A(G110), .B(n1325), .Z(n1324) );
XOR2_X1 U1051 ( .A(G128), .B(G119), .Z(n1325) );
NOR2_X1 U1052 ( .A1(KEYINPUT28), .A2(n1107), .ZN(n1321) );
XOR2_X1 U1053 ( .A(G125), .B(n1239), .Z(n1107) );
INV_X1 U1054 ( .A(G140), .ZN(n1239) );
XOR2_X1 U1055 ( .A(n1326), .B(n1327), .Z(n1319) );
AND3_X1 U1056 ( .A1(G221), .A2(n1065), .A3(G234), .ZN(n1327) );
NAND2_X1 U1057 ( .A1(KEYINPUT10), .A2(n1115), .ZN(n1326) );
INV_X1 U1058 ( .A(n1257), .ZN(n1253) );
XOR2_X1 U1059 ( .A(G472), .B(n1328), .Z(n1257) );
NOR2_X1 U1060 ( .A1(KEYINPUT62), .A2(n1056), .ZN(n1328) );
NAND2_X1 U1061 ( .A1(n1329), .A2(n1194), .ZN(n1056) );
INV_X1 U1062 ( .A(G902), .ZN(n1194) );
XOR2_X1 U1063 ( .A(n1330), .B(n1156), .Z(n1329) );
XOR2_X1 U1064 ( .A(n1331), .B(n1332), .Z(n1156) );
XOR2_X1 U1065 ( .A(G101), .B(n1333), .Z(n1332) );
AND3_X1 U1066 ( .A1(G210), .A2(n1065), .A3(n1303), .ZN(n1333) );
INV_X1 U1067 ( .A(G237), .ZN(n1303) );
INV_X1 U1068 ( .A(G953), .ZN(n1065) );
NAND2_X1 U1069 ( .A1(n1334), .A2(n1335), .ZN(n1331) );
NAND2_X1 U1070 ( .A1(n1336), .A2(n1260), .ZN(n1335) );
XOR2_X1 U1071 ( .A(n1337), .B(KEYINPUT49), .Z(n1334) );
OR2_X1 U1072 ( .A1(n1336), .A2(n1260), .ZN(n1337) );
INV_X1 U1073 ( .A(G113), .ZN(n1260) );
XNOR2_X1 U1074 ( .A(n1338), .B(G116), .ZN(n1336) );
NAND2_X1 U1075 ( .A1(KEYINPUT1), .A2(n1339), .ZN(n1338) );
INV_X1 U1076 ( .A(G119), .ZN(n1339) );
NAND2_X1 U1077 ( .A1(KEYINPUT41), .A2(n1157), .ZN(n1330) );
XOR2_X1 U1078 ( .A(n1190), .B(n1163), .Z(n1157) );
XNOR2_X1 U1079 ( .A(n1340), .B(n1341), .ZN(n1163) );
NOR2_X1 U1080 ( .A1(KEYINPUT57), .A2(n1115), .ZN(n1341) );
INV_X1 U1081 ( .A(G137), .ZN(n1115) );
XOR2_X1 U1082 ( .A(n1342), .B(G134), .Z(n1340) );
INV_X1 U1083 ( .A(G131), .ZN(n1342) );
INV_X1 U1084 ( .A(n1193), .ZN(n1190) );
XNOR2_X1 U1085 ( .A(G128), .B(n1300), .ZN(n1193) );
XOR2_X1 U1086 ( .A(G143), .B(G146), .Z(n1300) );
endmodule


