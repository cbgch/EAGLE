//Key = 0100011111110111100001111001110110001001001100010001010100101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362;

XNOR2_X1 U744 ( .A(G107), .B(n1037), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1039) );
NOR2_X1 U747 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U748 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR3_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NOR2_X1 U750 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U751 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U752 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U753 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U754 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U755 ( .A1(n1060), .A2(n1061), .ZN(n1054) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
AND2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1066), .A3(n1061), .ZN(n1050) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR3_X1 U760 ( .A1(n1053), .A2(n1069), .A3(n1061), .ZN(n1045) );
INV_X1 U761 ( .A(n1070), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U764 ( .A(n1075), .ZN(n1074) );
XNOR2_X1 U765 ( .A(n1076), .B(KEYINPUT59), .ZN(n1073) );
NOR3_X1 U766 ( .A1(n1077), .A2(n1047), .A3(n1057), .ZN(n1071) );
INV_X1 U767 ( .A(n1078), .ZN(n1053) );
NOR3_X1 U768 ( .A1(n1040), .A2(G953), .A3(G952), .ZN(n1038) );
AND4_X1 U769 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1040) );
NOR4_X1 U770 ( .A1(n1083), .A2(n1065), .A3(n1084), .A4(n1085), .ZN(n1082) );
INV_X1 U771 ( .A(n1086), .ZN(n1084) );
NAND3_X1 U772 ( .A1(n1087), .A2(n1077), .A3(n1088), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1081) );
NOR3_X1 U775 ( .A1(n1094), .A2(KEYINPUT57), .A3(n1095), .ZN(n1093) );
AND2_X1 U776 ( .A1(n1094), .A2(KEYINPUT57), .ZN(n1092) );
XNOR2_X1 U777 ( .A(n1096), .B(n1097), .ZN(n1091) );
XNOR2_X1 U778 ( .A(G475), .B(KEYINPUT33), .ZN(n1097) );
XNOR2_X1 U779 ( .A(n1098), .B(KEYINPUT54), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1099), .A2(n1100), .ZN(n1079) );
XOR2_X1 U781 ( .A(n1101), .B(KEYINPUT29), .Z(n1100) );
XOR2_X1 U782 ( .A(n1064), .B(KEYINPUT6), .Z(n1099) );
XOR2_X1 U783 ( .A(n1102), .B(n1103), .Z(G72) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR3_X1 U785 ( .A1(n1106), .A2(KEYINPUT50), .A3(G953), .ZN(n1105) );
NOR2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U788 ( .A(KEYINPUT48), .B(n1111), .ZN(n1110) );
XOR2_X1 U789 ( .A(n1112), .B(n1113), .Z(n1109) );
NAND2_X1 U790 ( .A1(KEYINPUT58), .A2(n1114), .ZN(n1112) );
INV_X1 U791 ( .A(G140), .ZN(n1114) );
NOR2_X1 U792 ( .A1(G900), .A2(n1115), .ZN(n1107) );
NOR2_X1 U793 ( .A1(n1116), .A2(n1115), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U795 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U797 ( .A1(n1115), .A2(n1123), .ZN(n1122) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U799 ( .A(n1126), .B(KEYINPUT43), .Z(n1124) );
NAND2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U801 ( .A(n1129), .B(KEYINPUT37), .Z(n1127) );
NAND2_X1 U802 ( .A1(n1130), .A2(n1131), .ZN(n1121) );
NAND2_X1 U803 ( .A1(G953), .A2(n1132), .ZN(n1131) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1130) );
NOR2_X1 U805 ( .A1(n1135), .A2(n1115), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U807 ( .A1(n1138), .A2(n1139), .ZN(G66) );
NOR3_X1 U808 ( .A1(n1089), .A2(n1140), .A3(n1141), .ZN(n1139) );
NOR4_X1 U809 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
INV_X1 U810 ( .A(n1146), .ZN(n1142) );
NOR2_X1 U811 ( .A1(n1147), .A2(n1146), .ZN(n1140) );
NOR3_X1 U812 ( .A1(n1145), .A2(n1148), .A3(n1144), .ZN(n1147) );
INV_X1 U813 ( .A(G217), .ZN(n1144) );
OR2_X1 U814 ( .A1(KEYINPUT38), .A2(n1149), .ZN(n1145) );
XOR2_X1 U815 ( .A(n1150), .B(KEYINPUT11), .Z(n1149) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1151), .ZN(G63) );
XOR2_X1 U817 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U818 ( .A1(n1094), .A2(n1143), .ZN(n1153) );
NOR2_X1 U819 ( .A1(n1138), .A2(n1154), .ZN(G60) );
NOR3_X1 U820 ( .A1(n1096), .A2(n1155), .A3(n1156), .ZN(n1154) );
NOR3_X1 U821 ( .A1(n1157), .A2(n1158), .A3(n1143), .ZN(n1156) );
NOR2_X1 U822 ( .A1(n1159), .A2(n1160), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1158), .ZN(n1159) );
INV_X1 U824 ( .A(n1042), .ZN(n1148) );
XNOR2_X1 U825 ( .A(n1161), .B(n1162), .ZN(G6) );
XOR2_X1 U826 ( .A(KEYINPUT25), .B(G104), .Z(n1162) );
NOR2_X1 U827 ( .A1(n1163), .A2(n1164), .ZN(G57) );
XOR2_X1 U828 ( .A(KEYINPUT17), .B(n1138), .Z(n1164) );
XOR2_X1 U829 ( .A(n1165), .B(n1166), .Z(n1163) );
NOR2_X1 U830 ( .A1(n1167), .A2(n1143), .ZN(n1165) );
NOR2_X1 U831 ( .A1(n1138), .A2(n1168), .ZN(G54) );
XNOR2_X1 U832 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U833 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U834 ( .A1(n1173), .A2(n1143), .ZN(n1172) );
NAND3_X1 U835 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1171) );
NAND2_X1 U836 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
OR3_X1 U837 ( .A1(n1178), .A2(n1177), .A3(n1179), .ZN(n1175) );
NOR2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
NAND2_X1 U839 ( .A1(n1179), .A2(n1178), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
XOR2_X1 U841 ( .A(KEYINPUT63), .B(n1180), .Z(n1183) );
NOR2_X1 U842 ( .A1(n1138), .A2(n1184), .ZN(G51) );
XOR2_X1 U843 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U844 ( .A1(n1187), .A2(n1143), .ZN(n1186) );
NAND2_X1 U845 ( .A1(G902), .A2(n1042), .ZN(n1143) );
NAND4_X1 U846 ( .A1(n1106), .A2(n1128), .A3(n1125), .A4(n1129), .ZN(n1042) );
NAND2_X1 U847 ( .A1(n1188), .A2(n1189), .ZN(n1129) );
XOR2_X1 U848 ( .A(KEYINPUT41), .B(n1190), .Z(n1189) );
NOR2_X1 U849 ( .A1(n1057), .A2(n1191), .ZN(n1190) );
AND4_X1 U850 ( .A1(n1161), .A2(n1192), .A3(n1193), .A4(n1037), .ZN(n1125) );
NAND3_X1 U851 ( .A1(n1067), .A2(n1070), .A3(n1194), .ZN(n1037) );
NAND3_X1 U852 ( .A1(n1194), .A2(n1070), .A3(n1068), .ZN(n1161) );
AND3_X1 U853 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1128) );
AND2_X1 U854 ( .A1(n1198), .A2(n1199), .ZN(n1106) );
NOR4_X1 U855 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U857 ( .A(KEYINPUT53), .B(n1206), .ZN(n1205) );
NOR4_X1 U858 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1198) );
AND4_X1 U859 ( .A1(n1068), .A2(n1059), .A3(n1211), .A4(n1076), .ZN(n1207) );
NAND2_X1 U860 ( .A1(KEYINPUT8), .A2(n1212), .ZN(n1185) );
XOR2_X1 U861 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U862 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U863 ( .A1(KEYINPUT62), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U864 ( .A(n1111), .B(n1218), .ZN(n1213) );
NOR3_X1 U865 ( .A1(n1137), .A2(KEYINPUT40), .A3(G953), .ZN(n1218) );
NOR2_X1 U866 ( .A1(n1115), .A2(G952), .ZN(n1138) );
NAND2_X1 U867 ( .A1(n1219), .A2(n1220), .ZN(G48) );
OR2_X1 U868 ( .A1(n1221), .A2(n1210), .ZN(n1220) );
XOR2_X1 U869 ( .A(n1222), .B(KEYINPUT61), .Z(n1219) );
NAND2_X1 U870 ( .A1(n1210), .A2(n1221), .ZN(n1222) );
NOR2_X1 U871 ( .A1(n1204), .A2(n1223), .ZN(n1210) );
INV_X1 U872 ( .A(n1068), .ZN(n1223) );
XNOR2_X1 U873 ( .A(G143), .B(n1224), .ZN(G45) );
NOR2_X1 U874 ( .A1(n1202), .A2(KEYINPUT12), .ZN(n1224) );
AND3_X1 U875 ( .A1(n1211), .A2(n1058), .A3(n1225), .ZN(n1202) );
AND3_X1 U876 ( .A1(n1063), .A2(n1226), .A3(n1227), .ZN(n1225) );
XNOR2_X1 U877 ( .A(n1201), .B(n1228), .ZN(G42) );
NAND2_X1 U878 ( .A1(KEYINPUT24), .A2(G140), .ZN(n1228) );
AND3_X1 U879 ( .A1(n1068), .A2(n1229), .A3(n1059), .ZN(n1201) );
XOR2_X1 U880 ( .A(G137), .B(n1209), .Z(G39) );
AND2_X1 U881 ( .A1(n1230), .A2(n1229), .ZN(n1209) );
XNOR2_X1 U882 ( .A(n1200), .B(n1231), .ZN(G36) );
XOR2_X1 U883 ( .A(KEYINPUT5), .B(G134), .Z(n1231) );
AND3_X1 U884 ( .A1(n1058), .A2(n1067), .A3(n1229), .ZN(n1200) );
XOR2_X1 U885 ( .A(G131), .B(n1208), .Z(G33) );
AND3_X1 U886 ( .A1(n1229), .A2(n1058), .A3(n1068), .ZN(n1208) );
AND4_X1 U887 ( .A1(n1232), .A2(n1063), .A3(n1233), .A4(n1077), .ZN(n1229) );
XNOR2_X1 U888 ( .A(n1234), .B(n1235), .ZN(G30) );
NOR2_X1 U889 ( .A1(n1206), .A2(n1204), .ZN(n1235) );
NAND4_X1 U890 ( .A1(n1211), .A2(n1063), .A3(n1098), .A4(n1236), .ZN(n1204) );
XNOR2_X1 U891 ( .A(G101), .B(n1192), .ZN(G3) );
NAND3_X1 U892 ( .A1(n1058), .A2(n1194), .A3(n1078), .ZN(n1192) );
XNOR2_X1 U893 ( .A(G125), .B(n1237), .ZN(G27) );
NAND4_X1 U894 ( .A1(n1076), .A2(n1211), .A3(n1068), .A4(n1238), .ZN(n1237) );
XOR2_X1 U895 ( .A(KEYINPUT49), .B(n1059), .Z(n1238) );
AND2_X1 U896 ( .A1(n1075), .A2(n1233), .ZN(n1211) );
NAND2_X1 U897 ( .A1(n1044), .A2(n1239), .ZN(n1233) );
NAND4_X1 U898 ( .A1(G953), .A2(G902), .A3(n1240), .A4(n1118), .ZN(n1239) );
INV_X1 U899 ( .A(G900), .ZN(n1118) );
XNOR2_X1 U900 ( .A(G122), .B(n1197), .ZN(G24) );
NAND4_X1 U901 ( .A1(n1241), .A2(n1070), .A3(n1227), .A4(n1226), .ZN(n1197) );
NOR2_X1 U902 ( .A1(n1236), .A2(n1098), .ZN(n1070) );
XNOR2_X1 U903 ( .A(G119), .B(n1195), .ZN(G21) );
NAND2_X1 U904 ( .A1(n1241), .A2(n1230), .ZN(n1195) );
AND3_X1 U905 ( .A1(n1098), .A2(n1236), .A3(n1078), .ZN(n1230) );
XNOR2_X1 U906 ( .A(G116), .B(n1196), .ZN(G18) );
NAND3_X1 U907 ( .A1(n1058), .A2(n1067), .A3(n1241), .ZN(n1196) );
AND3_X1 U908 ( .A1(n1075), .A2(n1242), .A3(n1076), .ZN(n1241) );
INV_X1 U909 ( .A(n1057), .ZN(n1076) );
INV_X1 U910 ( .A(n1206), .ZN(n1067) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1226), .ZN(n1206) );
XNOR2_X1 U912 ( .A(G113), .B(n1244), .ZN(G15) );
NAND3_X1 U913 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
XOR2_X1 U914 ( .A(n1188), .B(KEYINPUT0), .Z(n1247) );
XNOR2_X1 U915 ( .A(KEYINPUT20), .B(n1057), .ZN(n1246) );
NAND2_X1 U916 ( .A1(n1064), .A2(n1248), .ZN(n1057) );
INV_X1 U917 ( .A(n1191), .ZN(n1245) );
NAND3_X1 U918 ( .A1(n1058), .A2(n1242), .A3(n1068), .ZN(n1191) );
NOR2_X1 U919 ( .A1(n1226), .A2(n1243), .ZN(n1068) );
INV_X1 U920 ( .A(n1227), .ZN(n1243) );
NOR2_X1 U921 ( .A1(n1236), .A2(n1249), .ZN(n1058) );
XNOR2_X1 U922 ( .A(G110), .B(n1193), .ZN(G12) );
NAND3_X1 U923 ( .A1(n1059), .A2(n1194), .A3(n1078), .ZN(n1193) );
NOR2_X1 U924 ( .A1(n1226), .A2(n1227), .ZN(n1078) );
NAND2_X1 U925 ( .A1(n1250), .A2(n1251), .ZN(n1227) );
NAND2_X1 U926 ( .A1(n1096), .A2(n1158), .ZN(n1251) );
XOR2_X1 U927 ( .A(KEYINPUT16), .B(n1252), .Z(n1250) );
NOR2_X1 U928 ( .A1(n1096), .A2(n1158), .ZN(n1252) );
INV_X1 U929 ( .A(G475), .ZN(n1158) );
NOR2_X1 U930 ( .A1(n1160), .A2(G902), .ZN(n1096) );
INV_X1 U931 ( .A(n1157), .ZN(n1160) );
XNOR2_X1 U932 ( .A(n1253), .B(n1254), .ZN(n1157) );
XOR2_X1 U933 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U934 ( .A(G122), .B(n1257), .ZN(n1256) );
XNOR2_X1 U935 ( .A(n1258), .B(G131), .ZN(n1255) );
XOR2_X1 U936 ( .A(n1259), .B(n1260), .Z(n1253) );
XOR2_X1 U937 ( .A(G104), .B(n1261), .Z(n1260) );
AND3_X1 U938 ( .A1(G214), .A2(n1115), .A3(n1262), .ZN(n1261) );
NAND3_X1 U939 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1259) );
NAND2_X1 U940 ( .A1(KEYINPUT52), .A2(n1266), .ZN(n1265) );
NAND3_X1 U941 ( .A1(n1267), .A2(n1268), .A3(n1221), .ZN(n1264) );
NAND2_X1 U942 ( .A1(G146), .A2(n1269), .ZN(n1263) );
NAND2_X1 U943 ( .A1(n1270), .A2(n1268), .ZN(n1269) );
INV_X1 U944 ( .A(KEYINPUT52), .ZN(n1268) );
XNOR2_X1 U945 ( .A(KEYINPUT9), .B(n1267), .ZN(n1270) );
NAND2_X1 U946 ( .A1(n1271), .A2(n1086), .ZN(n1226) );
NAND2_X1 U947 ( .A1(n1095), .A2(n1094), .ZN(n1086) );
OR2_X1 U948 ( .A1(n1094), .A2(n1095), .ZN(n1271) );
NOR2_X1 U949 ( .A1(n1152), .A2(G902), .ZN(n1095) );
XOR2_X1 U950 ( .A(n1272), .B(n1273), .Z(n1152) );
AND3_X1 U951 ( .A1(G217), .A2(n1115), .A3(G234), .ZN(n1273) );
NAND2_X1 U952 ( .A1(n1274), .A2(KEYINPUT22), .ZN(n1272) );
XOR2_X1 U953 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U954 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U955 ( .A(n1234), .B(G122), .ZN(n1278) );
XOR2_X1 U956 ( .A(KEYINPUT55), .B(G134), .Z(n1277) );
XOR2_X1 U957 ( .A(n1279), .B(n1280), .Z(n1275) );
XNOR2_X1 U958 ( .A(n1281), .B(n1282), .ZN(n1279) );
NAND2_X1 U959 ( .A1(KEYINPUT42), .A2(n1258), .ZN(n1281) );
INV_X1 U960 ( .A(G143), .ZN(n1258) );
INV_X1 U961 ( .A(G478), .ZN(n1094) );
AND3_X1 U962 ( .A1(n1188), .A2(n1242), .A3(n1063), .ZN(n1194) );
NOR2_X1 U963 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U964 ( .A(n1248), .ZN(n1065) );
NAND2_X1 U965 ( .A1(G221), .A2(n1150), .ZN(n1248) );
XNOR2_X1 U966 ( .A(n1283), .B(n1173), .ZN(n1064) );
INV_X1 U967 ( .A(G469), .ZN(n1173) );
NAND2_X1 U968 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U969 ( .A(n1286), .B(n1287), .Z(n1284) );
XOR2_X1 U970 ( .A(n1181), .B(n1169), .Z(n1287) );
XNOR2_X1 U971 ( .A(n1288), .B(n1289), .ZN(n1169) );
XOR2_X1 U972 ( .A(G110), .B(n1290), .Z(n1289) );
NOR2_X1 U973 ( .A1(n1117), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U974 ( .A(KEYINPUT44), .B(n1115), .ZN(n1291) );
INV_X1 U975 ( .A(G227), .ZN(n1117) );
XNOR2_X1 U976 ( .A(G140), .B(KEYINPUT39), .ZN(n1288) );
INV_X1 U977 ( .A(n1182), .ZN(n1181) );
XOR2_X1 U978 ( .A(G101), .B(n1292), .Z(n1182) );
XNOR2_X1 U979 ( .A(n1282), .B(G104), .ZN(n1292) );
XNOR2_X1 U980 ( .A(n1113), .B(KEYINPUT31), .ZN(n1286) );
XOR2_X1 U981 ( .A(n1180), .B(n1178), .Z(n1113) );
NAND3_X1 U982 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1180) );
NAND2_X1 U983 ( .A1(KEYINPUT4), .A2(G128), .ZN(n1295) );
OR3_X1 U984 ( .A1(G128), .A2(KEYINPUT4), .A3(n1296), .ZN(n1294) );
NAND2_X1 U985 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
NAND2_X1 U986 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U987 ( .A(KEYINPUT4), .ZN(n1299) );
XNOR2_X1 U988 ( .A(G128), .B(KEYINPUT19), .ZN(n1298) );
XNOR2_X1 U989 ( .A(G143), .B(n1221), .ZN(n1296) );
NAND2_X1 U990 ( .A1(n1044), .A2(n1300), .ZN(n1242) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1132), .A4(n1240), .ZN(n1300) );
XNOR2_X1 U992 ( .A(KEYINPUT28), .B(n1136), .ZN(n1132) );
INV_X1 U993 ( .A(G898), .ZN(n1136) );
NAND3_X1 U994 ( .A1(n1240), .A2(n1115), .A3(G952), .ZN(n1044) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1240) );
XNOR2_X1 U996 ( .A(n1075), .B(KEYINPUT32), .ZN(n1188) );
NOR2_X1 U997 ( .A1(n1048), .A2(n1232), .ZN(n1075) );
INV_X1 U998 ( .A(n1047), .ZN(n1232) );
NAND2_X1 U999 ( .A1(n1301), .A2(n1101), .ZN(n1047) );
NAND2_X1 U1000 ( .A1(n1302), .A2(n1303), .ZN(n1101) );
XOR2_X1 U1001 ( .A(KEYINPUT51), .B(n1085), .Z(n1301) );
NOR2_X1 U1002 ( .A1(n1303), .A2(n1302), .ZN(n1085) );
INV_X1 U1003 ( .A(n1187), .ZN(n1302) );
NAND2_X1 U1004 ( .A1(G210), .A2(n1304), .ZN(n1187) );
NAND3_X1 U1005 ( .A1(n1305), .A2(n1306), .A3(n1285), .ZN(n1303) );
NAND2_X1 U1006 ( .A1(n1307), .A2(n1216), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1008 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
INV_X1 U1009 ( .A(KEYINPUT45), .ZN(n1311) );
NAND2_X1 U1010 ( .A1(KEYINPUT45), .A2(n1312), .ZN(n1308) );
OR2_X1 U1011 ( .A1(n1216), .A2(n1310), .ZN(n1305) );
NAND2_X1 U1012 ( .A1(KEYINPUT36), .A2(n1312), .ZN(n1310) );
XNOR2_X1 U1013 ( .A(n1313), .B(n1137), .ZN(n1312) );
INV_X1 U1014 ( .A(G224), .ZN(n1137) );
NAND3_X1 U1015 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1313) );
NAND2_X1 U1016 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
INV_X1 U1017 ( .A(KEYINPUT21), .ZN(n1318) );
NAND3_X1 U1018 ( .A1(KEYINPUT21), .A2(n1319), .A3(n1111), .ZN(n1315) );
OR2_X1 U1019 ( .A1(n1111), .A2(n1319), .ZN(n1314) );
NOR2_X1 U1020 ( .A1(KEYINPUT35), .A2(n1317), .ZN(n1319) );
XNOR2_X1 U1021 ( .A(n1320), .B(KEYINPUT10), .ZN(n1317) );
XOR2_X1 U1022 ( .A(n1321), .B(n1134), .Z(n1216) );
XOR2_X1 U1023 ( .A(G110), .B(G122), .Z(n1134) );
NAND2_X1 U1024 ( .A1(KEYINPUT60), .A2(n1133), .ZN(n1321) );
XOR2_X1 U1025 ( .A(n1322), .B(n1323), .Z(n1133) );
XOR2_X1 U1026 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1027 ( .A(G104), .B(n1326), .ZN(n1325) );
INV_X1 U1028 ( .A(G101), .ZN(n1326) );
NOR2_X1 U1029 ( .A1(KEYINPUT56), .A2(n1257), .ZN(n1324) );
INV_X1 U1030 ( .A(G113), .ZN(n1257) );
XOR2_X1 U1031 ( .A(n1327), .B(n1328), .Z(n1322) );
NAND2_X1 U1032 ( .A1(KEYINPUT27), .A2(n1282), .ZN(n1327) );
INV_X1 U1033 ( .A(G107), .ZN(n1282) );
INV_X1 U1034 ( .A(n1077), .ZN(n1048) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1304), .ZN(n1077) );
NAND2_X1 U1036 ( .A1(n1329), .A2(n1262), .ZN(n1304) );
AND2_X1 U1037 ( .A1(n1249), .A2(n1236), .ZN(n1059) );
NAND3_X1 U1038 ( .A1(n1330), .A2(n1331), .A3(n1087), .ZN(n1236) );
NAND2_X1 U1039 ( .A1(n1332), .A2(n1333), .ZN(n1087) );
NAND2_X1 U1040 ( .A1(KEYINPUT30), .A2(n1333), .ZN(n1331) );
OR3_X1 U1041 ( .A1(n1332), .A2(KEYINPUT30), .A3(n1333), .ZN(n1330) );
INV_X1 U1042 ( .A(n1089), .ZN(n1333) );
NOR2_X1 U1043 ( .A1(n1146), .A2(G902), .ZN(n1089) );
NAND2_X1 U1044 ( .A1(n1334), .A2(n1335), .ZN(n1146) );
NAND2_X1 U1045 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1046 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1047 ( .A(n1340), .B(KEYINPUT18), .Z(n1336) );
NAND2_X1 U1048 ( .A1(n1341), .A2(n1342), .ZN(n1334) );
XNOR2_X1 U1049 ( .A(n1339), .B(n1338), .ZN(n1342) );
NAND2_X1 U1050 ( .A1(KEYINPUT47), .A2(n1343), .ZN(n1338) );
INV_X1 U1051 ( .A(G137), .ZN(n1343) );
XOR2_X1 U1052 ( .A(n1344), .B(KEYINPUT2), .Z(n1339) );
NAND3_X1 U1053 ( .A1(G234), .A2(n1115), .A3(n1345), .ZN(n1344) );
XNOR2_X1 U1054 ( .A(G221), .B(KEYINPUT14), .ZN(n1345) );
XOR2_X1 U1055 ( .A(n1340), .B(KEYINPUT15), .Z(n1341) );
XOR2_X1 U1056 ( .A(n1346), .B(n1347), .Z(n1340) );
XNOR2_X1 U1057 ( .A(n1348), .B(n1267), .ZN(n1347) );
INV_X1 U1058 ( .A(n1266), .ZN(n1267) );
XNOR2_X1 U1059 ( .A(G140), .B(n1111), .ZN(n1266) );
INV_X1 U1060 ( .A(G125), .ZN(n1111) );
NOR2_X1 U1061 ( .A1(KEYINPUT26), .A2(n1234), .ZN(n1348) );
XNOR2_X1 U1062 ( .A(G110), .B(n1349), .ZN(n1346) );
XNOR2_X1 U1063 ( .A(n1221), .B(G119), .ZN(n1349) );
INV_X1 U1064 ( .A(n1090), .ZN(n1332) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1350), .ZN(n1090) );
XNOR2_X1 U1066 ( .A(KEYINPUT7), .B(n1150), .ZN(n1350) );
NAND2_X1 U1067 ( .A1(n1329), .A2(G234), .ZN(n1150) );
XNOR2_X1 U1068 ( .A(G902), .B(KEYINPUT3), .ZN(n1329) );
INV_X1 U1069 ( .A(n1098), .ZN(n1249) );
XOR2_X1 U1070 ( .A(n1351), .B(n1167), .Z(n1098) );
INV_X1 U1071 ( .A(G472), .ZN(n1167) );
NAND2_X1 U1072 ( .A1(n1352), .A2(n1285), .ZN(n1351) );
INV_X1 U1073 ( .A(G902), .ZN(n1285) );
XOR2_X1 U1074 ( .A(KEYINPUT13), .B(n1166), .Z(n1352) );
XNOR2_X1 U1075 ( .A(n1353), .B(n1354), .ZN(n1166) );
XOR2_X1 U1076 ( .A(n1355), .B(n1356), .Z(n1354) );
XNOR2_X1 U1077 ( .A(G101), .B(G113), .ZN(n1356) );
NAND3_X1 U1078 ( .A1(n1262), .A2(n1115), .A3(n1357), .ZN(n1355) );
XOR2_X1 U1079 ( .A(KEYINPUT34), .B(G210), .Z(n1357) );
INV_X1 U1080 ( .A(G953), .ZN(n1115) );
INV_X1 U1081 ( .A(G237), .ZN(n1262) );
XNOR2_X1 U1082 ( .A(n1358), .B(n1217), .ZN(n1353) );
INV_X1 U1083 ( .A(n1320), .ZN(n1217) );
XNOR2_X1 U1084 ( .A(n1359), .B(n1360), .ZN(n1320) );
XNOR2_X1 U1085 ( .A(n1221), .B(n1361), .ZN(n1360) );
NOR2_X1 U1086 ( .A1(G143), .A2(KEYINPUT46), .ZN(n1361) );
INV_X1 U1087 ( .A(G146), .ZN(n1221) );
NAND2_X1 U1088 ( .A1(KEYINPUT1), .A2(n1234), .ZN(n1359) );
INV_X1 U1089 ( .A(G128), .ZN(n1234) );
XOR2_X1 U1090 ( .A(n1328), .B(n1178), .Z(n1358) );
XNOR2_X1 U1091 ( .A(G131), .B(n1362), .ZN(n1178) );
XOR2_X1 U1092 ( .A(G137), .B(G134), .Z(n1362) );
XOR2_X1 U1093 ( .A(G119), .B(n1280), .Z(n1328) );
XOR2_X1 U1094 ( .A(G116), .B(KEYINPUT23), .Z(n1280) );
endmodule


