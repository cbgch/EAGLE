//Key = 0110110011110000000100011000110100111001001110100001001110011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;

XOR2_X1 U724 ( .A(n1000), .B(G107), .Z(G9) );
NAND2_X1 U725 ( .A1(KEYINPUT11), .A2(n1001), .ZN(n1000) );
NAND3_X1 U726 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1001) );
NOR2_X1 U727 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR4_X1 U728 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
XOR2_X1 U729 ( .A(KEYINPUT17), .B(n1011), .Z(n1010) );
NOR4_X1 U730 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
XOR2_X1 U731 ( .A(KEYINPUT14), .B(n1016), .Z(n1008) );
NOR2_X1 U732 ( .A1(n1017), .A2(n1012), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U734 ( .A1(n1020), .A2(n1014), .ZN(n1019) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
AND2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(n1021) );
NOR2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR3_X1 U740 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1027) );
NOR3_X1 U741 ( .A1(n1015), .A2(n1026), .A3(n1035), .ZN(n1018) );
NAND3_X1 U742 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1007) );
NAND3_X1 U743 ( .A1(n1039), .A2(n1040), .A3(n1003), .ZN(n1038) );
NAND2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U745 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U746 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND2_X1 U749 ( .A1(n1024), .A2(n1051), .ZN(n1041) );
INV_X1 U750 ( .A(n1015), .ZN(n1024) );
NAND2_X1 U751 ( .A1(n1047), .A2(n1049), .ZN(n1015) );
NOR3_X1 U752 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1005) );
INV_X1 U753 ( .A(n1036), .ZN(n1052) );
NAND4_X1 U754 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1036) );
NOR4_X1 U755 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
XNOR2_X1 U756 ( .A(n1061), .B(n1062), .ZN(n1060) );
XOR2_X1 U757 ( .A(KEYINPUT31), .B(G475), .Z(n1062) );
AND2_X1 U758 ( .A1(n1063), .A2(G478), .ZN(n1059) );
INV_X1 U759 ( .A(n1029), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1030), .A2(n1064), .ZN(n1055) );
INV_X1 U761 ( .A(n1049), .ZN(n1030) );
XOR2_X1 U762 ( .A(n1065), .B(n1066), .Z(n1054) );
NAND2_X1 U763 ( .A1(n1067), .A2(KEYINPUT56), .ZN(n1066) );
XNOR2_X1 U764 ( .A(n1068), .B(KEYINPUT0), .ZN(n1067) );
XOR2_X1 U765 ( .A(KEYINPUT29), .B(n1031), .Z(n1053) );
INV_X1 U766 ( .A(n1069), .ZN(n1031) );
XOR2_X1 U767 ( .A(n1070), .B(n1071), .Z(G72) );
XOR2_X1 U768 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR3_X1 U769 ( .A1(n1074), .A2(KEYINPUT18), .A3(G953), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XNOR2_X1 U771 ( .A(KEYINPUT62), .B(n1077), .ZN(n1076) );
NAND2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1072) );
NAND2_X1 U773 ( .A1(G953), .A2(n1080), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1078) );
XOR2_X1 U775 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR2_X1 U776 ( .A1(KEYINPUT13), .A2(n1085), .ZN(n1083) );
XOR2_X1 U777 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U778 ( .A1(KEYINPUT32), .A2(n1088), .ZN(n1087) );
XOR2_X1 U779 ( .A(G125), .B(n1089), .Z(n1081) );
XOR2_X1 U780 ( .A(KEYINPUT6), .B(G140), .Z(n1089) );
NAND2_X1 U781 ( .A1(G953), .A2(n1090), .ZN(n1070) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1091), .B(n1092), .Z(G69) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
INV_X1 U786 ( .A(n1097), .ZN(n1096) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1095) );
XOR2_X1 U788 ( .A(KEYINPUT54), .B(KEYINPUT19), .Z(n1099) );
NAND2_X1 U789 ( .A1(n1037), .A2(n1100), .ZN(n1093) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U791 ( .A(n1103), .B(KEYINPUT58), .Z(n1101) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1037), .ZN(n1091) );
AND2_X1 U793 ( .A1(G224), .A2(G898), .ZN(n1104) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(G66) );
NOR3_X1 U795 ( .A1(n1068), .A2(n1107), .A3(n1108), .ZN(n1106) );
NOR3_X1 U796 ( .A1(n1109), .A2(n1065), .A3(n1110), .ZN(n1108) );
INV_X1 U797 ( .A(n1111), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1111), .ZN(n1107) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1065), .ZN(n1112) );
INV_X1 U800 ( .A(n1009), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1105), .A2(n1114), .ZN(G63) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U803 ( .A(KEYINPUT7), .B(n1117), .Z(n1116) );
AND2_X1 U804 ( .A1(G478), .A2(n1118), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1105), .A2(n1119), .ZN(G60) );
XOR2_X1 U806 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U807 ( .A1(KEYINPUT52), .A2(n1122), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1118), .A2(G475), .ZN(n1120) );
XOR2_X1 U809 ( .A(G104), .B(n1123), .Z(G6) );
NOR2_X1 U810 ( .A1(n1105), .A2(n1124), .ZN(G57) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U812 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U813 ( .A(G101), .B(n1129), .Z(n1125) );
AND2_X1 U814 ( .A1(G472), .A2(n1118), .ZN(n1129) );
NOR2_X1 U815 ( .A1(n1105), .A2(n1130), .ZN(G54) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1133) );
AND2_X1 U819 ( .A1(G469), .A2(n1118), .ZN(n1136) );
NAND2_X1 U820 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
XOR2_X1 U821 ( .A(KEYINPUT49), .B(KEYINPUT36), .Z(n1138) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1131) );
XOR2_X1 U823 ( .A(KEYINPUT23), .B(G140), .Z(n1140) );
NOR3_X1 U824 ( .A1(n1105), .A2(n1141), .A3(n1142), .ZN(G51) );
NOR2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XNOR2_X1 U826 ( .A(KEYINPUT63), .B(n1145), .ZN(n1144) );
NOR2_X1 U827 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
XOR2_X1 U828 ( .A(n1145), .B(KEYINPUT44), .Z(n1147) );
NAND2_X1 U829 ( .A1(n1118), .A2(n1148), .ZN(n1145) );
INV_X1 U830 ( .A(n1110), .ZN(n1118) );
NAND2_X1 U831 ( .A1(G902), .A2(n1009), .ZN(n1110) );
NAND4_X1 U832 ( .A1(n1149), .A2(n1102), .A3(n1077), .A4(n1103), .ZN(n1009) );
AND4_X1 U833 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1102) );
NOR3_X1 U834 ( .A1(n1154), .A2(n1155), .A3(n1123), .ZN(n1153) );
AND3_X1 U835 ( .A1(n1003), .A2(n1051), .A3(n1002), .ZN(n1123) );
NOR4_X1 U836 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1154) );
XOR2_X1 U837 ( .A(n1160), .B(KEYINPUT16), .Z(n1159) );
NAND2_X1 U838 ( .A1(n1004), .A2(n1003), .ZN(n1156) );
NAND2_X1 U839 ( .A1(n1043), .A2(n1161), .ZN(n1151) );
NAND2_X1 U840 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U841 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U842 ( .A1(n1023), .A2(n1002), .ZN(n1162) );
INV_X1 U843 ( .A(n1075), .ZN(n1149) );
NAND4_X1 U844 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1075) );
NOR3_X1 U845 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
INV_X1 U846 ( .A(n1173), .ZN(n1170) );
NAND2_X1 U847 ( .A1(n1050), .A2(n1174), .ZN(n1168) );
NAND2_X1 U848 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U849 ( .A1(n1177), .A2(n1049), .ZN(n1176) );
NAND2_X1 U850 ( .A1(n1178), .A2(n1004), .ZN(n1175) );
NOR2_X1 U851 ( .A1(n1037), .A2(G952), .ZN(n1105) );
XOR2_X1 U852 ( .A(n1179), .B(G146), .Z(G48) );
NAND2_X1 U853 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
OR2_X1 U854 ( .A1(n1077), .A2(KEYINPUT53), .ZN(n1181) );
NAND3_X1 U855 ( .A1(n1050), .A2(n1051), .A3(n1178), .ZN(n1077) );
NAND4_X1 U856 ( .A1(n1051), .A2(n1160), .A3(n1178), .A4(KEYINPUT53), .ZN(n1180) );
XNOR2_X1 U857 ( .A(G143), .B(n1166), .ZN(G45) );
NAND4_X1 U858 ( .A1(n1182), .A2(n1183), .A3(n1050), .A4(n1184), .ZN(n1166) );
NOR3_X1 U859 ( .A1(n1185), .A2(n1157), .A3(n1013), .ZN(n1184) );
NAND2_X1 U860 ( .A1(n1186), .A2(n1187), .ZN(G42) );
NAND2_X1 U861 ( .A1(G140), .A2(n1167), .ZN(n1187) );
XOR2_X1 U862 ( .A(KEYINPUT51), .B(n1188), .Z(n1186) );
NOR2_X1 U863 ( .A1(G140), .A2(n1167), .ZN(n1188) );
NAND3_X1 U864 ( .A1(n1047), .A2(n1048), .A3(n1177), .ZN(n1167) );
XOR2_X1 U865 ( .A(n1189), .B(n1173), .Z(G39) );
NAND3_X1 U866 ( .A1(n1178), .A2(n1043), .A3(n1047), .ZN(n1173) );
INV_X1 U867 ( .A(n1033), .ZN(n1047) );
NOR3_X1 U868 ( .A1(n1157), .A2(n1190), .A3(n1191), .ZN(n1178) );
XOR2_X1 U869 ( .A(G134), .B(n1172), .Z(G36) );
AND2_X1 U870 ( .A1(n1192), .A2(n1004), .ZN(n1172) );
XOR2_X1 U871 ( .A(G131), .B(n1171), .Z(G33) );
AND2_X1 U872 ( .A1(n1192), .A2(n1051), .ZN(n1171) );
NOR4_X1 U873 ( .A1(n1033), .A2(n1013), .A3(n1157), .A4(n1190), .ZN(n1192) );
NAND2_X1 U874 ( .A1(n1069), .A2(n1029), .ZN(n1033) );
XOR2_X1 U875 ( .A(n1193), .B(n1194), .Z(G30) );
NAND4_X1 U876 ( .A1(n1195), .A2(n1196), .A3(n1048), .A4(n1197), .ZN(n1194) );
NOR2_X1 U877 ( .A1(n1035), .A2(n1191), .ZN(n1197) );
XOR2_X1 U878 ( .A(KEYINPUT28), .B(n1190), .Z(n1196) );
INV_X1 U879 ( .A(n1182), .ZN(n1190) );
XOR2_X1 U880 ( .A(KEYINPUT33), .B(n1050), .Z(n1195) );
XOR2_X1 U881 ( .A(G101), .B(n1155), .Z(G3) );
NOR3_X1 U882 ( .A1(n1013), .A2(n1198), .A3(n1014), .ZN(n1155) );
XNOR2_X1 U883 ( .A(G125), .B(n1199), .ZN(G27) );
NAND3_X1 U884 ( .A1(n1177), .A2(n1049), .A3(n1200), .ZN(n1199) );
XOR2_X1 U885 ( .A(n1160), .B(KEYINPUT8), .Z(n1200) );
AND3_X1 U886 ( .A1(n1051), .A2(n1182), .A3(n1023), .ZN(n1177) );
NAND2_X1 U887 ( .A1(n1012), .A2(n1201), .ZN(n1182) );
NAND4_X1 U888 ( .A1(G902), .A2(G953), .A3(n1202), .A4(n1080), .ZN(n1201) );
INV_X1 U889 ( .A(G900), .ZN(n1080) );
XOR2_X1 U890 ( .A(n1203), .B(n1152), .Z(G24) );
NAND4_X1 U891 ( .A1(n1204), .A2(n1165), .A3(n1003), .A4(n1183), .ZN(n1152) );
INV_X1 U892 ( .A(n1026), .ZN(n1003) );
NAND2_X1 U893 ( .A1(n1205), .A2(n1206), .ZN(n1026) );
XOR2_X1 U894 ( .A(n1207), .B(KEYINPUT3), .Z(n1205) );
NAND2_X1 U895 ( .A1(n1208), .A2(n1209), .ZN(G21) );
NAND2_X1 U896 ( .A1(G119), .A2(n1210), .ZN(n1209) );
XOR2_X1 U897 ( .A(KEYINPUT42), .B(n1211), .Z(n1208) );
NOR2_X1 U898 ( .A1(G119), .A2(n1210), .ZN(n1211) );
NAND4_X1 U899 ( .A1(n1212), .A2(n1213), .A3(n1049), .A4(n1214), .ZN(n1210) );
NOR2_X1 U900 ( .A1(n1191), .A2(n1014), .ZN(n1214) );
INV_X1 U901 ( .A(n1164), .ZN(n1191) );
NOR2_X1 U902 ( .A1(n1207), .A2(n1206), .ZN(n1164) );
XOR2_X1 U903 ( .A(KEYINPUT26), .B(n1050), .Z(n1212) );
INV_X1 U904 ( .A(n1160), .ZN(n1050) );
XOR2_X1 U905 ( .A(n1103), .B(n1215), .Z(G18) );
NAND2_X1 U906 ( .A1(KEYINPUT34), .A2(G116), .ZN(n1215) );
NAND3_X1 U907 ( .A1(n1165), .A2(n1004), .A3(n1216), .ZN(n1103) );
INV_X1 U908 ( .A(n1035), .ZN(n1004) );
NAND2_X1 U909 ( .A1(n1185), .A2(n1183), .ZN(n1035) );
INV_X1 U910 ( .A(n1217), .ZN(n1183) );
XNOR2_X1 U911 ( .A(G113), .B(n1218), .ZN(G15) );
NAND2_X1 U912 ( .A1(KEYINPUT5), .A2(n1219), .ZN(n1218) );
INV_X1 U913 ( .A(n1150), .ZN(n1219) );
NAND3_X1 U914 ( .A1(n1165), .A2(n1051), .A3(n1216), .ZN(n1150) );
INV_X1 U915 ( .A(n1013), .ZN(n1216) );
NAND2_X1 U916 ( .A1(n1207), .A2(n1064), .ZN(n1013) );
NAND2_X1 U917 ( .A1(n1220), .A2(n1221), .ZN(n1051) );
OR2_X1 U918 ( .A1(n1014), .A2(KEYINPUT59), .ZN(n1221) );
NAND3_X1 U919 ( .A1(n1217), .A2(n1204), .A3(KEYINPUT59), .ZN(n1220) );
AND2_X1 U920 ( .A1(n1049), .A2(n1222), .ZN(n1165) );
NOR2_X1 U921 ( .A1(n1034), .A2(n1223), .ZN(n1049) );
INV_X1 U922 ( .A(n1032), .ZN(n1223) );
XNOR2_X1 U923 ( .A(G110), .B(n1224), .ZN(G12) );
NAND4_X1 U924 ( .A1(n1023), .A2(n1043), .A3(n1225), .A4(n1226), .ZN(n1224) );
OR2_X1 U925 ( .A1(n1002), .A2(KEYINPUT40), .ZN(n1226) );
INV_X1 U926 ( .A(n1198), .ZN(n1002) );
NAND2_X1 U927 ( .A1(n1222), .A2(n1048), .ZN(n1198) );
INV_X1 U928 ( .A(n1157), .ZN(n1048) );
NAND2_X1 U929 ( .A1(KEYINPUT40), .A2(n1227), .ZN(n1225) );
NAND2_X1 U930 ( .A1(n1222), .A2(n1157), .ZN(n1227) );
NAND2_X1 U931 ( .A1(n1034), .A2(n1032), .ZN(n1157) );
NAND2_X1 U932 ( .A1(G221), .A2(n1228), .ZN(n1032) );
XNOR2_X1 U933 ( .A(n1229), .B(G469), .ZN(n1034) );
NAND2_X1 U934 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U935 ( .A(n1232), .B(n1233), .Z(n1230) );
XNOR2_X1 U936 ( .A(n1234), .B(n1235), .ZN(n1233) );
NOR2_X1 U937 ( .A1(KEYINPUT21), .A2(G140), .ZN(n1235) );
NAND2_X1 U938 ( .A1(KEYINPUT10), .A2(n1139), .ZN(n1234) );
NAND2_X1 U939 ( .A1(G227), .A2(n1037), .ZN(n1139) );
XOR2_X1 U940 ( .A(n1134), .B(n1137), .Z(n1232) );
XNOR2_X1 U941 ( .A(n1236), .B(n1237), .ZN(n1134) );
XNOR2_X1 U942 ( .A(G107), .B(n1238), .ZN(n1237) );
XNOR2_X1 U943 ( .A(KEYINPUT47), .B(KEYINPUT37), .ZN(n1238) );
XOR2_X1 U944 ( .A(n1239), .B(n1240), .Z(n1236) );
XOR2_X1 U945 ( .A(n1084), .B(n1241), .Z(n1239) );
NOR2_X1 U946 ( .A1(n1160), .A2(n1158), .ZN(n1222) );
INV_X1 U947 ( .A(n1213), .ZN(n1158) );
NAND2_X1 U948 ( .A1(n1242), .A2(n1243), .ZN(n1213) );
NAND3_X1 U949 ( .A1(n1097), .A2(n1202), .A3(G902), .ZN(n1243) );
NOR2_X1 U950 ( .A1(n1037), .A2(G898), .ZN(n1097) );
XOR2_X1 U951 ( .A(KEYINPUT39), .B(n1039), .Z(n1242) );
INV_X1 U952 ( .A(n1012), .ZN(n1039) );
NAND3_X1 U953 ( .A1(n1202), .A2(n1037), .A3(G952), .ZN(n1012) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1202) );
NAND2_X1 U955 ( .A1(n1244), .A2(n1029), .ZN(n1160) );
NAND2_X1 U956 ( .A1(G214), .A2(n1245), .ZN(n1029) );
XOR2_X1 U957 ( .A(n1069), .B(KEYINPUT4), .Z(n1244) );
XOR2_X1 U958 ( .A(n1246), .B(n1148), .Z(n1069) );
AND2_X1 U959 ( .A1(G210), .A2(n1245), .ZN(n1148) );
NAND2_X1 U960 ( .A1(n1247), .A2(n1231), .ZN(n1245) );
INV_X1 U961 ( .A(G237), .ZN(n1247) );
NAND2_X1 U962 ( .A1(n1146), .A2(n1231), .ZN(n1246) );
INV_X1 U963 ( .A(n1143), .ZN(n1146) );
XOR2_X1 U964 ( .A(n1248), .B(n1249), .Z(n1143) );
XOR2_X1 U965 ( .A(G125), .B(n1250), .Z(n1249) );
AND2_X1 U966 ( .A1(n1037), .A2(G224), .ZN(n1250) );
XNOR2_X1 U967 ( .A(n1251), .B(n1098), .ZN(n1248) );
XNOR2_X1 U968 ( .A(n1252), .B(n1253), .ZN(n1098) );
XOR2_X1 U969 ( .A(n1254), .B(n1240), .Z(n1253) );
XOR2_X1 U970 ( .A(G110), .B(G101), .Z(n1240) );
XOR2_X1 U971 ( .A(n1255), .B(n1256), .Z(n1252) );
XOR2_X1 U972 ( .A(n1203), .B(n1257), .Z(n1256) );
NAND2_X1 U973 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U974 ( .A1(G107), .A2(n1241), .ZN(n1259) );
XOR2_X1 U975 ( .A(KEYINPUT9), .B(n1260), .Z(n1258) );
NOR2_X1 U976 ( .A1(G107), .A2(n1241), .ZN(n1260) );
INV_X1 U977 ( .A(G104), .ZN(n1241) );
NAND2_X1 U978 ( .A1(KEYINPUT2), .A2(G116), .ZN(n1255) );
INV_X1 U979 ( .A(n1014), .ZN(n1043) );
NAND2_X1 U980 ( .A1(n1217), .A2(n1185), .ZN(n1014) );
INV_X1 U981 ( .A(n1204), .ZN(n1185) );
XOR2_X1 U982 ( .A(n1261), .B(n1262), .Z(n1204) );
NOR2_X1 U983 ( .A1(KEYINPUT22), .A2(n1061), .ZN(n1262) );
NOR2_X1 U984 ( .A1(n1122), .A2(G902), .ZN(n1061) );
XOR2_X1 U985 ( .A(n1263), .B(n1264), .Z(n1122) );
XOR2_X1 U986 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U987 ( .A(G131), .B(G122), .Z(n1266) );
XOR2_X1 U988 ( .A(n1267), .B(n1268), .Z(n1263) );
XOR2_X1 U989 ( .A(G113), .B(n1269), .Z(n1268) );
NOR2_X1 U990 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U991 ( .A(n1272), .B(KEYINPUT43), .Z(n1271) );
NAND2_X1 U992 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NOR2_X1 U993 ( .A1(n1274), .A2(n1273), .ZN(n1270) );
XOR2_X1 U994 ( .A(KEYINPUT15), .B(G125), .Z(n1273) );
INV_X1 U995 ( .A(G140), .ZN(n1274) );
XOR2_X1 U996 ( .A(n1275), .B(n1276), .Z(n1267) );
NOR2_X1 U997 ( .A1(G104), .A2(KEYINPUT61), .ZN(n1276) );
NAND2_X1 U998 ( .A1(G214), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U999 ( .A(G475), .B(KEYINPUT20), .ZN(n1261) );
NOR2_X1 U1000 ( .A1(n1057), .A2(n1278), .ZN(n1217) );
AND2_X1 U1001 ( .A1(n1279), .A2(n1063), .ZN(n1278) );
XOR2_X1 U1002 ( .A(KEYINPUT48), .B(G478), .Z(n1279) );
NOR2_X1 U1003 ( .A1(n1063), .A2(G478), .ZN(n1057) );
NAND2_X1 U1004 ( .A1(n1280), .A2(n1231), .ZN(n1063) );
XNOR2_X1 U1005 ( .A(n1115), .B(KEYINPUT41), .ZN(n1280) );
XNOR2_X1 U1006 ( .A(n1281), .B(n1282), .ZN(n1115) );
XOR2_X1 U1007 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1008 ( .A(n1285), .B(n1286), .Z(n1284) );
NOR2_X1 U1009 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
INV_X1 U1010 ( .A(G217), .ZN(n1288) );
NAND2_X1 U1011 ( .A1(KEYINPUT24), .A2(G107), .ZN(n1285) );
XOR2_X1 U1012 ( .A(n1289), .B(n1290), .Z(n1281) );
XOR2_X1 U1013 ( .A(G128), .B(G116), .Z(n1290) );
XNOR2_X1 U1014 ( .A(n1291), .B(n1292), .ZN(n1289) );
NOR2_X1 U1015 ( .A1(KEYINPUT30), .A2(n1203), .ZN(n1292) );
INV_X1 U1016 ( .A(G122), .ZN(n1203) );
NOR2_X1 U1017 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1291) );
NOR2_X1 U1018 ( .A1(n1064), .A2(n1207), .ZN(n1023) );
XOR2_X1 U1019 ( .A(n1068), .B(n1065), .Z(n1207) );
NAND2_X1 U1020 ( .A1(G217), .A2(n1228), .ZN(n1065) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1231), .ZN(n1228) );
NOR2_X1 U1022 ( .A1(n1111), .A2(G902), .ZN(n1068) );
XOR2_X1 U1023 ( .A(n1293), .B(n1294), .Z(n1111) );
XOR2_X1 U1024 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1025 ( .A(G137), .B(G110), .Z(n1296) );
NOR2_X1 U1026 ( .A1(KEYINPUT38), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1027 ( .A(G119), .B(n1193), .Z(n1297) );
XOR2_X1 U1028 ( .A(n1298), .B(n1299), .Z(n1293) );
NOR2_X1 U1029 ( .A1(n1287), .A2(n1300), .ZN(n1299) );
INV_X1 U1030 ( .A(G221), .ZN(n1300) );
NAND2_X1 U1031 ( .A1(n1301), .A2(n1037), .ZN(n1287) );
INV_X1 U1032 ( .A(G953), .ZN(n1037) );
XNOR2_X1 U1033 ( .A(G234), .B(KEYINPUT35), .ZN(n1301) );
NAND3_X1 U1034 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1298) );
NAND2_X1 U1035 ( .A1(KEYINPUT57), .A2(n1305), .ZN(n1304) );
OR3_X1 U1036 ( .A1(n1305), .A2(KEYINPUT57), .A3(G146), .ZN(n1303) );
NAND2_X1 U1037 ( .A1(G146), .A2(n1306), .ZN(n1302) );
NAND2_X1 U1038 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
INV_X1 U1039 ( .A(KEYINPUT57), .ZN(n1308) );
XNOR2_X1 U1040 ( .A(n1305), .B(KEYINPUT50), .ZN(n1307) );
XNOR2_X1 U1041 ( .A(n1309), .B(G125), .ZN(n1305) );
NAND2_X1 U1042 ( .A1(KEYINPUT55), .A2(G140), .ZN(n1309) );
INV_X1 U1043 ( .A(n1206), .ZN(n1064) );
XOR2_X1 U1044 ( .A(n1310), .B(G472), .Z(n1206) );
NAND2_X1 U1045 ( .A1(n1311), .A2(n1231), .ZN(n1310) );
INV_X1 U1046 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1047 ( .A(n1127), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1048 ( .A(n1313), .B(n1314), .ZN(n1312) );
NOR2_X1 U1049 ( .A1(KEYINPUT45), .A2(n1315), .ZN(n1314) );
INV_X1 U1050 ( .A(G101), .ZN(n1315) );
NOR2_X1 U1051 ( .A1(KEYINPUT27), .A2(n1128), .ZN(n1313) );
XNOR2_X1 U1052 ( .A(n1137), .B(n1251), .ZN(n1128) );
XOR2_X1 U1053 ( .A(n1084), .B(KEYINPUT60), .Z(n1251) );
XNOR2_X1 U1054 ( .A(n1193), .B(n1265), .ZN(n1084) );
XOR2_X1 U1055 ( .A(G146), .B(G143), .Z(n1265) );
INV_X1 U1056 ( .A(G128), .ZN(n1193) );
XOR2_X1 U1057 ( .A(n1086), .B(n1316), .Z(n1137) );
XOR2_X1 U1058 ( .A(KEYINPUT1), .B(n1088), .Z(n1316) );
INV_X1 U1059 ( .A(n1283), .ZN(n1088) );
XNOR2_X1 U1060 ( .A(G134), .B(KEYINPUT12), .ZN(n1283) );
XOR2_X1 U1061 ( .A(G131), .B(n1189), .Z(n1086) );
INV_X1 U1062 ( .A(G137), .ZN(n1189) );
XNOR2_X1 U1063 ( .A(n1317), .B(n1318), .ZN(n1127) );
XOR2_X1 U1064 ( .A(KEYINPUT46), .B(G116), .Z(n1318) );
XOR2_X1 U1065 ( .A(n1319), .B(n1254), .Z(n1317) );
XOR2_X1 U1066 ( .A(G113), .B(G119), .Z(n1254) );
NAND2_X1 U1067 ( .A1(G210), .A2(n1277), .ZN(n1319) );
NOR2_X1 U1068 ( .A1(G953), .A2(G237), .ZN(n1277) );
endmodule


