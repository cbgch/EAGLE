//Key = 0001111001000011010011001101110000010111010111100011111111111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357;

XNOR2_X1 U747 ( .A(n1027), .B(n1028), .ZN(G9) );
NAND2_X1 U748 ( .A1(KEYINPUT4), .A2(G107), .ZN(n1028) );
NAND3_X1 U749 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(G75) );
NAND2_X1 U750 ( .A1(G952), .A2(n1032), .ZN(n1031) );
NAND3_X1 U751 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NAND2_X1 U752 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND3_X1 U754 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U759 ( .A1(n1051), .A2(n1052), .ZN(n1043) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U762 ( .A(n1057), .B(KEYINPUT8), .Z(n1053) );
NAND4_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1051), .A4(n1060), .ZN(n1038) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U765 ( .A1(n1042), .A2(n1040), .ZN(n1062) );
NOR3_X1 U766 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1065), .ZN(n1067) );
XOR2_X1 U769 ( .A(KEYINPUT42), .B(n1045), .Z(n1068) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1058) );
NAND2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U772 ( .A1(n1073), .A2(n1065), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1045), .A2(n1074), .ZN(n1073) );
INV_X1 U774 ( .A(n1064), .ZN(n1045) );
NAND2_X1 U775 ( .A1(n1064), .A2(n1063), .ZN(n1071) );
INV_X1 U776 ( .A(KEYINPUT19), .ZN(n1063) );
NAND4_X1 U777 ( .A1(n1075), .A2(n1051), .A3(n1076), .A4(n1077), .ZN(n1029) );
NOR4_X1 U778 ( .A1(n1078), .A2(n1055), .A3(n1079), .A4(n1080), .ZN(n1077) );
XOR2_X1 U779 ( .A(n1056), .B(KEYINPUT28), .Z(n1080) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(n1079) );
NOR2_X1 U781 ( .A1(n1083), .A2(KEYINPUT32), .ZN(n1082) );
XOR2_X1 U782 ( .A(n1084), .B(n1085), .Z(n1076) );
XOR2_X1 U783 ( .A(n1069), .B(KEYINPUT18), .Z(n1075) );
XOR2_X1 U784 ( .A(n1086), .B(n1087), .Z(G72) );
NAND2_X1 U785 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U786 ( .A1(G900), .A2(n1089), .ZN(n1088) );
XOR2_X1 U787 ( .A(KEYINPUT31), .B(G227), .Z(n1089) );
NAND2_X1 U788 ( .A1(KEYINPUT38), .A2(n1090), .ZN(n1086) );
XOR2_X1 U789 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR3_X1 U790 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NOR2_X1 U791 ( .A1(G140), .A2(n1096), .ZN(n1095) );
XOR2_X1 U792 ( .A(KEYINPUT46), .B(n1097), .Z(n1096) );
NOR2_X1 U793 ( .A1(n1098), .A2(n1097), .ZN(n1094) );
XNOR2_X1 U794 ( .A(n1099), .B(n1100), .ZN(n1097) );
XOR2_X1 U795 ( .A(KEYINPUT49), .B(G125), .Z(n1100) );
NAND3_X1 U796 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1099) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1106), .A2(n1107), .ZN(n1102) );
INV_X1 U799 ( .A(KEYINPUT63), .ZN(n1107) );
NAND2_X1 U800 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
XOR2_X1 U801 ( .A(KEYINPUT50), .B(n1105), .Z(n1108) );
INV_X1 U802 ( .A(n1110), .ZN(n1105) );
NAND2_X1 U803 ( .A1(KEYINPUT63), .A2(n1111), .ZN(n1101) );
NAND2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U805 ( .A1(KEYINPUT50), .A2(n1109), .A3(n1110), .ZN(n1113) );
OR2_X1 U806 ( .A1(n1110), .A2(KEYINPUT50), .ZN(n1112) );
XOR2_X1 U807 ( .A(n1114), .B(n1115), .Z(n1110) );
NAND2_X1 U808 ( .A1(KEYINPUT17), .A2(n1116), .ZN(n1114) );
NOR2_X1 U809 ( .A1(G953), .A2(n1035), .ZN(n1091) );
XOR2_X1 U810 ( .A(n1117), .B(n1118), .Z(G69) );
NOR2_X1 U811 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR3_X1 U812 ( .A1(n1121), .A2(n1122), .A3(n1030), .ZN(n1120) );
NOR2_X1 U813 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U814 ( .A(KEYINPUT35), .ZN(n1121) );
NOR4_X1 U815 ( .A1(KEYINPUT35), .A2(n1124), .A3(n1030), .A4(n1123), .ZN(n1119) );
XOR2_X1 U816 ( .A(n1125), .B(n1126), .Z(n1117) );
NOR2_X1 U817 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U818 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U819 ( .A1(KEYINPUT39), .A2(n1131), .ZN(n1129) );
NOR2_X1 U820 ( .A1(G898), .A2(n1030), .ZN(n1127) );
NAND2_X1 U821 ( .A1(n1132), .A2(n1030), .ZN(n1125) );
NOR2_X1 U822 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U823 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U824 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U825 ( .A1(n1139), .A2(n1140), .ZN(G63) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U827 ( .A(KEYINPUT11), .B(n1143), .Z(n1142) );
NOR2_X1 U828 ( .A1(n1085), .A2(n1138), .ZN(n1143) );
NOR2_X1 U829 ( .A1(n1144), .A2(n1030), .ZN(n1139) );
XNOR2_X1 U830 ( .A(G952), .B(KEYINPUT44), .ZN(n1144) );
NOR2_X1 U831 ( .A1(n1133), .A2(n1145), .ZN(G60) );
NOR3_X1 U832 ( .A1(n1083), .A2(n1146), .A3(n1147), .ZN(n1145) );
NOR2_X1 U833 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1150), .A2(n1081), .ZN(n1148) );
NOR2_X1 U835 ( .A1(n1132), .A2(n1151), .ZN(n1150) );
NOR3_X1 U836 ( .A1(n1152), .A2(n1081), .A3(n1138), .ZN(n1146) );
INV_X1 U837 ( .A(G475), .ZN(n1081) );
XOR2_X1 U838 ( .A(G104), .B(n1153), .Z(G6) );
NOR3_X1 U839 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
NOR2_X1 U840 ( .A1(n1133), .A2(n1157), .ZN(G57) );
XOR2_X1 U841 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U842 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U843 ( .A(KEYINPUT24), .B(n1162), .Z(n1158) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1138), .ZN(n1162) );
XNOR2_X1 U845 ( .A(G472), .B(KEYINPUT30), .ZN(n1163) );
NOR2_X1 U846 ( .A1(n1133), .A2(n1164), .ZN(G54) );
XOR2_X1 U847 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U848 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U849 ( .A(n1169), .B(n1170), .Z(n1167) );
XOR2_X1 U850 ( .A(n1171), .B(n1172), .Z(n1165) );
XOR2_X1 U851 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U852 ( .A1(KEYINPUT16), .A2(n1109), .ZN(n1174) );
NOR2_X1 U853 ( .A1(n1175), .A2(n1138), .ZN(n1173) );
INV_X1 U854 ( .A(G469), .ZN(n1175) );
XOR2_X1 U855 ( .A(n1176), .B(KEYINPUT13), .Z(n1171) );
NOR2_X1 U856 ( .A1(n1133), .A2(n1177), .ZN(G51) );
XOR2_X1 U857 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U858 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U859 ( .A(G125), .B(n1182), .Z(n1181) );
NOR2_X1 U860 ( .A1(n1183), .A2(n1138), .ZN(n1180) );
NAND2_X1 U861 ( .A1(G902), .A2(n1184), .ZN(n1138) );
NAND2_X1 U862 ( .A1(n1035), .A2(n1033), .ZN(n1184) );
INV_X1 U863 ( .A(n1132), .ZN(n1033) );
NAND4_X1 U864 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1132) );
NOR4_X1 U865 ( .A1(n1027), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1188) );
INV_X1 U866 ( .A(n1192), .ZN(n1190) );
INV_X1 U867 ( .A(n1193), .ZN(n1189) );
NOR3_X1 U868 ( .A1(n1155), .A2(n1194), .A3(n1156), .ZN(n1027) );
NAND2_X1 U869 ( .A1(n1195), .A2(n1196), .ZN(n1187) );
NAND3_X1 U870 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
NAND2_X1 U871 ( .A1(KEYINPUT41), .A2(n1200), .ZN(n1199) );
NAND3_X1 U872 ( .A1(n1201), .A2(n1202), .A3(n1051), .ZN(n1198) );
NAND2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
INV_X1 U874 ( .A(KEYINPUT22), .ZN(n1204) );
NAND4_X1 U875 ( .A1(n1042), .A2(n1205), .A3(n1206), .A4(n1057), .ZN(n1186) );
INV_X1 U876 ( .A(n1207), .ZN(n1057) );
NAND2_X1 U877 ( .A1(n1208), .A2(n1209), .ZN(n1205) );
NAND2_X1 U878 ( .A1(KEYINPUT22), .A2(n1203), .ZN(n1209) );
NAND2_X1 U879 ( .A1(n1200), .A2(n1210), .ZN(n1208) );
INV_X1 U880 ( .A(KEYINPUT41), .ZN(n1210) );
NAND3_X1 U881 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1185) );
XOR2_X1 U882 ( .A(n1156), .B(KEYINPUT60), .Z(n1213) );
INV_X1 U883 ( .A(n1051), .ZN(n1156) );
INV_X1 U884 ( .A(n1151), .ZN(n1035) );
NAND4_X1 U885 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1151) );
NOR4_X1 U886 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
INV_X1 U887 ( .A(n1222), .ZN(n1220) );
NAND2_X1 U888 ( .A1(n1223), .A2(n1224), .ZN(n1216) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1074), .ZN(n1214) );
NAND2_X1 U890 ( .A1(n1194), .A2(n1154), .ZN(n1074) );
INV_X1 U891 ( .A(n1226), .ZN(n1194) );
XOR2_X1 U892 ( .A(n1227), .B(n1109), .Z(n1178) );
NOR2_X1 U893 ( .A1(n1030), .A2(G952), .ZN(n1133) );
XOR2_X1 U894 ( .A(n1228), .B(n1229), .Z(G48) );
NAND3_X1 U895 ( .A1(n1225), .A2(n1211), .A3(KEYINPUT56), .ZN(n1229) );
INV_X1 U896 ( .A(n1230), .ZN(n1225) );
XOR2_X1 U897 ( .A(n1231), .B(G143), .Z(G45) );
NAND2_X1 U898 ( .A1(KEYINPUT51), .A2(n1222), .ZN(n1231) );
NAND4_X1 U899 ( .A1(n1207), .A2(n1202), .A3(n1201), .A4(n1232), .ZN(n1222) );
NOR2_X1 U900 ( .A1(n1047), .A2(n1233), .ZN(n1232) );
NAND2_X1 U901 ( .A1(n1234), .A2(n1235), .ZN(G42) );
NAND2_X1 U902 ( .A1(G140), .A2(n1236), .ZN(n1235) );
XOR2_X1 U903 ( .A(KEYINPUT9), .B(n1237), .Z(n1234) );
NOR2_X1 U904 ( .A1(G140), .A2(n1236), .ZN(n1237) );
NAND3_X1 U905 ( .A1(n1223), .A2(n1238), .A3(n1239), .ZN(n1236) );
XOR2_X1 U906 ( .A(n1064), .B(KEYINPUT5), .Z(n1239) );
XOR2_X1 U907 ( .A(G137), .B(n1219), .Z(G39) );
AND2_X1 U908 ( .A1(n1200), .A2(n1224), .ZN(n1219) );
XOR2_X1 U909 ( .A(n1116), .B(n1215), .Z(G36) );
NAND3_X1 U910 ( .A1(n1240), .A2(n1226), .A3(n1224), .ZN(n1215) );
XOR2_X1 U911 ( .A(n1218), .B(n1241), .Z(G33) );
NOR2_X1 U912 ( .A1(KEYINPUT47), .A2(n1242), .ZN(n1241) );
INV_X1 U913 ( .A(G131), .ZN(n1242) );
AND2_X1 U914 ( .A1(n1203), .A2(n1224), .ZN(n1218) );
NOR2_X1 U915 ( .A1(n1233), .A2(n1064), .ZN(n1224) );
NAND2_X1 U916 ( .A1(n1056), .A2(n1243), .ZN(n1064) );
NOR2_X1 U917 ( .A1(n1047), .A2(n1154), .ZN(n1203) );
INV_X1 U918 ( .A(n1240), .ZN(n1047) );
XOR2_X1 U919 ( .A(G128), .B(n1244), .Z(G30) );
NOR2_X1 U920 ( .A1(n1230), .A2(n1245), .ZN(n1244) );
XOR2_X1 U921 ( .A(KEYINPUT27), .B(n1226), .Z(n1245) );
NAND4_X1 U922 ( .A1(n1238), .A2(n1207), .A3(n1050), .A4(n1246), .ZN(n1230) );
INV_X1 U923 ( .A(n1233), .ZN(n1238) );
NAND3_X1 U924 ( .A1(n1247), .A2(n1065), .A3(n1066), .ZN(n1233) );
XOR2_X1 U925 ( .A(G101), .B(n1191), .Z(G3) );
AND3_X1 U926 ( .A1(n1212), .A2(n1040), .A3(n1240), .ZN(n1191) );
XOR2_X1 U927 ( .A(G125), .B(n1221), .Z(G27) );
AND4_X1 U928 ( .A1(n1042), .A2(n1223), .A3(n1207), .A4(n1247), .ZN(n1221) );
NAND2_X1 U929 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND3_X1 U930 ( .A1(G902), .A2(n1037), .A3(n1093), .ZN(n1249) );
NOR2_X1 U931 ( .A1(n1030), .A2(G900), .ZN(n1093) );
AND3_X1 U932 ( .A1(n1049), .A2(n1050), .A3(n1211), .ZN(n1223) );
XNOR2_X1 U933 ( .A(G122), .B(n1250), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1201), .A2(n1195), .A3(n1251), .A4(n1202), .ZN(n1250) );
XOR2_X1 U935 ( .A(KEYINPUT34), .B(n1051), .Z(n1251) );
NOR2_X1 U936 ( .A1(n1246), .A2(n1050), .ZN(n1051) );
XOR2_X1 U937 ( .A(n1252), .B(n1253), .Z(G21) );
NAND3_X1 U938 ( .A1(n1195), .A2(n1200), .A3(KEYINPUT61), .ZN(n1253) );
AND3_X1 U939 ( .A1(n1050), .A2(n1246), .A3(n1040), .ZN(n1200) );
INV_X1 U940 ( .A(n1049), .ZN(n1246) );
XOR2_X1 U941 ( .A(n1254), .B(n1192), .Z(G18) );
NAND2_X1 U942 ( .A1(n1255), .A2(n1226), .ZN(n1192) );
XNOR2_X1 U943 ( .A(G113), .B(n1256), .ZN(G15) );
NAND2_X1 U944 ( .A1(n1255), .A2(n1211), .ZN(n1256) );
INV_X1 U945 ( .A(n1154), .ZN(n1211) );
NAND2_X1 U946 ( .A1(n1257), .A2(n1202), .ZN(n1154) );
XNOR2_X1 U947 ( .A(n1258), .B(KEYINPUT37), .ZN(n1202) );
XOR2_X1 U948 ( .A(KEYINPUT36), .B(n1259), .Z(n1257) );
AND2_X1 U949 ( .A1(n1195), .A2(n1240), .ZN(n1255) );
NOR2_X1 U950 ( .A1(n1050), .A2(n1049), .ZN(n1240) );
AND3_X1 U951 ( .A1(n1207), .A2(n1206), .A3(n1042), .ZN(n1195) );
NOR2_X1 U952 ( .A1(n1066), .A2(n1078), .ZN(n1042) );
INV_X1 U953 ( .A(n1065), .ZN(n1078) );
XOR2_X1 U954 ( .A(n1176), .B(n1193), .Z(G12) );
NAND4_X1 U955 ( .A1(n1049), .A2(n1212), .A3(n1040), .A4(n1050), .ZN(n1193) );
XOR2_X1 U956 ( .A(n1260), .B(n1137), .Z(n1050) );
NAND2_X1 U957 ( .A1(G217), .A2(n1261), .ZN(n1137) );
OR2_X1 U958 ( .A1(n1136), .A2(G902), .ZN(n1260) );
XNOR2_X1 U959 ( .A(n1262), .B(n1263), .ZN(n1136) );
XOR2_X1 U960 ( .A(G110), .B(n1264), .Z(n1263) );
XOR2_X1 U961 ( .A(G146), .B(G137), .Z(n1264) );
XOR2_X1 U962 ( .A(n1265), .B(n1266), .Z(n1262) );
XOR2_X1 U963 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U964 ( .A1(KEYINPUT25), .A2(n1269), .ZN(n1268) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1267) );
OR2_X1 U966 ( .A1(n1252), .A2(G128), .ZN(n1271) );
XOR2_X1 U967 ( .A(n1272), .B(KEYINPUT1), .Z(n1270) );
NAND2_X1 U968 ( .A1(G128), .A2(n1252), .ZN(n1272) );
INV_X1 U969 ( .A(G119), .ZN(n1252) );
NAND2_X1 U970 ( .A1(G221), .A2(n1273), .ZN(n1265) );
NAND2_X1 U971 ( .A1(n1274), .A2(n1275), .ZN(n1040) );
OR3_X1 U972 ( .A1(n1201), .A2(n1258), .A3(KEYINPUT36), .ZN(n1275) );
NAND2_X1 U973 ( .A1(KEYINPUT36), .A2(n1226), .ZN(n1274) );
NOR2_X1 U974 ( .A1(n1259), .A2(n1258), .ZN(n1226) );
XNOR2_X1 U975 ( .A(n1083), .B(n1276), .ZN(n1258) );
XOR2_X1 U976 ( .A(KEYINPUT29), .B(G475), .Z(n1276) );
NOR2_X1 U977 ( .A1(n1149), .A2(G902), .ZN(n1083) );
INV_X1 U978 ( .A(n1152), .ZN(n1149) );
XOR2_X1 U979 ( .A(n1277), .B(n1278), .Z(n1152) );
XNOR2_X1 U980 ( .A(G113), .B(n1279), .ZN(n1278) );
NAND2_X1 U981 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U982 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
INV_X1 U983 ( .A(G143), .ZN(n1283) );
XOR2_X1 U984 ( .A(KEYINPUT48), .B(n1284), .Z(n1282) );
NAND2_X1 U985 ( .A1(n1285), .A2(G143), .ZN(n1280) );
XOR2_X1 U986 ( .A(KEYINPUT53), .B(n1284), .Z(n1285) );
XNOR2_X1 U987 ( .A(n1286), .B(n1287), .ZN(n1284) );
XOR2_X1 U988 ( .A(G104), .B(n1288), .Z(n1287) );
AND3_X1 U989 ( .A1(G214), .A2(n1030), .A3(n1289), .ZN(n1288) );
NAND2_X1 U990 ( .A1(n1290), .A2(KEYINPUT14), .ZN(n1286) );
XOR2_X1 U991 ( .A(n1228), .B(n1269), .Z(n1290) );
XOR2_X1 U992 ( .A(G125), .B(G140), .Z(n1269) );
XNOR2_X1 U993 ( .A(G122), .B(n1291), .ZN(n1277) );
XOR2_X1 U994 ( .A(KEYINPUT55), .B(G131), .Z(n1291) );
INV_X1 U995 ( .A(n1201), .ZN(n1259) );
XOR2_X1 U996 ( .A(n1292), .B(n1084), .Z(n1201) );
NOR2_X1 U997 ( .A1(n1141), .A2(G902), .ZN(n1084) );
XNOR2_X1 U998 ( .A(n1293), .B(n1294), .ZN(n1141) );
XNOR2_X1 U999 ( .A(n1295), .B(n1296), .ZN(n1294) );
XNOR2_X1 U1000 ( .A(n1297), .B(n1298), .ZN(n1296) );
NOR2_X1 U1001 ( .A1(G122), .A2(KEYINPUT33), .ZN(n1298) );
NOR2_X1 U1002 ( .A1(G134), .A2(KEYINPUT0), .ZN(n1297) );
XOR2_X1 U1003 ( .A(n1299), .B(n1300), .Z(n1293) );
XOR2_X1 U1004 ( .A(n1254), .B(n1301), .Z(n1300) );
NAND2_X1 U1005 ( .A1(n1273), .A2(G217), .ZN(n1301) );
AND2_X1 U1006 ( .A1(G234), .A2(n1030), .ZN(n1273) );
NAND2_X1 U1007 ( .A1(KEYINPUT20), .A2(n1302), .ZN(n1299) );
INV_X1 U1008 ( .A(G107), .ZN(n1302) );
NAND2_X1 U1009 ( .A1(KEYINPUT54), .A2(n1085), .ZN(n1292) );
INV_X1 U1010 ( .A(G478), .ZN(n1085) );
INV_X1 U1011 ( .A(n1155), .ZN(n1212) );
NAND4_X1 U1012 ( .A1(n1207), .A2(n1066), .A3(n1206), .A4(n1065), .ZN(n1155) );
NAND2_X1 U1013 ( .A1(n1303), .A2(n1261), .ZN(n1065) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1304), .ZN(n1261) );
XOR2_X1 U1015 ( .A(KEYINPUT12), .B(G221), .Z(n1303) );
NAND2_X1 U1016 ( .A1(n1248), .A2(n1305), .ZN(n1206) );
NAND4_X1 U1017 ( .A1(G902), .A2(G953), .A3(n1037), .A4(n1124), .ZN(n1305) );
INV_X1 U1018 ( .A(G898), .ZN(n1124) );
NAND3_X1 U1019 ( .A1(n1306), .A2(n1030), .A3(G952), .ZN(n1248) );
XNOR2_X1 U1020 ( .A(KEYINPUT58), .B(n1037), .ZN(n1306) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1037) );
INV_X1 U1022 ( .A(n1069), .ZN(n1066) );
XOR2_X1 U1023 ( .A(n1307), .B(n1308), .Z(n1069) );
XOR2_X1 U1024 ( .A(KEYINPUT62), .B(G469), .Z(n1308) );
NAND2_X1 U1025 ( .A1(n1309), .A2(n1304), .ZN(n1307) );
XOR2_X1 U1026 ( .A(n1169), .B(n1310), .Z(n1309) );
XOR2_X1 U1027 ( .A(n1311), .B(n1312), .Z(n1310) );
NAND2_X1 U1028 ( .A1(KEYINPUT43), .A2(n1176), .ZN(n1312) );
NAND2_X1 U1029 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U1030 ( .A1(n1170), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1031 ( .A(n1316), .B(n1109), .Z(n1313) );
XNOR2_X1 U1032 ( .A(n1168), .B(n1317), .ZN(n1316) );
NOR2_X1 U1033 ( .A1(n1170), .A2(n1315), .ZN(n1317) );
INV_X1 U1034 ( .A(KEYINPUT57), .ZN(n1315) );
XNOR2_X1 U1035 ( .A(n1318), .B(n1319), .ZN(n1168) );
XOR2_X1 U1036 ( .A(G101), .B(n1320), .Z(n1319) );
NOR2_X1 U1037 ( .A1(G107), .A2(KEYINPUT26), .ZN(n1320) );
XNOR2_X1 U1038 ( .A(G104), .B(KEYINPUT59), .ZN(n1318) );
XOR2_X1 U1039 ( .A(n1098), .B(n1321), .Z(n1169) );
AND2_X1 U1040 ( .A1(n1030), .A2(G227), .ZN(n1321) );
INV_X1 U1041 ( .A(G953), .ZN(n1030) );
INV_X1 U1042 ( .A(G140), .ZN(n1098) );
NOR2_X1 U1043 ( .A1(n1056), .A2(n1055), .ZN(n1207) );
INV_X1 U1044 ( .A(n1243), .ZN(n1055) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1322), .ZN(n1243) );
XNOR2_X1 U1046 ( .A(n1323), .B(n1183), .ZN(n1056) );
NAND2_X1 U1047 ( .A1(G210), .A2(n1322), .ZN(n1183) );
NAND2_X1 U1048 ( .A1(n1289), .A2(n1304), .ZN(n1322) );
NAND2_X1 U1049 ( .A1(n1324), .A2(n1304), .ZN(n1323) );
XOR2_X1 U1050 ( .A(n1325), .B(n1326), .Z(n1324) );
INV_X1 U1051 ( .A(n1227), .ZN(n1326) );
XOR2_X1 U1052 ( .A(n1130), .B(n1131), .Z(n1227) );
XNOR2_X1 U1053 ( .A(n1327), .B(G101), .ZN(n1131) );
NAND2_X1 U1054 ( .A1(KEYINPUT15), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1055 ( .A(G107), .B(G104), .Z(n1328) );
XOR2_X1 U1056 ( .A(n1329), .B(n1330), .Z(n1130) );
XOR2_X1 U1057 ( .A(G122), .B(G116), .Z(n1330) );
XOR2_X1 U1058 ( .A(n1176), .B(n1331), .Z(n1329) );
NAND2_X1 U1059 ( .A1(n1332), .A2(n1333), .ZN(n1325) );
NAND2_X1 U1060 ( .A1(n1182), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1061 ( .A(n1335), .B(KEYINPUT7), .Z(n1332) );
OR2_X1 U1062 ( .A1(n1334), .A2(n1182), .ZN(n1335) );
NOR2_X1 U1063 ( .A1(n1123), .A2(G953), .ZN(n1182) );
INV_X1 U1064 ( .A(G224), .ZN(n1123) );
XNOR2_X1 U1065 ( .A(n1104), .B(n1336), .ZN(n1334) );
NOR2_X1 U1066 ( .A1(G125), .A2(KEYINPUT10), .ZN(n1336) );
XOR2_X1 U1067 ( .A(n1337), .B(G472), .Z(n1049) );
NAND4_X1 U1068 ( .A1(n1338), .A2(n1304), .A3(n1339), .A4(n1340), .ZN(n1337) );
NAND3_X1 U1069 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1340) );
NAND2_X1 U1070 ( .A1(KEYINPUT40), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1071 ( .A(KEYINPUT23), .B(KEYINPUT3), .ZN(n1341) );
NAND3_X1 U1072 ( .A1(n1345), .A2(n1346), .A3(n1160), .ZN(n1339) );
NAND2_X1 U1073 ( .A1(n1344), .A2(n1347), .ZN(n1346) );
INV_X1 U1074 ( .A(KEYINPUT40), .ZN(n1347) );
NAND2_X1 U1075 ( .A1(KEYINPUT21), .A2(n1161), .ZN(n1344) );
INV_X1 U1076 ( .A(n1348), .ZN(n1161) );
XOR2_X1 U1077 ( .A(KEYINPUT3), .B(KEYINPUT23), .Z(n1345) );
INV_X1 U1078 ( .A(G902), .ZN(n1304) );
NAND2_X1 U1079 ( .A1(n1348), .A2(n1349), .ZN(n1338) );
NAND2_X1 U1080 ( .A1(KEYINPUT21), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1081 ( .A(KEYINPUT40), .B(n1160), .Z(n1350) );
INV_X1 U1082 ( .A(n1343), .ZN(n1160) );
XOR2_X1 U1083 ( .A(n1351), .B(G101), .Z(n1343) );
NAND3_X1 U1084 ( .A1(n1352), .A2(n1289), .A3(G210), .ZN(n1351) );
INV_X1 U1085 ( .A(G237), .ZN(n1289) );
XOR2_X1 U1086 ( .A(KEYINPUT45), .B(G953), .Z(n1352) );
XOR2_X1 U1087 ( .A(n1353), .B(n1354), .Z(n1348) );
XOR2_X1 U1088 ( .A(n1109), .B(n1331), .Z(n1354) );
XOR2_X1 U1089 ( .A(G113), .B(G119), .Z(n1331) );
INV_X1 U1090 ( .A(n1104), .ZN(n1109) );
XOR2_X1 U1091 ( .A(n1228), .B(n1295), .Z(n1104) );
XOR2_X1 U1092 ( .A(G128), .B(G143), .Z(n1295) );
INV_X1 U1093 ( .A(G146), .ZN(n1228) );
XOR2_X1 U1094 ( .A(n1355), .B(n1170), .Z(n1353) );
XNOR2_X1 U1095 ( .A(n1356), .B(n1115), .ZN(n1170) );
XOR2_X1 U1096 ( .A(G131), .B(G137), .Z(n1115) );
XOR2_X1 U1097 ( .A(n1116), .B(KEYINPUT2), .Z(n1356) );
INV_X1 U1098 ( .A(G134), .ZN(n1116) );
XOR2_X1 U1099 ( .A(n1357), .B(KEYINPUT6), .Z(n1355) );
NAND2_X1 U1100 ( .A1(KEYINPUT52), .A2(n1254), .ZN(n1357) );
INV_X1 U1101 ( .A(G116), .ZN(n1254) );
INV_X1 U1102 ( .A(G110), .ZN(n1176) );
endmodule


