//Key = 0100001001001000011110010001010110110111011011010100100001110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334;

XOR2_X1 U736 ( .A(G107), .B(n1013), .Z(G9) );
NOR4_X1 U737 ( .A1(KEYINPUT15), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1013) );
NAND4_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(G75) );
NAND4_X1 U739 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1019) );
NOR4_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
INV_X1 U741 ( .A(n1029), .ZN(n1027) );
NAND3_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1025) );
NOR3_X1 U743 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1023) );
NOR2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1034) );
XOR2_X1 U746 ( .A(KEYINPUT39), .B(G475), .Z(n1039) );
XOR2_X1 U747 ( .A(n1040), .B(KEYINPUT22), .Z(n1033) );
XOR2_X1 U748 ( .A(n1041), .B(KEYINPUT33), .Z(n1021) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1018) );
NAND2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U751 ( .A1(n1041), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
NAND2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U755 ( .A1(n1055), .A2(n1029), .A3(n1028), .ZN(n1054) );
OR2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1049) );
NAND3_X1 U757 ( .A1(n1051), .A2(n1058), .A3(n1059), .ZN(n1044) );
NAND2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1041), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1026), .A2(n1014), .ZN(n1063) );
NAND3_X1 U761 ( .A1(n1064), .A2(n1065), .A3(n1048), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1046), .A2(n1066), .ZN(n1060) );
INV_X1 U763 ( .A(n1067), .ZN(n1042) );
XOR2_X1 U764 ( .A(n1068), .B(n1069), .Z(G72) );
NAND2_X1 U765 ( .A1(G953), .A2(n1070), .ZN(n1069) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1070) );
NAND2_X1 U767 ( .A1(KEYINPUT44), .A2(n1071), .ZN(n1068) );
XOR2_X1 U768 ( .A(n1072), .B(n1073), .Z(n1071) );
NAND2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U770 ( .A1(G953), .A2(n1076), .ZN(n1075) );
XNOR2_X1 U771 ( .A(n1077), .B(n1078), .ZN(n1074) );
XNOR2_X1 U772 ( .A(n1079), .B(n1080), .ZN(n1078) );
NOR2_X1 U773 ( .A1(KEYINPUT48), .A2(n1081), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR3_X1 U776 ( .A1(KEYINPUT41), .A2(G137), .A3(n1086), .ZN(n1085) );
INV_X1 U777 ( .A(G134), .ZN(n1086) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
INV_X1 U779 ( .A(KEYINPUT41), .ZN(n1088) );
INV_X1 U780 ( .A(G131), .ZN(n1082) );
NAND2_X1 U781 ( .A1(KEYINPUT12), .A2(n1089), .ZN(n1079) );
NAND3_X1 U782 ( .A1(KEYINPUT42), .A2(n1090), .A3(n1091), .ZN(n1072) );
XOR2_X1 U783 ( .A(n1020), .B(KEYINPUT28), .Z(n1091) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(G69) );
NAND2_X1 U785 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NAND2_X1 U786 ( .A1(G898), .A2(n1095), .ZN(n1094) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U788 ( .A(n1098), .B(KEYINPUT30), .Z(n1092) );
NAND2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U790 ( .A1(G953), .A2(n1097), .ZN(n1100) );
XNOR2_X1 U791 ( .A(n1101), .B(n1096), .ZN(n1099) );
XNOR2_X1 U792 ( .A(n1102), .B(KEYINPUT14), .ZN(n1096) );
NOR3_X1 U793 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(G66) );
NOR3_X1 U794 ( .A1(n1106), .A2(G953), .A3(G952), .ZN(n1105) );
AND2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
INV_X1 U796 ( .A(KEYINPUT25), .ZN(n1106) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1103) );
NOR2_X1 U798 ( .A1(n1037), .A2(n1110), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(G63) );
XNOR2_X1 U800 ( .A(n1107), .B(KEYINPUT59), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1111) );
AND2_X1 U802 ( .A1(G478), .A2(n1115), .ZN(n1114) );
NAND2_X1 U803 ( .A1(KEYINPUT35), .A2(n1116), .ZN(n1113) );
NOR2_X1 U804 ( .A1(n1107), .A2(n1117), .ZN(G60) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1110), .ZN(n1119) );
NAND2_X1 U807 ( .A1(KEYINPUT38), .A2(n1121), .ZN(n1118) );
XNOR2_X1 U808 ( .A(G104), .B(n1122), .ZN(G6) );
NAND4_X1 U809 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1014), .A2(n1127), .ZN(n1126) );
XOR2_X1 U811 ( .A(KEYINPUT10), .B(n1066), .Z(n1123) );
NOR2_X1 U812 ( .A1(n1107), .A2(n1128), .ZN(G57) );
XNOR2_X1 U813 ( .A(n1129), .B(n1130), .ZN(n1128) );
NAND3_X1 U814 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1129) );
NAND2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND3_X1 U816 ( .A1(n1115), .A2(G472), .A3(KEYINPUT1), .ZN(n1135) );
OR4_X1 U817 ( .A1(n1134), .A2(n1136), .A3(n1137), .A4(KEYINPUT60), .ZN(n1132) );
INV_X1 U818 ( .A(KEYINPUT1), .ZN(n1137) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1134) );
NAND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NAND2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U822 ( .A(n1144), .B(KEYINPUT6), .Z(n1143) );
XOR2_X1 U823 ( .A(n1145), .B(KEYINPUT29), .Z(n1142) );
XOR2_X1 U824 ( .A(n1146), .B(KEYINPUT62), .Z(n1140) );
NAND2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1146) );
XOR2_X1 U826 ( .A(n1147), .B(KEYINPUT26), .Z(n1144) );
NAND2_X1 U827 ( .A1(KEYINPUT60), .A2(n1136), .ZN(n1131) );
NAND2_X1 U828 ( .A1(n1115), .A2(G472), .ZN(n1136) );
NOR2_X1 U829 ( .A1(n1107), .A2(n1148), .ZN(G54) );
XOR2_X1 U830 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U831 ( .A1(n1151), .A2(n1110), .ZN(n1150) );
NOR2_X1 U832 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
XOR2_X1 U833 ( .A(KEYINPUT11), .B(n1154), .Z(n1153) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
AND2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
XNOR2_X1 U836 ( .A(n1145), .B(n1157), .ZN(n1156) );
NOR2_X1 U837 ( .A1(n1107), .A2(n1158), .ZN(G51) );
XOR2_X1 U838 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U839 ( .A(n1161), .B(n1162), .Z(n1159) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1110), .ZN(n1162) );
INV_X1 U841 ( .A(n1115), .ZN(n1110) );
NOR2_X1 U842 ( .A1(n1164), .A2(n1017), .ZN(n1115) );
NOR2_X1 U843 ( .A1(n1101), .A2(n1090), .ZN(n1017) );
NAND4_X1 U844 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1090) );
NOR4_X1 U845 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
NOR3_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1167) );
NOR4_X1 U847 ( .A1(n1176), .A2(n1177), .A3(n1056), .A4(n1178), .ZN(n1175) );
NAND2_X1 U848 ( .A1(n1179), .A2(n1127), .ZN(n1177) );
INV_X1 U849 ( .A(KEYINPUT21), .ZN(n1176) );
NOR2_X1 U850 ( .A1(KEYINPUT21), .A2(n1180), .ZN(n1174) );
NOR3_X1 U851 ( .A1(n1181), .A2(n1065), .A3(n1182), .ZN(n1173) );
XOR2_X1 U852 ( .A(KEYINPUT32), .B(n1183), .Z(n1181) );
NAND4_X1 U853 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1101) );
NOR3_X1 U854 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NOR3_X1 U855 ( .A1(n1015), .A2(n1057), .A3(n1014), .ZN(n1190) );
NOR2_X1 U856 ( .A1(n1183), .A2(n1191), .ZN(n1057) );
NOR4_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1022), .A4(n1194), .ZN(n1189) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
XOR2_X1 U859 ( .A(n1014), .B(KEYINPUT23), .Z(n1196) );
AND2_X1 U860 ( .A1(n1065), .A2(n1195), .ZN(n1192) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1188) );
XOR2_X1 U862 ( .A(n1065), .B(KEYINPUT3), .Z(n1197) );
XOR2_X1 U863 ( .A(KEYINPUT13), .B(n1199), .Z(n1164) );
XOR2_X1 U864 ( .A(n1200), .B(KEYINPUT2), .Z(n1163) );
NAND2_X1 U865 ( .A1(KEYINPUT52), .A2(n1201), .ZN(n1161) );
XOR2_X1 U866 ( .A(n1202), .B(n1203), .Z(n1201) );
NAND2_X1 U867 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
OR3_X1 U868 ( .A1(n1206), .A2(n1147), .A3(KEYINPUT58), .ZN(n1205) );
NAND2_X1 U869 ( .A1(n1207), .A2(KEYINPUT58), .ZN(n1204) );
NOR2_X1 U870 ( .A1(n1020), .A2(G952), .ZN(n1107) );
XOR2_X1 U871 ( .A(G146), .B(n1172), .Z(G48) );
AND2_X1 U872 ( .A1(n1208), .A2(n1183), .ZN(n1172) );
XOR2_X1 U873 ( .A(n1209), .B(n1165), .Z(G45) );
NAND4_X1 U874 ( .A1(n1210), .A2(n1211), .A3(n1125), .A4(n1212), .ZN(n1165) );
XOR2_X1 U875 ( .A(G140), .B(n1171), .Z(G42) );
NOR3_X1 U876 ( .A1(n1127), .A2(n1064), .A3(n1182), .ZN(n1171) );
XOR2_X1 U877 ( .A(G137), .B(n1170), .Z(G39) );
AND4_X1 U878 ( .A1(n1213), .A2(n1051), .A3(n1040), .A4(n1214), .ZN(n1170) );
NAND2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(G36) );
NAND2_X1 U880 ( .A1(G134), .A2(n1166), .ZN(n1216) );
XOR2_X1 U881 ( .A(KEYINPUT9), .B(n1217), .Z(n1215) );
NOR2_X1 U882 ( .A1(G134), .A2(n1166), .ZN(n1217) );
NAND3_X1 U883 ( .A1(n1213), .A2(n1195), .A3(n1210), .ZN(n1166) );
XOR2_X1 U884 ( .A(G131), .B(n1218), .Z(G33) );
AND2_X1 U885 ( .A1(n1219), .A2(n1213), .ZN(n1218) );
INV_X1 U886 ( .A(n1182), .ZN(n1213) );
NAND4_X1 U887 ( .A1(n1041), .A2(n1125), .A3(n1220), .A4(n1048), .ZN(n1182) );
XOR2_X1 U888 ( .A(n1169), .B(n1221), .Z(G30) );
NOR2_X1 U889 ( .A1(KEYINPUT16), .A2(n1222), .ZN(n1221) );
AND2_X1 U890 ( .A1(n1208), .A2(n1191), .ZN(n1169) );
INV_X1 U891 ( .A(n1016), .ZN(n1191) );
NAND2_X1 U892 ( .A1(n1195), .A2(n1223), .ZN(n1016) );
NOR4_X1 U893 ( .A1(n1224), .A2(n1178), .A3(n1053), .A4(n1225), .ZN(n1208) );
XOR2_X1 U894 ( .A(G101), .B(n1226), .Z(G3) );
NOR2_X1 U895 ( .A1(n1198), .A2(n1065), .ZN(n1226) );
XOR2_X1 U896 ( .A(n1180), .B(n1227), .Z(G27) );
XNOR2_X1 U897 ( .A(KEYINPUT37), .B(n1206), .ZN(n1227) );
INV_X1 U898 ( .A(G125), .ZN(n1206) );
NAND4_X1 U899 ( .A1(n1211), .A2(n1183), .A3(n1059), .A4(n1179), .ZN(n1180) );
INV_X1 U900 ( .A(n1064), .ZN(n1179) );
INV_X1 U901 ( .A(n1127), .ZN(n1183) );
INV_X1 U902 ( .A(n1178), .ZN(n1211) );
NAND2_X1 U903 ( .A1(n1066), .A2(n1220), .ZN(n1178) );
NAND2_X1 U904 ( .A1(n1067), .A2(n1228), .ZN(n1220) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1076), .ZN(n1228) );
INV_X1 U906 ( .A(G900), .ZN(n1076) );
XOR2_X1 U907 ( .A(n1230), .B(n1231), .Z(G24) );
NAND4_X1 U908 ( .A1(n1232), .A2(n1046), .A3(n1223), .A4(n1212), .ZN(n1231) );
INV_X1 U909 ( .A(n1014), .ZN(n1046) );
NAND2_X1 U910 ( .A1(n1233), .A2(n1225), .ZN(n1014) );
XOR2_X1 U911 ( .A(n1040), .B(KEYINPUT31), .Z(n1233) );
XNOR2_X1 U912 ( .A(n1186), .B(n1234), .ZN(G21) );
NOR2_X1 U913 ( .A1(KEYINPUT4), .A2(n1235), .ZN(n1234) );
NAND4_X1 U914 ( .A1(n1232), .A2(n1051), .A3(n1040), .A4(n1214), .ZN(n1186) );
NAND2_X1 U915 ( .A1(n1236), .A2(n1237), .ZN(G18) );
NAND2_X1 U916 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U917 ( .A1(n1240), .A2(G116), .ZN(n1236) );
NAND2_X1 U918 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U919 ( .A1(KEYINPUT0), .A2(n1243), .ZN(n1242) );
OR2_X1 U920 ( .A1(n1238), .A2(KEYINPUT0), .ZN(n1241) );
AND2_X1 U921 ( .A1(KEYINPUT20), .A2(n1243), .ZN(n1238) );
AND3_X1 U922 ( .A1(n1244), .A2(n1210), .A3(n1245), .ZN(n1243) );
AND3_X1 U923 ( .A1(n1066), .A2(n1124), .A3(n1195), .ZN(n1245) );
INV_X1 U924 ( .A(n1212), .ZN(n1195) );
NOR2_X1 U925 ( .A1(n1065), .A2(n1022), .ZN(n1210) );
XOR2_X1 U926 ( .A(n1056), .B(KEYINPUT57), .Z(n1244) );
XOR2_X1 U927 ( .A(n1246), .B(n1184), .Z(G15) );
NAND2_X1 U928 ( .A1(n1232), .A2(n1219), .ZN(n1184) );
NOR2_X1 U929 ( .A1(n1127), .A2(n1065), .ZN(n1219) );
NAND2_X1 U930 ( .A1(n1225), .A2(n1040), .ZN(n1065) );
INV_X1 U931 ( .A(n1214), .ZN(n1225) );
NAND2_X1 U932 ( .A1(n1022), .A2(n1212), .ZN(n1127) );
INV_X1 U933 ( .A(n1194), .ZN(n1232) );
NAND3_X1 U934 ( .A1(n1066), .A2(n1124), .A3(n1059), .ZN(n1194) );
INV_X1 U935 ( .A(n1056), .ZN(n1059) );
NAND3_X1 U936 ( .A1(n1247), .A2(n1029), .A3(n1055), .ZN(n1056) );
XNOR2_X1 U937 ( .A(G110), .B(n1185), .ZN(G12) );
OR2_X1 U938 ( .A1(n1064), .A2(n1198), .ZN(n1185) );
NAND2_X1 U939 ( .A1(n1051), .A2(n1248), .ZN(n1198) );
INV_X1 U940 ( .A(n1015), .ZN(n1248) );
NAND3_X1 U941 ( .A1(n1066), .A2(n1124), .A3(n1125), .ZN(n1015) );
INV_X1 U942 ( .A(n1053), .ZN(n1125) );
NAND2_X1 U943 ( .A1(n1247), .A2(n1249), .ZN(n1053) );
NAND2_X1 U944 ( .A1(n1055), .A2(n1029), .ZN(n1249) );
NAND3_X1 U945 ( .A1(n1151), .A2(n1199), .A3(n1250), .ZN(n1029) );
INV_X1 U946 ( .A(G469), .ZN(n1151) );
XOR2_X1 U947 ( .A(n1032), .B(KEYINPUT61), .Z(n1055) );
NAND2_X1 U948 ( .A1(G469), .A2(n1251), .ZN(n1032) );
NAND2_X1 U949 ( .A1(n1250), .A2(n1199), .ZN(n1251) );
XOR2_X1 U950 ( .A(n1155), .B(n1252), .Z(n1250) );
XOR2_X1 U951 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U952 ( .A1(KEYINPUT7), .A2(n1157), .ZN(n1254) );
XNOR2_X1 U953 ( .A(n1255), .B(n1077), .ZN(n1157) );
XNOR2_X1 U954 ( .A(n1222), .B(n1256), .ZN(n1077) );
NOR2_X1 U955 ( .A1(KEYINPUT54), .A2(n1257), .ZN(n1256) );
XOR2_X1 U956 ( .A(n1209), .B(n1258), .Z(n1257) );
INV_X1 U957 ( .A(G143), .ZN(n1209) );
XOR2_X1 U958 ( .A(n1259), .B(n1260), .Z(n1255) );
NOR3_X1 U959 ( .A1(n1261), .A2(KEYINPUT5), .A3(n1262), .ZN(n1260) );
NOR2_X1 U960 ( .A1(G104), .A2(n1263), .ZN(n1262) );
XOR2_X1 U961 ( .A(KEYINPUT53), .B(n1264), .Z(n1261) );
AND2_X1 U962 ( .A1(n1263), .A2(G104), .ZN(n1264) );
INV_X1 U963 ( .A(G107), .ZN(n1263) );
XNOR2_X1 U964 ( .A(n1265), .B(n1266), .ZN(n1155) );
XOR2_X1 U965 ( .A(G140), .B(G110), .Z(n1266) );
NAND2_X1 U966 ( .A1(G227), .A2(n1020), .ZN(n1265) );
XOR2_X1 U967 ( .A(n1028), .B(KEYINPUT49), .Z(n1247) );
AND2_X1 U968 ( .A1(G221), .A2(n1267), .ZN(n1028) );
XOR2_X1 U969 ( .A(KEYINPUT47), .B(n1268), .Z(n1267) );
AND2_X1 U970 ( .A1(n1199), .A2(G234), .ZN(n1268) );
NAND2_X1 U971 ( .A1(n1067), .A2(n1269), .ZN(n1124) );
NAND4_X1 U972 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1270), .ZN(n1269) );
INV_X1 U973 ( .A(G898), .ZN(n1270) );
NAND3_X1 U974 ( .A1(n1229), .A2(n1020), .A3(G952), .ZN(n1067) );
NAND2_X1 U975 ( .A1(G234), .A2(G237), .ZN(n1229) );
NOR2_X1 U976 ( .A1(n1041), .A2(n1026), .ZN(n1066) );
INV_X1 U977 ( .A(n1048), .ZN(n1026) );
NAND2_X1 U978 ( .A1(G214), .A2(n1271), .ZN(n1048) );
XNOR2_X1 U979 ( .A(n1272), .B(n1200), .ZN(n1041) );
NAND2_X1 U980 ( .A1(G210), .A2(n1271), .ZN(n1200) );
NAND2_X1 U981 ( .A1(n1273), .A2(n1199), .ZN(n1271) );
NAND2_X1 U982 ( .A1(n1274), .A2(n1199), .ZN(n1272) );
XOR2_X1 U983 ( .A(n1160), .B(n1275), .Z(n1274) );
XOR2_X1 U984 ( .A(n1203), .B(n1207), .Z(n1275) );
XNOR2_X1 U985 ( .A(G125), .B(n1147), .ZN(n1207) );
NOR2_X1 U986 ( .A1(n1097), .A2(G953), .ZN(n1203) );
INV_X1 U987 ( .A(G224), .ZN(n1097) );
XNOR2_X1 U988 ( .A(n1102), .B(KEYINPUT27), .ZN(n1160) );
XOR2_X1 U989 ( .A(n1276), .B(n1277), .Z(n1102) );
XOR2_X1 U990 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U991 ( .A(n1280), .B(n1281), .Z(n1279) );
NOR2_X1 U992 ( .A1(G104), .A2(KEYINPUT43), .ZN(n1281) );
NAND3_X1 U993 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1280) );
NAND2_X1 U994 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
INV_X1 U995 ( .A(n1287), .ZN(n1286) );
NAND3_X1 U996 ( .A1(n1287), .A2(n1239), .A3(n1235), .ZN(n1283) );
INV_X1 U997 ( .A(G119), .ZN(n1235) );
NAND2_X1 U998 ( .A1(n1288), .A2(G119), .ZN(n1282) );
XOR2_X1 U999 ( .A(n1239), .B(n1287), .Z(n1288) );
NOR2_X1 U1000 ( .A1(KEYINPUT63), .A2(G113), .ZN(n1287) );
NAND2_X1 U1001 ( .A1(KEYINPUT18), .A2(n1230), .ZN(n1278) );
INV_X1 U1002 ( .A(G122), .ZN(n1230) );
XOR2_X1 U1003 ( .A(n1259), .B(n1289), .Z(n1276) );
XOR2_X1 U1004 ( .A(G110), .B(G107), .Z(n1289) );
INV_X1 U1005 ( .A(G101), .ZN(n1259) );
NOR2_X1 U1006 ( .A1(n1223), .A2(n1212), .ZN(n1051) );
NAND2_X1 U1007 ( .A1(n1290), .A2(n1030), .ZN(n1212) );
NAND2_X1 U1008 ( .A1(n1038), .A2(n1120), .ZN(n1030) );
INV_X1 U1009 ( .A(G475), .ZN(n1120) );
INV_X1 U1010 ( .A(n1291), .ZN(n1038) );
NAND2_X1 U1011 ( .A1(G475), .A2(n1291), .ZN(n1290) );
NAND2_X1 U1012 ( .A1(n1121), .A2(n1199), .ZN(n1291) );
XNOR2_X1 U1013 ( .A(n1292), .B(n1293), .ZN(n1121) );
XOR2_X1 U1014 ( .A(G122), .B(G113), .Z(n1293) );
XNOR2_X1 U1015 ( .A(n1294), .B(n1295), .ZN(n1292) );
NOR2_X1 U1016 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1295) );
NOR2_X1 U1017 ( .A1(KEYINPUT51), .A2(n1296), .ZN(n1294) );
XOR2_X1 U1018 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1019 ( .A(n1089), .B(n1258), .Z(n1298) );
XOR2_X1 U1020 ( .A(n1299), .B(n1300), .Z(n1297) );
NOR2_X1 U1021 ( .A1(G143), .A2(KEYINPUT40), .ZN(n1300) );
XOR2_X1 U1022 ( .A(n1301), .B(G131), .Z(n1299) );
NAND3_X1 U1023 ( .A1(G214), .A2(n1020), .A3(n1302), .ZN(n1301) );
XOR2_X1 U1024 ( .A(n1273), .B(KEYINPUT24), .Z(n1302) );
INV_X1 U1025 ( .A(n1022), .ZN(n1223) );
XOR2_X1 U1026 ( .A(n1303), .B(G478), .Z(n1022) );
NAND2_X1 U1027 ( .A1(n1116), .A2(n1199), .ZN(n1303) );
XNOR2_X1 U1028 ( .A(n1304), .B(n1305), .ZN(n1116) );
XOR2_X1 U1029 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1030 ( .A(G128), .B(G122), .Z(n1307) );
XOR2_X1 U1031 ( .A(G143), .B(G134), .Z(n1306) );
XOR2_X1 U1032 ( .A(n1308), .B(n1309), .Z(n1304) );
XOR2_X1 U1033 ( .A(G116), .B(G107), .Z(n1309) );
NAND3_X1 U1034 ( .A1(G217), .A2(n1020), .A3(G234), .ZN(n1308) );
NAND2_X1 U1035 ( .A1(n1224), .A2(n1214), .ZN(n1064) );
NAND2_X1 U1036 ( .A1(n1310), .A2(n1311), .ZN(n1214) );
OR2_X1 U1037 ( .A1(n1037), .A2(n1036), .ZN(n1311) );
XOR2_X1 U1038 ( .A(n1031), .B(KEYINPUT50), .Z(n1310) );
NAND2_X1 U1039 ( .A1(n1036), .A2(n1037), .ZN(n1031) );
NAND2_X1 U1040 ( .A1(G217), .A2(n1312), .ZN(n1037) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1199), .ZN(n1312) );
NOR2_X1 U1042 ( .A1(n1109), .A2(G902), .ZN(n1036) );
XNOR2_X1 U1043 ( .A(n1313), .B(n1314), .ZN(n1109) );
XOR2_X1 U1044 ( .A(G110), .B(n1315), .Z(n1314) );
XOR2_X1 U1045 ( .A(G137), .B(G119), .Z(n1315) );
XOR2_X1 U1046 ( .A(n1316), .B(n1317), .Z(n1313) );
XOR2_X1 U1047 ( .A(n1318), .B(n1319), .Z(n1316) );
NOR2_X1 U1048 ( .A1(KEYINPUT55), .A2(n1089), .ZN(n1319) );
XNOR2_X1 U1049 ( .A(G140), .B(G125), .ZN(n1089) );
NAND3_X1 U1050 ( .A1(G234), .A2(n1020), .A3(G221), .ZN(n1318) );
INV_X1 U1051 ( .A(n1040), .ZN(n1224) );
XOR2_X1 U1052 ( .A(n1320), .B(n1321), .Z(n1040) );
XOR2_X1 U1053 ( .A(KEYINPUT17), .B(G472), .Z(n1321) );
NAND2_X1 U1054 ( .A1(n1322), .A2(n1199), .ZN(n1320) );
INV_X1 U1055 ( .A(G902), .ZN(n1199) );
XOR2_X1 U1056 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1057 ( .A(n1253), .B(n1130), .Z(n1324) );
XNOR2_X1 U1058 ( .A(n1325), .B(G101), .ZN(n1130) );
NAND3_X1 U1059 ( .A1(n1273), .A2(n1020), .A3(G210), .ZN(n1325) );
INV_X1 U1060 ( .A(G953), .ZN(n1020) );
INV_X1 U1061 ( .A(G237), .ZN(n1273) );
INV_X1 U1062 ( .A(n1145), .ZN(n1253) );
XNOR2_X1 U1063 ( .A(n1087), .B(n1326), .ZN(n1145) );
NOR2_X1 U1064 ( .A1(G131), .A2(KEYINPUT56), .ZN(n1326) );
XOR2_X1 U1065 ( .A(G134), .B(G137), .Z(n1087) );
XOR2_X1 U1066 ( .A(n1139), .B(n1147), .Z(n1323) );
XNOR2_X1 U1067 ( .A(n1317), .B(n1327), .ZN(n1147) );
NOR2_X1 U1068 ( .A1(KEYINPUT46), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1069 ( .A(KEYINPUT45), .B(G143), .Z(n1328) );
XNOR2_X1 U1070 ( .A(n1222), .B(n1258), .ZN(n1317) );
XOR2_X1 U1071 ( .A(G146), .B(KEYINPUT19), .Z(n1258) );
INV_X1 U1072 ( .A(G128), .ZN(n1222) );
NAND2_X1 U1073 ( .A1(n1329), .A2(n1330), .ZN(n1139) );
OR3_X1 U1074 ( .A1(n1285), .A2(G113), .A3(n1331), .ZN(n1330) );
XOR2_X1 U1075 ( .A(KEYINPUT34), .B(n1332), .Z(n1329) );
NOR2_X1 U1076 ( .A1(n1333), .A2(n1246), .ZN(n1332) );
INV_X1 U1077 ( .A(G113), .ZN(n1246) );
NOR2_X1 U1078 ( .A1(n1285), .A2(n1331), .ZN(n1333) );
XNOR2_X1 U1079 ( .A(n1334), .B(KEYINPUT36), .ZN(n1331) );
NAND2_X1 U1080 ( .A1(G119), .A2(n1239), .ZN(n1334) );
NOR2_X1 U1081 ( .A1(n1239), .A2(G119), .ZN(n1285) );
INV_X1 U1082 ( .A(G116), .ZN(n1239) );
endmodule


