//Key = 0010000110001110010001111101010111001110101001000011100011000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333;

XNOR2_X1 U731 ( .A(G107), .B(n1009), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1012), .A2(n1013), .A3(G953), .A4(n1014), .ZN(n1011) );
NOR3_X1 U734 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1013) );
INV_X1 U735 ( .A(n1018), .ZN(n1017) );
NOR2_X1 U736 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NOR2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
INV_X1 U738 ( .A(n1023), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NOR2_X1 U740 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U742 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR3_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1024) );
AND3_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1019) );
NAND2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1012) );
NAND2_X1 U746 ( .A1(n1035), .A2(n1040), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1023), .ZN(n1042) );
NAND2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1047), .ZN(n1046) );
NAND2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
INV_X1 U753 ( .A(n1052), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1018), .A2(n1053), .ZN(n1045) );
XOR2_X1 U755 ( .A(n1054), .B(KEYINPUT58), .Z(n1041) );
NAND4_X1 U756 ( .A1(n1055), .A2(n1043), .A3(n1037), .A4(n1018), .ZN(n1054) );
NOR3_X1 U757 ( .A1(n1014), .A2(G953), .A3(G952), .ZN(n1010) );
AND4_X1 U758 ( .A1(n1050), .A2(n1056), .A3(n1037), .A4(n1057), .ZN(n1014) );
NOR4_X1 U759 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
XOR2_X1 U760 ( .A(n1062), .B(n1063), .Z(n1061) );
NOR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XNOR2_X1 U762 ( .A(KEYINPUT61), .B(KEYINPUT25), .ZN(n1065) );
XNOR2_X1 U763 ( .A(G478), .B(n1066), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1067), .A2(KEYINPUT6), .ZN(n1066) );
XNOR2_X1 U765 ( .A(n1068), .B(n1069), .ZN(n1059) );
NAND2_X1 U766 ( .A1(KEYINPUT33), .A2(n1070), .ZN(n1068) );
XOR2_X1 U767 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U769 ( .A(n1075), .ZN(n1074) );
AND2_X1 U770 ( .A1(G227), .A2(G900), .ZN(n1073) );
NOR2_X1 U771 ( .A1(KEYINPUT10), .A2(n1076), .ZN(n1071) );
XOR2_X1 U772 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U775 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(n1081) );
XNOR2_X1 U777 ( .A(KEYINPUT49), .B(n1087), .ZN(n1086) );
NOR2_X1 U778 ( .A1(KEYINPUT44), .A2(n1088), .ZN(n1087) );
XNOR2_X1 U779 ( .A(KEYINPUT54), .B(n1089), .ZN(n1088) );
INV_X1 U780 ( .A(G134), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1085) );
NAND2_X1 U782 ( .A1(G140), .A2(n1092), .ZN(n1091) );
XOR2_X1 U783 ( .A(KEYINPUT56), .B(n1093), .Z(n1090) );
NOR2_X1 U784 ( .A1(G140), .A2(n1092), .ZN(n1093) );
NOR2_X1 U785 ( .A1(G900), .A2(n1094), .ZN(n1079) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1077) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(G69) );
NAND2_X1 U788 ( .A1(n1075), .A2(n1098), .ZN(n1097) );
NAND2_X1 U789 ( .A1(G898), .A2(G224), .ZN(n1098) );
XOR2_X1 U790 ( .A(G953), .B(KEYINPUT43), .Z(n1075) );
NAND2_X1 U791 ( .A1(KEYINPUT40), .A2(n1099), .ZN(n1096) );
XOR2_X1 U792 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U793 ( .A1(n1094), .A2(n1102), .ZN(n1101) );
NAND2_X1 U794 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U795 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1103) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1106) );
NAND2_X1 U798 ( .A1(KEYINPUT51), .A2(n1110), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(G66) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1114) );
AND2_X1 U802 ( .A1(n1117), .A2(KEYINPUT63), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NOR2_X1 U804 ( .A1(KEYINPUT63), .A2(n1117), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1120), .ZN(G63) );
NOR3_X1 U806 ( .A1(n1067), .A2(n1121), .A3(n1122), .ZN(n1120) );
AND3_X1 U807 ( .A1(n1123), .A2(G478), .A3(n1118), .ZN(n1122) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1123), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1038), .A2(n1125), .ZN(n1124) );
NOR3_X1 U810 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(G60) );
AND3_X1 U811 ( .A1(KEYINPUT35), .A2(G953), .A3(G952), .ZN(n1128) );
NOR2_X1 U812 ( .A1(KEYINPUT35), .A2(n1129), .ZN(n1127) );
INV_X1 U813 ( .A(n1111), .ZN(n1129) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1126) );
NAND2_X1 U815 ( .A1(n1118), .A2(G475), .ZN(n1130) );
XNOR2_X1 U816 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1111), .A2(n1133), .ZN(G57) );
XOR2_X1 U818 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U819 ( .A(G101), .B(n1136), .ZN(n1135) );
NAND2_X1 U820 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND2_X1 U821 ( .A1(KEYINPUT20), .A2(n1139), .ZN(n1138) );
XOR2_X1 U822 ( .A(n1140), .B(n1141), .Z(n1137) );
NOR2_X1 U823 ( .A1(KEYINPUT20), .A2(n1139), .ZN(n1141) );
NAND3_X1 U824 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1139) );
NAND2_X1 U825 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
INV_X1 U826 ( .A(KEYINPUT57), .ZN(n1146) );
NAND3_X1 U827 ( .A1(KEYINPUT57), .A2(n1147), .A3(n1148), .ZN(n1143) );
OR2_X1 U828 ( .A1(n1148), .A2(n1147), .ZN(n1142) );
NOR2_X1 U829 ( .A1(KEYINPUT60), .A2(n1145), .ZN(n1147) );
XNOR2_X1 U830 ( .A(n1149), .B(n1150), .ZN(n1145) );
NAND2_X1 U831 ( .A1(KEYINPUT21), .A2(n1151), .ZN(n1149) );
NAND2_X1 U832 ( .A1(n1118), .A2(G472), .ZN(n1140) );
NOR2_X1 U833 ( .A1(n1111), .A2(n1152), .ZN(G54) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U835 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND3_X1 U836 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
OR2_X1 U837 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND3_X1 U838 ( .A1(n1161), .A2(n1160), .A3(n1162), .ZN(n1158) );
NAND2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1157) );
NAND2_X1 U840 ( .A1(n1165), .A2(n1160), .ZN(n1164) );
INV_X1 U841 ( .A(KEYINPUT4), .ZN(n1160) );
XNOR2_X1 U842 ( .A(n1161), .B(KEYINPUT36), .ZN(n1165) );
XNOR2_X1 U843 ( .A(n1166), .B(KEYINPUT55), .ZN(n1161) );
INV_X1 U844 ( .A(n1162), .ZN(n1163) );
NAND3_X1 U845 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1155) );
NAND2_X1 U846 ( .A1(KEYINPUT0), .A2(n1170), .ZN(n1169) );
INV_X1 U847 ( .A(n1171), .ZN(n1170) );
OR3_X1 U848 ( .A1(n1172), .A2(KEYINPUT0), .A3(n1150), .ZN(n1168) );
NAND2_X1 U849 ( .A1(n1150), .A2(n1172), .ZN(n1167) );
NAND2_X1 U850 ( .A1(KEYINPUT13), .A2(n1171), .ZN(n1172) );
XOR2_X1 U851 ( .A(G101), .B(n1173), .Z(n1171) );
NAND2_X1 U852 ( .A1(n1118), .A2(G469), .ZN(n1153) );
NOR2_X1 U853 ( .A1(n1111), .A2(n1174), .ZN(G51) );
XOR2_X1 U854 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U855 ( .A1(n1118), .A2(n1064), .ZN(n1176) );
NOR2_X1 U856 ( .A1(n1177), .A2(n1038), .ZN(n1118) );
NOR2_X1 U857 ( .A1(n1095), .A2(n1102), .ZN(n1038) );
NAND4_X1 U858 ( .A1(n1132), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1102) );
AND4_X1 U859 ( .A1(n1009), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1180) );
NAND3_X1 U860 ( .A1(n1036), .A2(n1018), .A3(n1184), .ZN(n1009) );
NAND2_X1 U861 ( .A1(n1029), .A2(n1185), .ZN(n1179) );
NAND2_X1 U862 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U863 ( .A(n1188), .B(KEYINPUT59), .Z(n1186) );
NAND3_X1 U864 ( .A1(n1184), .A2(n1018), .A3(n1055), .ZN(n1132) );
NAND4_X1 U865 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1095) );
NOR4_X1 U866 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
INV_X1 U867 ( .A(n1197), .ZN(n1196) );
NAND2_X1 U868 ( .A1(n1053), .A2(n1198), .ZN(n1191) );
NAND2_X1 U869 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND4_X1 U870 ( .A1(n1035), .A2(n1052), .A3(n1036), .A4(n1201), .ZN(n1200) );
NAND2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
XNOR2_X1 U872 ( .A(n1035), .B(KEYINPUT8), .ZN(n1202) );
NAND3_X1 U873 ( .A1(n1037), .A2(n1029), .A3(n1203), .ZN(n1189) );
INV_X1 U874 ( .A(n1204), .ZN(n1203) );
NAND3_X1 U875 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1175) );
OR2_X1 U876 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND3_X1 U877 ( .A1(n1209), .A2(n1208), .A3(n1210), .ZN(n1206) );
NAND2_X1 U878 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND2_X1 U879 ( .A1(n1213), .A2(n1208), .ZN(n1212) );
INV_X1 U880 ( .A(KEYINPUT41), .ZN(n1208) );
XNOR2_X1 U881 ( .A(KEYINPUT7), .B(n1209), .ZN(n1213) );
NAND2_X1 U882 ( .A1(n1214), .A2(n1215), .ZN(n1209) );
NAND2_X1 U883 ( .A1(n1216), .A2(n1092), .ZN(n1215) );
XOR2_X1 U884 ( .A(KEYINPUT32), .B(n1217), .Z(n1216) );
NAND2_X1 U885 ( .A1(n1217), .A2(G125), .ZN(n1214) );
NOR2_X1 U886 ( .A1(n1094), .A2(G952), .ZN(n1111) );
XNOR2_X1 U887 ( .A(G146), .B(n1190), .ZN(G48) );
NAND3_X1 U888 ( .A1(n1218), .A2(n1029), .A3(n1055), .ZN(n1190) );
XNOR2_X1 U889 ( .A(G143), .B(n1197), .ZN(G45) );
NAND4_X1 U890 ( .A1(n1219), .A2(n1220), .A3(n1029), .A4(n1221), .ZN(n1197) );
XOR2_X1 U891 ( .A(G140), .B(n1222), .Z(G42) );
NOR3_X1 U892 ( .A1(n1204), .A2(n1223), .A3(n1033), .ZN(n1222) );
INV_X1 U893 ( .A(n1035), .ZN(n1033) );
XNOR2_X1 U894 ( .A(G137), .B(n1224), .ZN(G39) );
NAND2_X1 U895 ( .A1(KEYINPUT23), .A2(n1195), .ZN(n1224) );
AND3_X1 U896 ( .A1(n1035), .A2(n1218), .A3(n1023), .ZN(n1195) );
XNOR2_X1 U897 ( .A(G134), .B(n1225), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1220), .A2(n1036), .A3(n1226), .ZN(n1225) );
XNOR2_X1 U899 ( .A(n1035), .B(KEYINPUT42), .ZN(n1226) );
XOR2_X1 U900 ( .A(G131), .B(n1194), .Z(G33) );
AND3_X1 U901 ( .A1(n1055), .A2(n1220), .A3(n1035), .ZN(n1194) );
NOR2_X1 U902 ( .A1(n1030), .A2(n1058), .ZN(n1035) );
AND3_X1 U903 ( .A1(n1053), .A2(n1201), .A3(n1052), .ZN(n1220) );
XNOR2_X1 U904 ( .A(n1227), .B(n1193), .ZN(G30) );
AND3_X1 U905 ( .A1(n1036), .A2(n1029), .A3(n1218), .ZN(n1193) );
AND4_X1 U906 ( .A1(n1053), .A2(n1051), .A3(n1228), .A4(n1201), .ZN(n1218) );
XNOR2_X1 U907 ( .A(G101), .B(n1178), .ZN(G3) );
NAND3_X1 U908 ( .A1(n1052), .A2(n1184), .A3(n1023), .ZN(n1178) );
XNOR2_X1 U909 ( .A(n1092), .B(n1229), .ZN(G27) );
NOR3_X1 U910 ( .A1(n1204), .A2(n1230), .A3(n1027), .ZN(n1229) );
XNOR2_X1 U911 ( .A(n1029), .B(KEYINPUT53), .ZN(n1230) );
NAND4_X1 U912 ( .A1(n1050), .A2(n1055), .A3(n1051), .A4(n1201), .ZN(n1204) );
NAND2_X1 U913 ( .A1(n1231), .A2(n1232), .ZN(n1201) );
NAND4_X1 U914 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1234), .ZN(n1232) );
INV_X1 U915 ( .A(G900), .ZN(n1234) );
XNOR2_X1 U916 ( .A(n1043), .B(KEYINPUT18), .ZN(n1231) );
INV_X1 U917 ( .A(n1015), .ZN(n1043) );
XNOR2_X1 U918 ( .A(n1235), .B(n1236), .ZN(G24) );
NOR2_X1 U919 ( .A1(n1237), .A2(n1188), .ZN(n1236) );
NAND4_X1 U920 ( .A1(n1238), .A2(n1018), .A3(n1219), .A4(n1221), .ZN(n1188) );
NOR2_X1 U921 ( .A1(n1228), .A2(n1051), .ZN(n1018) );
INV_X1 U922 ( .A(n1029), .ZN(n1237) );
XNOR2_X1 U923 ( .A(G119), .B(n1183), .ZN(G21) );
NAND3_X1 U924 ( .A1(n1238), .A2(n1023), .A3(n1239), .ZN(n1183) );
AND3_X1 U925 ( .A1(n1029), .A2(n1228), .A3(n1051), .ZN(n1239) );
NAND2_X1 U926 ( .A1(n1240), .A2(n1241), .ZN(G18) );
NAND2_X1 U927 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U928 ( .A1(G116), .A2(n1244), .ZN(n1240) );
NAND2_X1 U929 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
OR2_X1 U930 ( .A1(n1182), .A2(KEYINPUT52), .ZN(n1246) );
NAND2_X1 U931 ( .A1(KEYINPUT52), .A2(n1247), .ZN(n1245) );
INV_X1 U932 ( .A(n1242), .ZN(n1247) );
NOR2_X1 U933 ( .A1(KEYINPUT1), .A2(n1182), .ZN(n1242) );
NAND4_X1 U934 ( .A1(n1238), .A2(n1052), .A3(n1036), .A4(n1029), .ZN(n1182) );
NOR2_X1 U935 ( .A1(n1221), .A2(n1248), .ZN(n1036) );
NAND2_X1 U936 ( .A1(n1249), .A2(n1250), .ZN(G15) );
OR2_X1 U937 ( .A1(n1251), .A2(G113), .ZN(n1250) );
XOR2_X1 U938 ( .A(n1252), .B(KEYINPUT47), .Z(n1249) );
NAND2_X1 U939 ( .A1(G113), .A2(n1251), .ZN(n1252) );
NAND2_X1 U940 ( .A1(n1029), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U941 ( .A(KEYINPUT5), .B(n1187), .ZN(n1253) );
NAND3_X1 U942 ( .A1(n1055), .A2(n1052), .A3(n1238), .ZN(n1187) );
AND2_X1 U943 ( .A1(n1037), .A2(n1254), .ZN(n1238) );
INV_X1 U944 ( .A(n1027), .ZN(n1037) );
NAND2_X1 U945 ( .A1(n1255), .A2(n1032), .ZN(n1027) );
INV_X1 U946 ( .A(n1034), .ZN(n1255) );
NOR2_X1 U947 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
AND2_X1 U948 ( .A1(n1256), .A2(n1221), .ZN(n1055) );
XNOR2_X1 U949 ( .A(n1248), .B(KEYINPUT24), .ZN(n1256) );
XNOR2_X1 U950 ( .A(G110), .B(n1181), .ZN(G12) );
NAND4_X1 U951 ( .A1(n1023), .A2(n1184), .A3(n1050), .A4(n1051), .ZN(n1181) );
XNOR2_X1 U952 ( .A(n1056), .B(KEYINPUT19), .ZN(n1051) );
XOR2_X1 U953 ( .A(n1257), .B(n1119), .Z(n1056) );
AND2_X1 U954 ( .A1(G217), .A2(n1258), .ZN(n1119) );
OR2_X1 U955 ( .A1(n1117), .A2(G902), .ZN(n1257) );
XNOR2_X1 U956 ( .A(n1259), .B(n1260), .ZN(n1117) );
XNOR2_X1 U957 ( .A(n1261), .B(n1262), .ZN(n1260) );
NAND2_X1 U958 ( .A1(KEYINPUT45), .A2(n1263), .ZN(n1261) );
XOR2_X1 U959 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U960 ( .A(n1227), .B(G119), .ZN(n1265) );
XOR2_X1 U961 ( .A(n1266), .B(n1267), .Z(n1259) );
XNOR2_X1 U962 ( .A(n1268), .B(G125), .ZN(n1267) );
INV_X1 U963 ( .A(G137), .ZN(n1268) );
NAND2_X1 U964 ( .A1(n1269), .A2(G221), .ZN(n1266) );
INV_X1 U965 ( .A(n1228), .ZN(n1050) );
XNOR2_X1 U966 ( .A(n1270), .B(G472), .ZN(n1228) );
NAND2_X1 U967 ( .A1(n1271), .A2(n1177), .ZN(n1270) );
XOR2_X1 U968 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U969 ( .A(n1274), .B(n1148), .ZN(n1273) );
XOR2_X1 U970 ( .A(n1275), .B(n1276), .Z(n1148) );
NOR2_X1 U971 ( .A1(KEYINPUT9), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U972 ( .A(G116), .B(G119), .ZN(n1275) );
XOR2_X1 U973 ( .A(n1136), .B(n1151), .Z(n1272) );
NAND3_X1 U974 ( .A1(G210), .A2(n1094), .A3(n1278), .ZN(n1136) );
AND3_X1 U975 ( .A1(n1053), .A2(n1254), .A3(n1029), .ZN(n1184) );
NOR2_X1 U976 ( .A1(n1279), .A2(n1058), .ZN(n1029) );
INV_X1 U977 ( .A(n1031), .ZN(n1058) );
NAND2_X1 U978 ( .A1(G214), .A2(n1280), .ZN(n1031) );
INV_X1 U979 ( .A(n1030), .ZN(n1279) );
XNOR2_X1 U980 ( .A(n1062), .B(n1064), .ZN(n1030) );
AND2_X1 U981 ( .A1(G210), .A2(n1280), .ZN(n1064) );
NAND2_X1 U982 ( .A1(n1281), .A2(n1177), .ZN(n1280) );
NAND2_X1 U983 ( .A1(n1282), .A2(n1177), .ZN(n1062) );
XNOR2_X1 U984 ( .A(n1283), .B(n1210), .ZN(n1282) );
INV_X1 U985 ( .A(n1211), .ZN(n1210) );
XNOR2_X1 U986 ( .A(n1284), .B(n1109), .ZN(n1211) );
XNOR2_X1 U987 ( .A(n1235), .B(n1264), .ZN(n1109) );
NAND2_X1 U988 ( .A1(n1285), .A2(KEYINPUT29), .ZN(n1284) );
XOR2_X1 U989 ( .A(n1110), .B(n1107), .Z(n1285) );
XNOR2_X1 U990 ( .A(n1286), .B(n1287), .ZN(n1107) );
NAND2_X1 U991 ( .A1(KEYINPUT12), .A2(G101), .ZN(n1286) );
XNOR2_X1 U992 ( .A(n1288), .B(n1277), .ZN(n1110) );
XOR2_X1 U993 ( .A(n1289), .B(G119), .Z(n1288) );
NAND2_X1 U994 ( .A1(KEYINPUT37), .A2(n1243), .ZN(n1289) );
INV_X1 U995 ( .A(G116), .ZN(n1243) );
NAND2_X1 U996 ( .A1(KEYINPUT31), .A2(n1290), .ZN(n1283) );
XOR2_X1 U997 ( .A(n1291), .B(n1292), .Z(n1290) );
XNOR2_X1 U998 ( .A(n1092), .B(n1217), .ZN(n1292) );
XNOR2_X1 U999 ( .A(n1293), .B(n1151), .ZN(n1217) );
XNOR2_X1 U1000 ( .A(n1294), .B(G128), .ZN(n1151) );
NAND3_X1 U1001 ( .A1(KEYINPUT27), .A2(n1295), .A3(n1296), .ZN(n1294) );
XNOR2_X1 U1002 ( .A(n1297), .B(KEYINPUT30), .ZN(n1296) );
NAND2_X1 U1003 ( .A1(G143), .A2(n1298), .ZN(n1295) );
NAND2_X1 U1004 ( .A1(G224), .A2(n1094), .ZN(n1293) );
INV_X1 U1005 ( .A(G125), .ZN(n1092) );
XOR2_X1 U1006 ( .A(KEYINPUT28), .B(KEYINPUT26), .Z(n1291) );
NAND2_X1 U1007 ( .A1(n1015), .A2(n1299), .ZN(n1254) );
NAND4_X1 U1008 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1105), .ZN(n1299) );
INV_X1 U1009 ( .A(G898), .ZN(n1105) );
NAND3_X1 U1010 ( .A1(n1233), .A2(n1094), .A3(G952), .ZN(n1015) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1233) );
INV_X1 U1012 ( .A(n1223), .ZN(n1053) );
NAND2_X1 U1013 ( .A1(n1034), .A2(n1032), .ZN(n1223) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1258), .ZN(n1032) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1177), .ZN(n1258) );
XNOR2_X1 U1016 ( .A(n1300), .B(G469), .ZN(n1034) );
NAND2_X1 U1017 ( .A1(n1301), .A2(n1177), .ZN(n1300) );
XOR2_X1 U1018 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1019 ( .A(n1166), .B(n1304), .ZN(n1303) );
NOR2_X1 U1020 ( .A1(KEYINPUT11), .A2(n1162), .ZN(n1304) );
XOR2_X1 U1021 ( .A(G140), .B(n1264), .Z(n1162) );
XOR2_X1 U1022 ( .A(G110), .B(KEYINPUT38), .Z(n1264) );
NAND2_X1 U1023 ( .A1(G227), .A2(n1094), .ZN(n1166) );
XOR2_X1 U1024 ( .A(n1274), .B(n1173), .Z(n1302) );
XOR2_X1 U1025 ( .A(n1287), .B(n1305), .Z(n1173) );
XOR2_X1 U1026 ( .A(KEYINPUT2), .B(n1084), .Z(n1305) );
XNOR2_X1 U1027 ( .A(n1306), .B(n1307), .ZN(n1084) );
NOR2_X1 U1028 ( .A1(n1297), .A2(n1308), .ZN(n1307) );
NOR2_X1 U1029 ( .A1(G146), .A2(n1309), .ZN(n1308) );
NOR2_X1 U1030 ( .A1(n1298), .A2(G143), .ZN(n1297) );
NAND2_X1 U1031 ( .A1(KEYINPUT50), .A2(n1227), .ZN(n1306) );
INV_X1 U1032 ( .A(G128), .ZN(n1227) );
XNOR2_X1 U1033 ( .A(G104), .B(n1310), .ZN(n1287) );
INV_X1 U1034 ( .A(G107), .ZN(n1310) );
XOR2_X1 U1035 ( .A(G101), .B(n1150), .Z(n1274) );
XNOR2_X1 U1036 ( .A(G134), .B(n1083), .ZN(n1150) );
XOR2_X1 U1037 ( .A(G131), .B(G137), .Z(n1083) );
NOR2_X1 U1038 ( .A1(n1221), .A2(n1219), .ZN(n1023) );
INV_X1 U1039 ( .A(n1248), .ZN(n1219) );
XOR2_X1 U1040 ( .A(n1067), .B(n1311), .Z(n1248) );
NOR2_X1 U1041 ( .A1(KEYINPUT34), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1042 ( .A(KEYINPUT16), .B(n1125), .ZN(n1312) );
INV_X1 U1043 ( .A(G478), .ZN(n1125) );
NOR2_X1 U1044 ( .A1(n1123), .A2(G902), .ZN(n1067) );
XNOR2_X1 U1045 ( .A(n1313), .B(n1314), .ZN(n1123) );
XOR2_X1 U1046 ( .A(n1315), .B(n1316), .Z(n1314) );
AND2_X1 U1047 ( .A1(n1269), .A2(G217), .ZN(n1316) );
AND2_X1 U1048 ( .A1(G234), .A2(n1094), .ZN(n1269) );
NOR2_X1 U1049 ( .A1(KEYINPUT3), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1050 ( .A(n1318), .B(n1319), .Z(n1317) );
NOR2_X1 U1051 ( .A1(KEYINPUT48), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1052 ( .A(KEYINPUT15), .B(n1309), .ZN(n1320) );
INV_X1 U1053 ( .A(G143), .ZN(n1309) );
XNOR2_X1 U1054 ( .A(G128), .B(G134), .ZN(n1318) );
XNOR2_X1 U1055 ( .A(G107), .B(n1321), .ZN(n1313) );
XNOR2_X1 U1056 ( .A(n1235), .B(G116), .ZN(n1321) );
XNOR2_X1 U1057 ( .A(n1069), .B(n1322), .ZN(n1221) );
XNOR2_X1 U1058 ( .A(KEYINPUT62), .B(n1070), .ZN(n1322) );
INV_X1 U1059 ( .A(G475), .ZN(n1070) );
NAND2_X1 U1060 ( .A1(n1131), .A2(n1177), .ZN(n1069) );
INV_X1 U1061 ( .A(G902), .ZN(n1177) );
XNOR2_X1 U1062 ( .A(n1323), .B(n1324), .ZN(n1131) );
XOR2_X1 U1063 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1064 ( .A(n1327), .B(n1328), .Z(n1326) );
AND3_X1 U1065 ( .A1(n1278), .A2(n1094), .A3(G214), .ZN(n1328) );
INV_X1 U1066 ( .A(G953), .ZN(n1094) );
XOR2_X1 U1067 ( .A(n1281), .B(KEYINPUT46), .Z(n1278) );
INV_X1 U1068 ( .A(G237), .ZN(n1281) );
NAND2_X1 U1069 ( .A1(KEYINPUT17), .A2(n1235), .ZN(n1327) );
INV_X1 U1070 ( .A(G122), .ZN(n1235) );
XNOR2_X1 U1071 ( .A(G131), .B(G143), .ZN(n1325) );
XOR2_X1 U1072 ( .A(n1329), .B(n1330), .Z(n1323) );
XNOR2_X1 U1073 ( .A(n1262), .B(n1277), .ZN(n1330) );
XNOR2_X1 U1074 ( .A(G113), .B(KEYINPUT14), .ZN(n1277) );
XNOR2_X1 U1075 ( .A(G140), .B(n1298), .ZN(n1262) );
INV_X1 U1076 ( .A(G146), .ZN(n1298) );
XOR2_X1 U1077 ( .A(n1331), .B(n1332), .Z(n1329) );
NOR2_X1 U1078 ( .A1(G125), .A2(KEYINPUT39), .ZN(n1332) );
NAND2_X1 U1079 ( .A1(KEYINPUT22), .A2(n1333), .ZN(n1331) );
INV_X1 U1080 ( .A(G104), .ZN(n1333) );
endmodule


