//Key = 0110101000101010000001111010000111000000101000111011100110100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U737 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
NAND3_X1 U741 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND3_X1 U743 ( .A1(n1042), .A2(n1043), .A3(KEYINPUT29), .ZN(n1040) );
NAND3_X1 U744 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1037) );
NAND2_X1 U745 ( .A1(n1042), .A2(n1047), .ZN(n1045) );
NAND2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
OR2_X1 U747 ( .A1(n1050), .A2(KEYINPUT29), .ZN(n1049) );
NAND2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1044) );
NAND2_X1 U749 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U753 ( .A(n1061), .ZN(n1057) );
NAND2_X1 U754 ( .A1(n1062), .A2(n1063), .ZN(n1053) );
NAND2_X1 U755 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U756 ( .A1(KEYINPUT22), .A2(n1066), .ZN(n1065) );
NAND2_X1 U757 ( .A1(n1067), .A2(n1068), .ZN(n1035) );
INV_X1 U758 ( .A(KEYINPUT22), .ZN(n1068) );
NAND4_X1 U759 ( .A1(n1039), .A2(n1069), .A3(n1070), .A4(n1046), .ZN(n1067) );
NAND4_X1 U760 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1031) );
NAND3_X1 U761 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1072) );
NAND2_X1 U762 ( .A1(n1078), .A2(n1079), .ZN(n1071) );
XOR2_X1 U763 ( .A(KEYINPUT62), .B(n1077), .Z(n1079) );
AND3_X1 U764 ( .A1(n1042), .A2(n1051), .A3(n1039), .ZN(n1077) );
INV_X1 U765 ( .A(n1080), .ZN(n1039) );
NOR3_X1 U766 ( .A1(n1081), .A2(G953), .A3(G952), .ZN(n1029) );
INV_X1 U767 ( .A(n1073), .ZN(n1081) );
NAND4_X1 U768 ( .A1(n1082), .A2(n1075), .A3(n1083), .A4(n1084), .ZN(n1073) );
NOR4_X1 U769 ( .A1(n1085), .A2(n1086), .A3(n1059), .A4(n1076), .ZN(n1084) );
NAND2_X1 U770 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
INV_X1 U771 ( .A(n1089), .ZN(n1085) );
NOR3_X1 U772 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1083) );
XNOR2_X1 U773 ( .A(G469), .B(n1093), .ZN(n1092) );
NOR2_X1 U774 ( .A1(n1094), .A2(KEYINPUT49), .ZN(n1093) );
NOR2_X1 U775 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
XNOR2_X1 U776 ( .A(n1097), .B(KEYINPUT51), .ZN(n1090) );
XNOR2_X1 U777 ( .A(n1098), .B(KEYINPUT37), .ZN(n1082) );
XOR2_X1 U778 ( .A(n1099), .B(n1100), .Z(G72) );
XOR2_X1 U779 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U780 ( .A1(G953), .A2(n1103), .ZN(n1102) );
NAND2_X1 U781 ( .A1(n1104), .A2(G900), .ZN(n1103) );
XNOR2_X1 U782 ( .A(G227), .B(KEYINPUT55), .ZN(n1104) );
NAND2_X1 U783 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
NAND2_X1 U784 ( .A1(G953), .A2(n1107), .ZN(n1106) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(n1105) );
XNOR2_X1 U786 ( .A(n1110), .B(n1111), .ZN(n1109) );
XOR2_X1 U787 ( .A(n1112), .B(n1113), .Z(n1108) );
XNOR2_X1 U788 ( .A(G140), .B(n1114), .ZN(n1112) );
NOR2_X1 U789 ( .A1(KEYINPUT53), .A2(n1115), .ZN(n1114) );
NOR2_X1 U790 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U791 ( .A(KEYINPUT5), .B(n1118), .Z(n1117) );
AND2_X1 U792 ( .A1(n1119), .A2(G137), .ZN(n1118) );
NOR2_X1 U793 ( .A1(G137), .A2(n1119), .ZN(n1116) );
AND2_X1 U794 ( .A1(n1034), .A2(n1074), .ZN(n1099) );
NAND2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(G69) );
NAND2_X1 U796 ( .A1(G953), .A2(n1122), .ZN(n1121) );
NAND2_X1 U797 ( .A1(G898), .A2(n1123), .ZN(n1122) );
XOR2_X1 U798 ( .A(G224), .B(n1124), .Z(n1123) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1074), .ZN(n1120) );
XOR2_X1 U800 ( .A(n1033), .B(n1124), .Z(n1125) );
XNOR2_X1 U801 ( .A(n1126), .B(n1127), .ZN(n1124) );
XOR2_X1 U802 ( .A(KEYINPUT63), .B(KEYINPUT14), .Z(n1127) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1126) );
NOR2_X1 U804 ( .A1(KEYINPUT18), .A2(n1130), .ZN(n1129) );
NOR2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR3_X1 U807 ( .A1(n1135), .A2(KEYINPUT17), .A3(n1136), .ZN(n1133) );
INV_X1 U808 ( .A(G217), .ZN(n1136) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1137), .ZN(G63) );
XOR2_X1 U810 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U811 ( .A1(n1140), .A2(n1135), .ZN(n1139) );
NAND2_X1 U812 ( .A1(KEYINPUT42), .A2(n1141), .ZN(n1138) );
NOR2_X1 U813 ( .A1(n1131), .A2(n1142), .ZN(G60) );
XOR2_X1 U814 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U815 ( .A1(n1145), .A2(G475), .ZN(n1144) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(G6) );
XOR2_X1 U817 ( .A(KEYINPUT23), .B(G104), .Z(n1147) );
NOR2_X1 U818 ( .A1(n1131), .A2(n1148), .ZN(G57) );
XOR2_X1 U819 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U821 ( .A1(n1145), .A2(G472), .ZN(n1151) );
XOR2_X1 U822 ( .A(n1153), .B(n1154), .Z(n1149) );
NAND2_X1 U823 ( .A1(KEYINPUT50), .A2(n1155), .ZN(n1154) );
NOR2_X1 U824 ( .A1(n1131), .A2(n1156), .ZN(G54) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U826 ( .A(n1159), .B(n1160), .ZN(n1158) );
XNOR2_X1 U827 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U828 ( .A(n1163), .B(n1164), .Z(n1157) );
XNOR2_X1 U829 ( .A(KEYINPUT46), .B(n1165), .ZN(n1164) );
NOR2_X1 U830 ( .A1(KEYINPUT34), .A2(n1166), .ZN(n1165) );
NAND2_X1 U831 ( .A1(n1145), .A2(G469), .ZN(n1163) );
NOR2_X1 U832 ( .A1(n1131), .A2(n1167), .ZN(G51) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U834 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U835 ( .A1(n1145), .A2(n1172), .ZN(n1170) );
INV_X1 U836 ( .A(n1135), .ZN(n1145) );
NAND2_X1 U837 ( .A1(G902), .A2(n1173), .ZN(n1135) );
OR2_X1 U838 ( .A1(n1034), .A2(n1033), .ZN(n1173) );
NAND4_X1 U839 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1033) );
NOR4_X1 U840 ( .A1(n1178), .A2(n1179), .A3(n1146), .A4(n1180), .ZN(n1177) );
INV_X1 U841 ( .A(n1028), .ZN(n1180) );
NAND3_X1 U842 ( .A1(n1055), .A2(n1043), .A3(n1181), .ZN(n1028) );
AND3_X1 U843 ( .A1(n1181), .A2(n1055), .A3(n1182), .ZN(n1146) );
NAND2_X1 U844 ( .A1(n1078), .A2(n1183), .ZN(n1176) );
NAND2_X1 U845 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U846 ( .A(n1186), .B(KEYINPUT44), .Z(n1184) );
NAND2_X1 U847 ( .A1(n1187), .A2(n1188), .ZN(n1034) );
AND4_X1 U848 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NOR4_X1 U849 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1187) );
NOR3_X1 U850 ( .A1(n1197), .A2(n1198), .A3(n1050), .ZN(n1196) );
NOR3_X1 U851 ( .A1(n1199), .A2(n1041), .A3(n1200), .ZN(n1195) );
XNOR2_X1 U852 ( .A(KEYINPUT20), .B(n1201), .ZN(n1200) );
NAND3_X1 U853 ( .A1(n1182), .A2(n1061), .A3(n1066), .ZN(n1199) );
XNOR2_X1 U854 ( .A(n1202), .B(n1203), .ZN(n1168) );
NOR2_X1 U855 ( .A1(KEYINPUT36), .A2(n1204), .ZN(n1203) );
NOR2_X1 U856 ( .A1(n1074), .A2(G952), .ZN(n1131) );
XOR2_X1 U857 ( .A(n1192), .B(n1205), .Z(G48) );
XOR2_X1 U858 ( .A(KEYINPUT48), .B(G146), .Z(n1205) );
NAND2_X1 U859 ( .A1(n1206), .A2(n1207), .ZN(n1192) );
NAND3_X1 U860 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(G45) );
NAND2_X1 U861 ( .A1(G143), .A2(n1211), .ZN(n1210) );
NAND2_X1 U862 ( .A1(KEYINPUT0), .A2(n1212), .ZN(n1209) );
NAND2_X1 U863 ( .A1(n1194), .A2(n1213), .ZN(n1212) );
XNOR2_X1 U864 ( .A(KEYINPUT52), .B(n1214), .ZN(n1213) );
NAND2_X1 U865 ( .A1(n1215), .A2(n1216), .ZN(n1208) );
INV_X1 U866 ( .A(KEYINPUT0), .ZN(n1216) );
NAND2_X1 U867 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NAND3_X1 U868 ( .A1(KEYINPUT52), .A2(n1194), .A3(n1214), .ZN(n1218) );
INV_X1 U869 ( .A(n1211), .ZN(n1194) );
NAND3_X1 U870 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1211) );
AND3_X1 U871 ( .A1(n1078), .A2(n1222), .A3(n1097), .ZN(n1221) );
OR2_X1 U872 ( .A1(n1214), .A2(KEYINPUT52), .ZN(n1217) );
XNOR2_X1 U873 ( .A(n1223), .B(n1224), .ZN(G42) );
NOR4_X1 U874 ( .A1(n1225), .A2(n1048), .A3(n1226), .A4(n1227), .ZN(n1224) );
XNOR2_X1 U875 ( .A(n1046), .B(KEYINPUT9), .ZN(n1225) );
XNOR2_X1 U876 ( .A(G137), .B(n1191), .ZN(G39) );
NAND3_X1 U877 ( .A1(n1046), .A2(n1051), .A3(n1206), .ZN(n1191) );
INV_X1 U878 ( .A(n1197), .ZN(n1206) );
XNOR2_X1 U879 ( .A(n1119), .B(n1193), .ZN(G36) );
NOR4_X1 U880 ( .A1(n1064), .A2(n1227), .A3(n1041), .A4(n1050), .ZN(n1193) );
INV_X1 U881 ( .A(n1219), .ZN(n1064) );
XNOR2_X1 U882 ( .A(G131), .B(n1190), .ZN(G33) );
NAND4_X1 U883 ( .A1(n1219), .A2(n1220), .A3(n1046), .A4(n1182), .ZN(n1190) );
INV_X1 U884 ( .A(n1041), .ZN(n1046) );
NAND2_X1 U885 ( .A1(n1075), .A2(n1228), .ZN(n1041) );
INV_X1 U886 ( .A(n1229), .ZN(n1228) );
XOR2_X1 U887 ( .A(G128), .B(n1230), .Z(G30) );
NOR3_X1 U888 ( .A1(n1231), .A2(n1050), .A3(n1197), .ZN(n1230) );
NAND3_X1 U889 ( .A1(n1098), .A2(n1232), .A3(n1220), .ZN(n1197) );
INV_X1 U890 ( .A(n1227), .ZN(n1220) );
NAND2_X1 U891 ( .A1(n1061), .A2(n1201), .ZN(n1227) );
XNOR2_X1 U892 ( .A(KEYINPUT26), .B(n1198), .ZN(n1231) );
XNOR2_X1 U893 ( .A(G101), .B(n1174), .ZN(G3) );
NAND3_X1 U894 ( .A1(n1181), .A2(n1051), .A3(n1219), .ZN(n1174) );
XNOR2_X1 U895 ( .A(G125), .B(n1189), .ZN(G27) );
NAND4_X1 U896 ( .A1(n1062), .A2(n1066), .A3(n1207), .A4(n1201), .ZN(n1189) );
NAND2_X1 U897 ( .A1(n1080), .A2(n1233), .ZN(n1201) );
NAND4_X1 U898 ( .A1(G902), .A2(G953), .A3(n1234), .A4(n1107), .ZN(n1233) );
INV_X1 U899 ( .A(G900), .ZN(n1107) );
XNOR2_X1 U900 ( .A(n1235), .B(n1236), .ZN(G24) );
NOR2_X1 U901 ( .A1(n1237), .A2(n1185), .ZN(n1236) );
NAND4_X1 U902 ( .A1(n1042), .A2(n1097), .A3(n1222), .A4(n1238), .ZN(n1185) );
AND2_X1 U903 ( .A1(n1062), .A2(n1055), .ZN(n1042) );
NOR2_X1 U904 ( .A1(n1232), .A2(n1098), .ZN(n1055) );
XNOR2_X1 U905 ( .A(n1078), .B(KEYINPUT35), .ZN(n1237) );
XNOR2_X1 U906 ( .A(G119), .B(n1175), .ZN(G21) );
NAND4_X1 U907 ( .A1(n1069), .A2(n1078), .A3(n1098), .A4(n1238), .ZN(n1175) );
AND3_X1 U908 ( .A1(n1051), .A2(n1232), .A3(n1062), .ZN(n1069) );
XNOR2_X1 U909 ( .A(G116), .B(n1239), .ZN(G18) );
NOR2_X1 U910 ( .A1(n1240), .A2(KEYINPUT41), .ZN(n1239) );
NOR2_X1 U911 ( .A1(n1198), .A2(n1186), .ZN(n1240) );
NAND4_X1 U912 ( .A1(n1219), .A2(n1062), .A3(n1043), .A4(n1238), .ZN(n1186) );
INV_X1 U913 ( .A(n1050), .ZN(n1043) );
NAND2_X1 U914 ( .A1(n1241), .A2(n1242), .ZN(n1050) );
XNOR2_X1 U915 ( .A(KEYINPUT1), .B(n1222), .ZN(n1242) );
XNOR2_X1 U916 ( .A(KEYINPUT13), .B(n1097), .ZN(n1241) );
XNOR2_X1 U917 ( .A(G113), .B(n1243), .ZN(G15) );
NOR2_X1 U918 ( .A1(n1179), .A2(KEYINPUT8), .ZN(n1243) );
AND4_X1 U919 ( .A1(n1219), .A2(n1062), .A3(n1207), .A4(n1238), .ZN(n1179) );
NOR2_X1 U920 ( .A1(n1048), .A2(n1198), .ZN(n1207) );
INV_X1 U921 ( .A(n1078), .ZN(n1198) );
INV_X1 U922 ( .A(n1182), .ZN(n1048) );
NOR2_X1 U923 ( .A1(n1244), .A2(n1059), .ZN(n1062) );
NOR2_X1 U924 ( .A1(n1232), .A2(n1070), .ZN(n1219) );
XOR2_X1 U925 ( .A(n1178), .B(n1245), .Z(G12) );
NOR2_X1 U926 ( .A1(KEYINPUT25), .A2(n1246), .ZN(n1245) );
AND3_X1 U927 ( .A1(n1181), .A2(n1051), .A3(n1066), .ZN(n1178) );
INV_X1 U928 ( .A(n1226), .ZN(n1066) );
NAND2_X1 U929 ( .A1(n1070), .A2(n1232), .ZN(n1226) );
NAND3_X1 U930 ( .A1(n1247), .A2(n1248), .A3(n1089), .ZN(n1232) );
NAND2_X1 U931 ( .A1(n1095), .A2(n1096), .ZN(n1089) );
NAND2_X1 U932 ( .A1(n1096), .A2(n1249), .ZN(n1248) );
OR3_X1 U933 ( .A1(n1096), .A2(n1095), .A3(n1249), .ZN(n1247) );
INV_X1 U934 ( .A(KEYINPUT47), .ZN(n1249) );
NOR2_X1 U935 ( .A1(n1134), .A2(G902), .ZN(n1095) );
XNOR2_X1 U936 ( .A(n1250), .B(n1251), .ZN(n1134) );
XOR2_X1 U937 ( .A(G119), .B(n1252), .Z(n1251) );
XOR2_X1 U938 ( .A(KEYINPUT30), .B(G137), .Z(n1252) );
XOR2_X1 U939 ( .A(n1253), .B(n1162), .Z(n1250) );
XOR2_X1 U940 ( .A(n1110), .B(n1254), .Z(n1253) );
AND4_X1 U941 ( .A1(n1255), .A2(n1256), .A3(G234), .A4(G221), .ZN(n1254) );
INV_X1 U942 ( .A(KEYINPUT16), .ZN(n1255) );
NAND2_X1 U943 ( .A1(n1257), .A2(G217), .ZN(n1096) );
XOR2_X1 U944 ( .A(n1258), .B(KEYINPUT57), .Z(n1257) );
INV_X1 U945 ( .A(n1098), .ZN(n1070) );
XNOR2_X1 U946 ( .A(n1259), .B(G472), .ZN(n1098) );
NAND2_X1 U947 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U948 ( .A(n1262), .B(n1263), .Z(n1260) );
XNOR2_X1 U949 ( .A(G101), .B(n1153), .ZN(n1263) );
NAND3_X1 U950 ( .A1(n1256), .A2(n1264), .A3(G210), .ZN(n1153) );
NOR2_X1 U951 ( .A1(KEYINPUT39), .A2(n1152), .ZN(n1262) );
XOR2_X1 U952 ( .A(n1265), .B(n1266), .Z(n1152) );
XNOR2_X1 U953 ( .A(n1267), .B(n1268), .ZN(n1266) );
XOR2_X1 U954 ( .A(n1269), .B(G119), .Z(n1268) );
XOR2_X1 U955 ( .A(n1270), .B(n1271), .Z(n1265) );
NAND2_X1 U956 ( .A1(n1272), .A2(n1273), .ZN(n1051) );
OR3_X1 U957 ( .A1(n1222), .A2(n1097), .A3(KEYINPUT13), .ZN(n1273) );
NAND2_X1 U958 ( .A1(KEYINPUT13), .A2(n1182), .ZN(n1272) );
NOR2_X1 U959 ( .A1(n1222), .A2(n1274), .ZN(n1182) );
INV_X1 U960 ( .A(n1097), .ZN(n1274) );
XNOR2_X1 U961 ( .A(n1275), .B(G475), .ZN(n1097) );
NAND2_X1 U962 ( .A1(n1261), .A2(n1143), .ZN(n1275) );
NAND2_X1 U963 ( .A1(n1276), .A2(n1277), .ZN(n1143) );
NAND2_X1 U964 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U965 ( .A(n1280), .B(KEYINPUT54), .Z(n1276) );
OR2_X1 U966 ( .A1(n1279), .A2(n1278), .ZN(n1280) );
XOR2_X1 U967 ( .A(n1281), .B(n1282), .Z(n1278) );
NOR2_X1 U968 ( .A1(KEYINPUT43), .A2(G113), .ZN(n1282) );
XNOR2_X1 U969 ( .A(G104), .B(G122), .ZN(n1281) );
XNOR2_X1 U970 ( .A(n1283), .B(n1284), .ZN(n1279) );
XNOR2_X1 U971 ( .A(n1223), .B(G125), .ZN(n1284) );
XOR2_X1 U972 ( .A(n1285), .B(n1286), .Z(n1283) );
NAND2_X1 U973 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
NAND2_X1 U974 ( .A1(n1289), .A2(n1113), .ZN(n1288) );
XOR2_X1 U975 ( .A(n1290), .B(KEYINPUT59), .Z(n1287) );
OR2_X1 U976 ( .A1(n1289), .A2(n1113), .ZN(n1290) );
XOR2_X1 U977 ( .A(n1291), .B(n1214), .Z(n1289) );
NAND3_X1 U978 ( .A1(G214), .A2(n1256), .A3(n1292), .ZN(n1291) );
XNOR2_X1 U979 ( .A(G237), .B(KEYINPUT15), .ZN(n1292) );
NAND2_X1 U980 ( .A1(n1293), .A2(n1087), .ZN(n1222) );
NAND3_X1 U981 ( .A1(n1140), .A2(n1261), .A3(n1141), .ZN(n1087) );
INV_X1 U982 ( .A(G478), .ZN(n1140) );
XOR2_X1 U983 ( .A(n1088), .B(KEYINPUT28), .Z(n1293) );
NAND2_X1 U984 ( .A1(G478), .A2(n1294), .ZN(n1088) );
NAND2_X1 U985 ( .A1(n1141), .A2(n1261), .ZN(n1294) );
XNOR2_X1 U986 ( .A(n1295), .B(n1296), .ZN(n1141) );
XNOR2_X1 U987 ( .A(n1297), .B(n1298), .ZN(n1296) );
XNOR2_X1 U988 ( .A(n1119), .B(G128), .ZN(n1298) );
INV_X1 U989 ( .A(G134), .ZN(n1119) );
XOR2_X1 U990 ( .A(n1299), .B(n1300), .Z(n1295) );
XOR2_X1 U991 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U992 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U993 ( .A1(G116), .A2(n1235), .ZN(n1304) );
XOR2_X1 U994 ( .A(n1305), .B(KEYINPUT3), .Z(n1303) );
OR2_X1 U995 ( .A1(n1235), .A2(G116), .ZN(n1305) );
NAND3_X1 U996 ( .A1(G217), .A2(n1256), .A3(n1306), .ZN(n1301) );
XNOR2_X1 U997 ( .A(G234), .B(KEYINPUT2), .ZN(n1306) );
NAND2_X1 U998 ( .A1(KEYINPUT32), .A2(n1214), .ZN(n1299) );
AND3_X1 U999 ( .A1(n1078), .A2(n1238), .A3(n1061), .ZN(n1181) );
NOR2_X1 U1000 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
AND2_X1 U1001 ( .A1(G221), .A2(n1258), .ZN(n1059) );
NAND2_X1 U1002 ( .A1(n1307), .A2(n1261), .ZN(n1258) );
INV_X1 U1003 ( .A(n1244), .ZN(n1060) );
XNOR2_X1 U1004 ( .A(n1308), .B(n1094), .ZN(n1244) );
AND2_X1 U1005 ( .A1(n1309), .A2(n1261), .ZN(n1094) );
XOR2_X1 U1006 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1007 ( .A(n1312), .B(n1166), .ZN(n1311) );
AND2_X1 U1008 ( .A1(n1313), .A2(n1314), .ZN(n1166) );
NAND2_X1 U1009 ( .A1(n1315), .A2(G107), .ZN(n1314) );
NAND2_X1 U1010 ( .A1(n1316), .A2(n1297), .ZN(n1313) );
INV_X1 U1011 ( .A(G107), .ZN(n1297) );
XNOR2_X1 U1012 ( .A(n1315), .B(KEYINPUT45), .ZN(n1316) );
INV_X1 U1013 ( .A(n1159), .ZN(n1312) );
XNOR2_X1 U1014 ( .A(n1317), .B(n1271), .ZN(n1159) );
XNOR2_X1 U1015 ( .A(n1318), .B(n1113), .ZN(n1271) );
XOR2_X1 U1016 ( .A(G131), .B(KEYINPUT21), .Z(n1113) );
XNOR2_X1 U1017 ( .A(G134), .B(G137), .ZN(n1318) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1256), .ZN(n1317) );
XOR2_X1 U1019 ( .A(n1319), .B(n1320), .Z(n1310) );
XNOR2_X1 U1020 ( .A(KEYINPUT38), .B(n1321), .ZN(n1320) );
NOR2_X1 U1021 ( .A1(KEYINPUT11), .A2(n1161), .ZN(n1321) );
XOR2_X1 U1022 ( .A(n1270), .B(n1322), .Z(n1161) );
INV_X1 U1023 ( .A(n1111), .ZN(n1322) );
XOR2_X1 U1024 ( .A(G143), .B(KEYINPUT24), .Z(n1111) );
NAND2_X1 U1025 ( .A1(KEYINPUT12), .A2(n1162), .ZN(n1319) );
XNOR2_X1 U1026 ( .A(n1223), .B(n1323), .ZN(n1162) );
INV_X1 U1027 ( .A(G140), .ZN(n1223) );
NAND2_X1 U1028 ( .A1(KEYINPUT58), .A2(G469), .ZN(n1308) );
NAND2_X1 U1029 ( .A1(n1080), .A2(n1324), .ZN(n1238) );
NAND4_X1 U1030 ( .A1(G902), .A2(G953), .A3(n1234), .A4(n1325), .ZN(n1324) );
INV_X1 U1031 ( .A(G898), .ZN(n1325) );
NAND3_X1 U1032 ( .A1(n1234), .A2(n1074), .A3(G952), .ZN(n1080) );
INV_X1 U1033 ( .A(G953), .ZN(n1074) );
NAND2_X1 U1034 ( .A1(G237), .A2(n1307), .ZN(n1234) );
XNOR2_X1 U1035 ( .A(G234), .B(KEYINPUT31), .ZN(n1307) );
NOR2_X1 U1036 ( .A1(n1229), .A2(n1075), .ZN(n1078) );
XOR2_X1 U1037 ( .A(n1326), .B(n1172), .Z(n1075) );
AND2_X1 U1038 ( .A1(G210), .A2(n1327), .ZN(n1172) );
NAND2_X1 U1039 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
XOR2_X1 U1040 ( .A(n1171), .B(n1330), .Z(n1329) );
XNOR2_X1 U1041 ( .A(KEYINPUT40), .B(n1331), .ZN(n1330) );
NOR2_X1 U1042 ( .A1(KEYINPUT60), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1043 ( .A(n1202), .B(n1204), .ZN(n1332) );
XOR2_X1 U1044 ( .A(n1110), .B(n1269), .Z(n1204) );
NAND2_X1 U1045 ( .A1(KEYINPUT56), .A2(n1214), .ZN(n1269) );
INV_X1 U1046 ( .A(G143), .ZN(n1214) );
XOR2_X1 U1047 ( .A(n1270), .B(G125), .Z(n1110) );
XNOR2_X1 U1048 ( .A(G128), .B(n1286), .ZN(n1270) );
XOR2_X1 U1049 ( .A(G146), .B(KEYINPUT27), .Z(n1286) );
NAND2_X1 U1050 ( .A1(G224), .A2(n1256), .ZN(n1202) );
XOR2_X1 U1051 ( .A(G953), .B(KEYINPUT6), .Z(n1256) );
XOR2_X1 U1052 ( .A(n1333), .B(n1334), .Z(n1171) );
XOR2_X1 U1053 ( .A(KEYINPUT7), .B(KEYINPUT10), .Z(n1334) );
XNOR2_X1 U1054 ( .A(n1128), .B(n1130), .ZN(n1333) );
XOR2_X1 U1055 ( .A(n1235), .B(n1323), .Z(n1130) );
XNOR2_X1 U1056 ( .A(n1246), .B(KEYINPUT4), .ZN(n1323) );
INV_X1 U1057 ( .A(G110), .ZN(n1246) );
INV_X1 U1058 ( .A(G122), .ZN(n1235) );
XOR2_X1 U1059 ( .A(n1335), .B(n1336), .Z(n1128) );
XOR2_X1 U1060 ( .A(n1267), .B(n1315), .Z(n1336) );
XNOR2_X1 U1061 ( .A(G104), .B(n1155), .ZN(n1315) );
INV_X1 U1062 ( .A(G101), .ZN(n1155) );
XOR2_X1 U1063 ( .A(G113), .B(G116), .Z(n1267) );
XNOR2_X1 U1064 ( .A(G107), .B(n1337), .ZN(n1335) );
NOR2_X1 U1065 ( .A1(G119), .A2(KEYINPUT61), .ZN(n1337) );
XNOR2_X1 U1066 ( .A(KEYINPUT33), .B(n1261), .ZN(n1328) );
XOR2_X1 U1067 ( .A(n1076), .B(KEYINPUT19), .Z(n1229) );
AND2_X1 U1068 ( .A1(G214), .A2(n1327), .ZN(n1076) );
NAND2_X1 U1069 ( .A1(n1261), .A2(n1264), .ZN(n1327) );
INV_X1 U1070 ( .A(G237), .ZN(n1264) );
INV_X1 U1071 ( .A(G902), .ZN(n1261) );
endmodule


