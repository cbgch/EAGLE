//Key = 0101000101110101111010010110110010010111101101100110010100001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277;

XOR2_X1 U711 ( .A(G107), .B(n973), .Z(G9) );
NAND3_X1 U712 ( .A1(n974), .A2(n975), .A3(n976), .ZN(G75) );
NAND2_X1 U713 ( .A1(G952), .A2(n977), .ZN(n976) );
NAND2_X1 U714 ( .A1(n978), .A2(n979), .ZN(n977) );
NAND2_X1 U715 ( .A1(n980), .A2(n981), .ZN(n979) );
NAND2_X1 U716 ( .A1(n982), .A2(n983), .ZN(n980) );
NAND3_X1 U717 ( .A1(n984), .A2(n985), .A3(n986), .ZN(n983) );
NAND2_X1 U718 ( .A1(n987), .A2(n988), .ZN(n985) );
NAND2_X1 U719 ( .A1(n989), .A2(n990), .ZN(n988) );
OR2_X1 U720 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U721 ( .A1(n993), .A2(n994), .ZN(n987) );
NAND3_X1 U722 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
OR2_X1 U723 ( .A1(n998), .A2(KEYINPUT7), .ZN(n996) );
NAND3_X1 U724 ( .A1(n999), .A2(n1000), .A3(KEYINPUT7), .ZN(n995) );
NAND3_X1 U725 ( .A1(n989), .A2(n1001), .A3(n993), .ZN(n982) );
NAND3_X1 U726 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1001) );
NAND2_X1 U727 ( .A1(n986), .A2(n1005), .ZN(n1004) );
NAND2_X1 U728 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U729 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
XNOR2_X1 U730 ( .A(n1010), .B(KEYINPUT24), .ZN(n1006) );
NAND3_X1 U731 ( .A1(n1011), .A2(n984), .A3(n1012), .ZN(n1003) );
NAND2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(n1002) );
XNOR2_X1 U733 ( .A(KEYINPUT33), .B(n1015), .ZN(n1014) );
NAND4_X1 U734 ( .A1(n1016), .A2(n989), .A3(n1017), .A4(n1018), .ZN(n974) );
NOR3_X1 U735 ( .A1(n1015), .A2(n1012), .A3(n1019), .ZN(n1018) );
XNOR2_X1 U736 ( .A(n1020), .B(n1021), .ZN(n1019) );
NAND2_X1 U737 ( .A1(KEYINPUT17), .A2(n1022), .ZN(n1020) );
INV_X1 U738 ( .A(n984), .ZN(n1015) );
XNOR2_X1 U739 ( .A(n1023), .B(n1024), .ZN(n1017) );
NAND2_X1 U740 ( .A1(KEYINPUT37), .A2(n1025), .ZN(n1023) );
XNOR2_X1 U741 ( .A(n1026), .B(G475), .ZN(n1016) );
XOR2_X1 U742 ( .A(n1027), .B(n1028), .Z(G72) );
NOR2_X1 U743 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
XOR2_X1 U744 ( .A(KEYINPUT57), .B(n1031), .Z(n1030) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
AND2_X1 U746 ( .A1(n1033), .A2(n1032), .ZN(n1029) );
AND2_X1 U747 ( .A1(n1034), .A2(n975), .ZN(n1032) );
NAND2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XOR2_X1 U749 ( .A(KEYINPUT30), .B(n1037), .Z(n1036) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1033) );
XOR2_X1 U751 ( .A(KEYINPUT63), .B(n1040), .Z(n1039) );
NOR2_X1 U752 ( .A1(G900), .A2(n975), .ZN(n1040) );
XOR2_X1 U753 ( .A(n1041), .B(n1042), .Z(n1038) );
XOR2_X1 U754 ( .A(n1043), .B(n1044), .Z(n1042) );
XNOR2_X1 U755 ( .A(G131), .B(n1045), .ZN(n1044) );
XNOR2_X1 U756 ( .A(KEYINPUT18), .B(n1046), .ZN(n1043) );
XOR2_X1 U757 ( .A(n1047), .B(n1048), .Z(n1041) );
NOR2_X1 U758 ( .A1(G140), .A2(KEYINPUT5), .ZN(n1048) );
XNOR2_X1 U759 ( .A(n1049), .B(n1050), .ZN(n1047) );
NOR2_X1 U760 ( .A1(KEYINPUT6), .A2(n1051), .ZN(n1050) );
NOR2_X1 U761 ( .A1(KEYINPUT34), .A2(n1052), .ZN(n1049) );
NOR2_X1 U762 ( .A1(KEYINPUT14), .A2(n1053), .ZN(n1027) );
NOR2_X1 U763 ( .A1(n1054), .A2(n975), .ZN(n1053) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1054) );
NAND2_X1 U765 ( .A1(n1055), .A2(n1056), .ZN(G69) );
NAND2_X1 U766 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U767 ( .A1(G953), .A2(n1059), .ZN(n1058) );
NAND3_X1 U768 ( .A1(G953), .A2(n1060), .A3(n1061), .ZN(n1055) );
XNOR2_X1 U769 ( .A(n1057), .B(KEYINPUT52), .ZN(n1061) );
XNOR2_X1 U770 ( .A(n1062), .B(n1063), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1064), .A2(G953), .ZN(n1063) );
NAND2_X1 U772 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U773 ( .A1(G953), .A2(n1067), .ZN(n1066) );
XOR2_X1 U774 ( .A(n1068), .B(n1069), .Z(n1065) );
XNOR2_X1 U775 ( .A(n1070), .B(KEYINPUT15), .ZN(n1069) );
NAND2_X1 U776 ( .A1(KEYINPUT29), .A2(n1071), .ZN(n1070) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1060) );
NOR2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XOR2_X1 U779 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U780 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U781 ( .A1(n1072), .A2(n1078), .ZN(G63) );
XNOR2_X1 U782 ( .A(n1079), .B(n1080), .ZN(n1078) );
NOR2_X1 U783 ( .A1(n1024), .A2(n1077), .ZN(n1080) );
NOR2_X1 U784 ( .A1(n1072), .A2(n1081), .ZN(G60) );
NOR3_X1 U785 ( .A1(n1026), .A2(n1082), .A3(n1083), .ZN(n1081) );
NOR3_X1 U786 ( .A1(n1084), .A2(n1085), .A3(n1077), .ZN(n1083) );
NOR2_X1 U787 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NOR2_X1 U788 ( .A1(n978), .A2(n1085), .ZN(n1086) );
INV_X1 U789 ( .A(n1088), .ZN(n978) );
NAND2_X1 U790 ( .A1(n1089), .A2(n1090), .ZN(G6) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U792 ( .A(n1093), .B(KEYINPUT19), .Z(n1089) );
OR2_X1 U793 ( .A1(n1092), .A2(n1091), .ZN(n1093) );
INV_X1 U794 ( .A(n1094), .ZN(n1091) );
XOR2_X1 U795 ( .A(G104), .B(KEYINPUT9), .Z(n1092) );
NOR2_X1 U796 ( .A1(n1072), .A2(n1095), .ZN(G57) );
XOR2_X1 U797 ( .A(n1096), .B(n1097), .Z(n1095) );
XNOR2_X1 U798 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR3_X1 U799 ( .A1(n1077), .A2(KEYINPUT54), .A3(n1100), .ZN(n1099) );
NAND2_X1 U800 ( .A1(KEYINPUT28), .A2(n1101), .ZN(n1098) );
NOR2_X1 U801 ( .A1(n1072), .A2(n1102), .ZN(G54) );
XOR2_X1 U802 ( .A(n1103), .B(n1104), .Z(n1102) );
XNOR2_X1 U803 ( .A(n1101), .B(n1105), .ZN(n1104) );
XNOR2_X1 U804 ( .A(n1106), .B(n1107), .ZN(n1105) );
NAND2_X1 U805 ( .A1(KEYINPUT23), .A2(n1108), .ZN(n1106) );
XOR2_X1 U806 ( .A(n1109), .B(n1110), .Z(n1103) );
XOR2_X1 U807 ( .A(G140), .B(n1111), .Z(n1110) );
NOR2_X1 U808 ( .A1(n1112), .A2(n1077), .ZN(n1109) );
NOR2_X1 U809 ( .A1(n1072), .A2(n1113), .ZN(G51) );
XOR2_X1 U810 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U811 ( .A(n1052), .B(n1116), .ZN(n1115) );
XOR2_X1 U812 ( .A(n1117), .B(n1118), .Z(n1114) );
XNOR2_X1 U813 ( .A(n1045), .B(n1119), .ZN(n1118) );
NOR2_X1 U814 ( .A1(n1021), .A2(n1077), .ZN(n1117) );
NAND2_X1 U815 ( .A1(G902), .A2(n1088), .ZN(n1077) );
NAND3_X1 U816 ( .A1(n1064), .A2(n1035), .A3(n1037), .ZN(n1088) );
AND4_X1 U817 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1037) );
AND3_X1 U818 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1035) );
NAND2_X1 U819 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U820 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U821 ( .A1(n1131), .A2(n993), .ZN(n1130) );
XNOR2_X1 U822 ( .A(n986), .B(KEYINPUT60), .ZN(n1131) );
NAND2_X1 U823 ( .A1(n991), .A2(n1013), .ZN(n1129) );
NAND2_X1 U824 ( .A1(n1132), .A2(n1133), .ZN(n1124) );
INV_X1 U825 ( .A(n1134), .ZN(n1133) );
XNOR2_X1 U826 ( .A(n1135), .B(KEYINPUT39), .ZN(n1132) );
AND4_X1 U827 ( .A1(n1136), .A2(n1094), .A3(n1137), .A4(n1138), .ZN(n1064) );
NOR4_X1 U828 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n973), .ZN(n1138) );
AND3_X1 U829 ( .A1(n984), .A2(n1142), .A3(n992), .ZN(n973) );
AND2_X1 U830 ( .A1(n1143), .A2(n1144), .ZN(n1137) );
NAND3_X1 U831 ( .A1(n984), .A2(n1142), .A3(n991), .ZN(n1094) );
NAND4_X1 U832 ( .A1(n1145), .A2(n1146), .A3(n989), .A4(n1147), .ZN(n1136) );
XNOR2_X1 U833 ( .A(n993), .B(KEYINPUT38), .ZN(n1145) );
NOR2_X1 U834 ( .A1(n975), .A2(G952), .ZN(n1072) );
XNOR2_X1 U835 ( .A(G146), .B(n1148), .ZN(G48) );
NAND3_X1 U836 ( .A1(n991), .A2(n1149), .A3(n1127), .ZN(n1148) );
XOR2_X1 U837 ( .A(KEYINPUT2), .B(n1013), .Z(n1149) );
XNOR2_X1 U838 ( .A(n1150), .B(n1151), .ZN(G45) );
NOR2_X1 U839 ( .A1(n997), .A2(n1134), .ZN(n1151) );
NAND4_X1 U840 ( .A1(n1152), .A2(n1010), .A3(n1153), .A4(n1013), .ZN(n1134) );
NOR2_X1 U841 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XNOR2_X1 U842 ( .A(G140), .B(n1125), .ZN(G42) );
NAND3_X1 U843 ( .A1(n1156), .A2(n1135), .A3(n986), .ZN(n1125) );
XOR2_X1 U844 ( .A(G137), .B(n1157), .Z(G39) );
AND3_X1 U845 ( .A1(n993), .A2(n1127), .A3(n986), .ZN(n1157) );
XNOR2_X1 U846 ( .A(G134), .B(n1121), .ZN(G36) );
NAND4_X1 U847 ( .A1(n1010), .A2(n986), .A3(n1158), .A4(n992), .ZN(n1121) );
NOR2_X1 U848 ( .A1(n1154), .A2(n997), .ZN(n1158) );
INV_X1 U849 ( .A(n1135), .ZN(n997) );
INV_X1 U850 ( .A(n1159), .ZN(n1154) );
XOR2_X1 U851 ( .A(n1160), .B(G131), .Z(G33) );
NAND2_X1 U852 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
OR2_X1 U853 ( .A1(n1120), .A2(KEYINPUT0), .ZN(n1162) );
OR2_X1 U854 ( .A1(n1163), .A2(n1164), .ZN(n1120) );
NAND3_X1 U855 ( .A1(n986), .A2(n1163), .A3(KEYINPUT0), .ZN(n1161) );
NAND4_X1 U856 ( .A1(n1010), .A2(n991), .A3(n1135), .A4(n1159), .ZN(n1163) );
INV_X1 U857 ( .A(n1164), .ZN(n986) );
NAND2_X1 U858 ( .A1(n1011), .A2(n1165), .ZN(n1164) );
XNOR2_X1 U859 ( .A(G128), .B(n1122), .ZN(G30) );
NAND3_X1 U860 ( .A1(n992), .A2(n1013), .A3(n1127), .ZN(n1122) );
AND3_X1 U861 ( .A1(n1135), .A2(n1159), .A3(n1146), .ZN(n1127) );
XNOR2_X1 U862 ( .A(G101), .B(n1144), .ZN(G3) );
NAND3_X1 U863 ( .A1(n1010), .A2(n1142), .A3(n993), .ZN(n1144) );
XNOR2_X1 U864 ( .A(G125), .B(n1123), .ZN(G27) );
NAND3_X1 U865 ( .A1(n989), .A2(n1013), .A3(n1156), .ZN(n1123) );
AND4_X1 U866 ( .A1(n1008), .A2(n991), .A3(n1009), .A4(n1159), .ZN(n1156) );
NAND2_X1 U867 ( .A1(n1166), .A2(n1167), .ZN(n1159) );
NAND4_X1 U868 ( .A1(n1168), .A2(G953), .A3(G902), .A4(n981), .ZN(n1167) );
XNOR2_X1 U869 ( .A(G900), .B(KEYINPUT61), .ZN(n1168) );
XNOR2_X1 U870 ( .A(G122), .B(n1143), .ZN(G24) );
NAND4_X1 U871 ( .A1(n1169), .A2(n1147), .A3(n984), .A4(n1170), .ZN(n1143) );
AND2_X1 U872 ( .A1(n989), .A2(n1152), .ZN(n1170) );
NOR2_X1 U873 ( .A1(n1009), .A2(n1171), .ZN(n984) );
XNOR2_X1 U874 ( .A(G119), .B(n1172), .ZN(G21) );
NAND4_X1 U875 ( .A1(n1173), .A2(n993), .A3(n1146), .A4(n1147), .ZN(n1172) );
AND2_X1 U876 ( .A1(n1174), .A2(n1009), .ZN(n1146) );
XNOR2_X1 U877 ( .A(n1171), .B(KEYINPUT32), .ZN(n1174) );
XNOR2_X1 U878 ( .A(n989), .B(KEYINPUT55), .ZN(n1173) );
XOR2_X1 U879 ( .A(G116), .B(n1141), .Z(G18) );
AND2_X1 U880 ( .A1(n1175), .A2(n992), .ZN(n1141) );
NOR2_X1 U881 ( .A1(n1155), .A2(n1152), .ZN(n992) );
XOR2_X1 U882 ( .A(n1140), .B(n1176), .Z(G15) );
NOR2_X1 U883 ( .A1(KEYINPUT12), .A2(n1177), .ZN(n1176) );
AND2_X1 U884 ( .A1(n1175), .A2(n991), .ZN(n1140) );
AND2_X1 U885 ( .A1(n1152), .A2(n1155), .ZN(n991) );
AND3_X1 U886 ( .A1(n989), .A2(n1147), .A3(n1010), .ZN(n1175) );
NOR2_X1 U887 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
INV_X1 U888 ( .A(n998), .ZN(n989) );
NAND2_X1 U889 ( .A1(n1000), .A2(n1178), .ZN(n998) );
XNOR2_X1 U890 ( .A(G110), .B(n1179), .ZN(G12) );
NAND2_X1 U891 ( .A1(KEYINPUT62), .A2(n1139), .ZN(n1179) );
AND4_X1 U892 ( .A1(n993), .A2(n1142), .A3(n1008), .A4(n1009), .ZN(n1139) );
XNOR2_X1 U893 ( .A(n1180), .B(n1181), .ZN(n1009) );
NOR2_X1 U894 ( .A1(G902), .A2(n1075), .ZN(n1181) );
XNOR2_X1 U895 ( .A(n1182), .B(n1183), .ZN(n1075) );
XOR2_X1 U896 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U897 ( .A(G119), .B(n1108), .ZN(n1185) );
NOR3_X1 U898 ( .A1(n1186), .A2(KEYINPUT31), .A3(n1187), .ZN(n1184) );
NOR2_X1 U899 ( .A1(n1188), .A2(n1051), .ZN(n1187) );
AND2_X1 U900 ( .A1(n1189), .A2(G221), .ZN(n1188) );
XOR2_X1 U901 ( .A(n1190), .B(KEYINPUT25), .Z(n1186) );
NAND3_X1 U902 ( .A1(n1189), .A2(n1051), .A3(G221), .ZN(n1190) );
INV_X1 U903 ( .A(n1191), .ZN(n1189) );
XNOR2_X1 U904 ( .A(n1192), .B(n1193), .ZN(n1182) );
NAND2_X1 U905 ( .A1(G217), .A2(n1194), .ZN(n1180) );
XOR2_X1 U906 ( .A(KEYINPUT43), .B(n1195), .Z(n1194) );
AND2_X1 U907 ( .A1(n1196), .A2(G234), .ZN(n1195) );
INV_X1 U908 ( .A(n1171), .ZN(n1008) );
XOR2_X1 U909 ( .A(n1197), .B(n1100), .Z(n1171) );
INV_X1 U910 ( .A(G472), .ZN(n1100) );
NAND2_X1 U911 ( .A1(n1198), .A2(n1196), .ZN(n1197) );
XOR2_X1 U912 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U913 ( .A(n1096), .B(n1101), .ZN(n1200) );
XNOR2_X1 U914 ( .A(n1052), .B(n1201), .ZN(n1101) );
XNOR2_X1 U915 ( .A(n1202), .B(n1203), .ZN(n1096) );
XOR2_X1 U916 ( .A(G101), .B(n1204), .Z(n1203) );
XNOR2_X1 U917 ( .A(KEYINPUT27), .B(n1177), .ZN(n1204) );
INV_X1 U918 ( .A(G113), .ZN(n1177) );
XOR2_X1 U919 ( .A(n1205), .B(n1206), .Z(n1202) );
NAND3_X1 U920 ( .A1(n1207), .A2(n975), .A3(G210), .ZN(n1205) );
XOR2_X1 U921 ( .A(KEYINPUT16), .B(n1208), .Z(n1199) );
XOR2_X1 U922 ( .A(KEYINPUT35), .B(KEYINPUT21), .Z(n1208) );
AND2_X1 U923 ( .A1(n1147), .A2(n1135), .ZN(n1142) );
NOR2_X1 U924 ( .A1(n1000), .A2(n999), .ZN(n1135) );
INV_X1 U925 ( .A(n1178), .ZN(n999) );
NAND2_X1 U926 ( .A1(G221), .A2(n1209), .ZN(n1178) );
NAND2_X1 U927 ( .A1(G234), .A2(n1196), .ZN(n1209) );
XNOR2_X1 U928 ( .A(n1210), .B(n1112), .ZN(n1000) );
INV_X1 U929 ( .A(G469), .ZN(n1112) );
NAND2_X1 U930 ( .A1(n1211), .A2(n1196), .ZN(n1210) );
XOR2_X1 U931 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U932 ( .A(n1214), .B(n1215), .Z(n1213) );
NAND2_X1 U933 ( .A1(KEYINPUT13), .A2(n1201), .ZN(n1215) );
XNOR2_X1 U934 ( .A(n1051), .B(n1216), .ZN(n1201) );
XNOR2_X1 U935 ( .A(n1046), .B(n1217), .ZN(n1216) );
NOR2_X1 U936 ( .A1(G131), .A2(KEYINPUT8), .ZN(n1217) );
INV_X1 U937 ( .A(G134), .ZN(n1046) );
XOR2_X1 U938 ( .A(G137), .B(KEYINPUT22), .Z(n1051) );
NAND2_X1 U939 ( .A1(n1218), .A2(n1219), .ZN(n1214) );
XNOR2_X1 U940 ( .A(n1108), .B(n1220), .ZN(n1219) );
XOR2_X1 U941 ( .A(KEYINPUT56), .B(G140), .Z(n1220) );
XNOR2_X1 U942 ( .A(KEYINPUT58), .B(KEYINPUT4), .ZN(n1218) );
XNOR2_X1 U943 ( .A(n1111), .B(n1221), .ZN(n1212) );
NAND2_X1 U944 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U945 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U946 ( .A(n1226), .B(KEYINPUT36), .Z(n1222) );
NAND2_X1 U947 ( .A1(n1052), .A2(n1107), .ZN(n1226) );
INV_X1 U948 ( .A(n1225), .ZN(n1052) );
AND2_X1 U949 ( .A1(G227), .A2(n975), .ZN(n1111) );
AND2_X1 U950 ( .A1(n1013), .A2(n1227), .ZN(n1147) );
NAND2_X1 U951 ( .A1(n1228), .A2(n1166), .ZN(n1227) );
NAND3_X1 U952 ( .A1(n1229), .A2(n975), .A3(G952), .ZN(n1166) );
XNOR2_X1 U953 ( .A(KEYINPUT50), .B(n981), .ZN(n1229) );
XOR2_X1 U954 ( .A(n1230), .B(KEYINPUT51), .Z(n1228) );
NAND4_X1 U955 ( .A1(G953), .A2(G902), .A3(n981), .A4(n1067), .ZN(n1230) );
INV_X1 U956 ( .A(G898), .ZN(n1067) );
NAND2_X1 U957 ( .A1(G237), .A2(G234), .ZN(n981) );
NOR2_X1 U958 ( .A1(n1011), .A2(n1012), .ZN(n1013) );
INV_X1 U959 ( .A(n1165), .ZN(n1012) );
NAND2_X1 U960 ( .A1(G214), .A2(n1231), .ZN(n1165) );
XNOR2_X1 U961 ( .A(n1022), .B(n1021), .ZN(n1011) );
NAND2_X1 U962 ( .A1(G210), .A2(n1231), .ZN(n1021) );
NAND2_X1 U963 ( .A1(n1207), .A2(n1196), .ZN(n1231) );
NAND2_X1 U964 ( .A1(n1232), .A2(n1196), .ZN(n1022) );
INV_X1 U965 ( .A(G902), .ZN(n1196) );
XOR2_X1 U966 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U967 ( .A(n1119), .B(n1235), .ZN(n1234) );
NAND3_X1 U968 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
OR2_X1 U969 ( .A1(n1225), .A2(KEYINPUT11), .ZN(n1238) );
NAND3_X1 U970 ( .A1(KEYINPUT11), .A2(n1225), .A3(G125), .ZN(n1237) );
NAND2_X1 U971 ( .A1(n1239), .A2(n1045), .ZN(n1236) );
NAND2_X1 U972 ( .A1(n1240), .A2(KEYINPUT11), .ZN(n1239) );
XNOR2_X1 U973 ( .A(n1225), .B(KEYINPUT1), .ZN(n1240) );
XNOR2_X1 U974 ( .A(n1241), .B(n1192), .ZN(n1225) );
XOR2_X1 U975 ( .A(G146), .B(n1242), .Z(n1192) );
XNOR2_X1 U976 ( .A(G143), .B(KEYINPUT44), .ZN(n1241) );
NOR2_X1 U977 ( .A1(n1059), .A2(G953), .ZN(n1119) );
INV_X1 U978 ( .A(G224), .ZN(n1059) );
NAND2_X1 U979 ( .A1(KEYINPUT20), .A2(n1116), .ZN(n1233) );
XNOR2_X1 U980 ( .A(n1068), .B(n1243), .ZN(n1116) );
XNOR2_X1 U981 ( .A(KEYINPUT59), .B(n1071), .ZN(n1243) );
XNOR2_X1 U982 ( .A(n1108), .B(n1244), .ZN(n1071) );
INV_X1 U983 ( .A(G110), .ZN(n1108) );
XOR2_X1 U984 ( .A(n1245), .B(n1206), .Z(n1068) );
XOR2_X1 U985 ( .A(G116), .B(G119), .Z(n1206) );
XNOR2_X1 U986 ( .A(n1246), .B(n1224), .ZN(n1245) );
INV_X1 U987 ( .A(n1107), .ZN(n1224) );
XOR2_X1 U988 ( .A(G101), .B(n1247), .Z(n1107) );
XOR2_X1 U989 ( .A(G107), .B(G104), .Z(n1247) );
NAND2_X1 U990 ( .A1(KEYINPUT26), .A2(G113), .ZN(n1246) );
NOR2_X1 U991 ( .A1(n1169), .A2(n1152), .ZN(n993) );
XNOR2_X1 U992 ( .A(n1248), .B(n1249), .ZN(n1152) );
INV_X1 U993 ( .A(n1026), .ZN(n1249) );
NOR2_X1 U994 ( .A1(n1087), .A2(G902), .ZN(n1026) );
INV_X1 U995 ( .A(n1084), .ZN(n1087) );
XNOR2_X1 U996 ( .A(n1250), .B(n1251), .ZN(n1084) );
XNOR2_X1 U997 ( .A(n1193), .B(n1252), .ZN(n1251) );
XNOR2_X1 U998 ( .A(n1253), .B(n1254), .ZN(n1252) );
NAND2_X1 U999 ( .A1(KEYINPUT49), .A2(G104), .ZN(n1254) );
NAND2_X1 U1000 ( .A1(KEYINPUT46), .A2(n1255), .ZN(n1253) );
NAND2_X1 U1001 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND3_X1 U1002 ( .A1(n1258), .A2(n1259), .A3(G131), .ZN(n1257) );
XOR2_X1 U1003 ( .A(KEYINPUT42), .B(n1260), .Z(n1256) );
NOR2_X1 U1004 ( .A1(G131), .A2(n1261), .ZN(n1260) );
AND2_X1 U1005 ( .A1(n1258), .A2(n1259), .ZN(n1261) );
NAND2_X1 U1006 ( .A1(G143), .A2(n1262), .ZN(n1259) );
XOR2_X1 U1007 ( .A(KEYINPUT53), .B(n1263), .Z(n1262) );
NAND2_X1 U1008 ( .A1(n1263), .A2(n1150), .ZN(n1258) );
AND3_X1 U1009 ( .A1(n1207), .A2(n975), .A3(G214), .ZN(n1263) );
INV_X1 U1010 ( .A(G237), .ZN(n1207) );
XNOR2_X1 U1011 ( .A(G140), .B(n1045), .ZN(n1193) );
INV_X1 U1012 ( .A(G125), .ZN(n1045) );
XOR2_X1 U1013 ( .A(n1264), .B(n1265), .Z(n1250) );
XNOR2_X1 U1014 ( .A(n1244), .B(G113), .ZN(n1265) );
XNOR2_X1 U1015 ( .A(G146), .B(KEYINPUT41), .ZN(n1264) );
NAND2_X1 U1016 ( .A1(KEYINPUT40), .A2(n1085), .ZN(n1248) );
INV_X1 U1017 ( .A(G475), .ZN(n1085) );
INV_X1 U1018 ( .A(n1155), .ZN(n1169) );
XOR2_X1 U1019 ( .A(n1266), .B(n1024), .Z(n1155) );
INV_X1 U1020 ( .A(G478), .ZN(n1024) );
NAND2_X1 U1021 ( .A1(KEYINPUT3), .A2(n1267), .ZN(n1266) );
INV_X1 U1022 ( .A(n1025), .ZN(n1267) );
NOR2_X1 U1023 ( .A1(n1268), .A2(G902), .ZN(n1025) );
INV_X1 U1024 ( .A(n1079), .ZN(n1268) );
XNOR2_X1 U1025 ( .A(n1269), .B(n1270), .ZN(n1079) );
XOR2_X1 U1026 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U1027 ( .A1(G107), .A2(KEYINPUT47), .ZN(n1272) );
NOR2_X1 U1028 ( .A1(n1191), .A2(n1076), .ZN(n1271) );
INV_X1 U1029 ( .A(G217), .ZN(n1076) );
NAND2_X1 U1030 ( .A1(G234), .A2(n975), .ZN(n1191) );
INV_X1 U1031 ( .A(G953), .ZN(n975) );
XOR2_X1 U1032 ( .A(n1273), .B(n1274), .Z(n1269) );
XNOR2_X1 U1033 ( .A(n1244), .B(G116), .ZN(n1274) );
INV_X1 U1034 ( .A(G122), .ZN(n1244) );
NAND2_X1 U1035 ( .A1(n1275), .A2(KEYINPUT10), .ZN(n1273) );
XNOR2_X1 U1036 ( .A(G134), .B(n1276), .ZN(n1275) );
NOR2_X1 U1037 ( .A1(KEYINPUT48), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U1038 ( .A(n1150), .B(n1242), .ZN(n1277) );
XOR2_X1 U1039 ( .A(G128), .B(KEYINPUT45), .Z(n1242) );
INV_X1 U1040 ( .A(G143), .ZN(n1150) );
endmodule


