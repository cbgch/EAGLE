//Key = 0011100001010110100101111010111001110101000111000110110110111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;

XOR2_X1 U740 ( .A(G107), .B(n1025), .Z(G9) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(G75) );
XOR2_X1 U742 ( .A(KEYINPUT6), .B(n1028), .Z(n1027) );
AND3_X1 U743 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR4_X1 U744 ( .A1(n1032), .A2(n1033), .A3(n1030), .A4(n1034), .ZN(n1026) );
INV_X1 U745 ( .A(G952), .ZN(n1030) );
NAND3_X1 U746 ( .A1(n1035), .A2(n1031), .A3(n1036), .ZN(n1032) );
NAND2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
INV_X1 U750 ( .A(KEYINPUT4), .ZN(n1043) );
NAND4_X1 U751 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1042) );
NAND3_X1 U752 ( .A1(n1045), .A2(n1048), .A3(n1044), .ZN(n1040) );
NAND3_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1052), .ZN(n1051) );
NAND3_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U756 ( .A1(KEYINPUT4), .A2(n1046), .ZN(n1055) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND2_X1 U758 ( .A1(KEYINPUT19), .A2(KEYINPUT39), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1056), .A2(n1058), .ZN(n1050) );
NAND2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U761 ( .A1(KEYINPUT19), .A2(n1061), .A3(n1062), .ZN(n1060) );
NAND2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
INV_X1 U763 ( .A(KEYINPUT48), .ZN(n1064) );
NAND3_X1 U764 ( .A1(KEYINPUT48), .A2(n1063), .A3(n1065), .ZN(n1049) );
NAND2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1039) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND4_X1 U767 ( .A1(n1070), .A2(n1037), .A3(n1071), .A4(n1072), .ZN(n1031) );
NOR4_X1 U768 ( .A1(n1062), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XOR2_X1 U769 ( .A(G478), .B(n1076), .Z(n1071) );
NAND3_X1 U770 ( .A1(n1045), .A2(n1077), .A3(n1066), .ZN(n1035) );
AND3_X1 U771 ( .A1(n1047), .A2(n1056), .A3(n1044), .ZN(n1066) );
INV_X1 U772 ( .A(n1078), .ZN(n1044) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND3_X1 U774 ( .A1(n1081), .A2(n1082), .A3(KEYINPUT39), .ZN(n1080) );
XOR2_X1 U775 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U777 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1088) );
NOR2_X1 U779 ( .A1(KEYINPUT32), .A2(n1091), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1092), .B(G137), .Z(n1091) );
NAND2_X1 U781 ( .A1(KEYINPUT58), .A2(G134), .ZN(n1092) );
XNOR2_X1 U782 ( .A(n1093), .B(n1094), .ZN(n1087) );
NAND3_X1 U783 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1083) );
INV_X1 U784 ( .A(n1085), .ZN(n1097) );
NAND2_X1 U785 ( .A1(G953), .A2(n1098), .ZN(n1096) );
NAND2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
NAND3_X1 U787 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1104), .B(KEYINPUT1), .Z(n1103) );
NAND2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(G69) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
XOR2_X1 U792 ( .A(n1108), .B(KEYINPUT35), .Z(n1110) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U794 ( .A1(G953), .A2(n1113), .ZN(n1112) );
INV_X1 U795 ( .A(n1107), .ZN(n1109) );
NAND2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(n1107) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U798 ( .A(n1118), .B(KEYINPUT47), .Z(n1116) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
INV_X1 U800 ( .A(n1117), .ZN(n1120) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1111), .ZN(n1117) );
INV_X1 U802 ( .A(n1122), .ZN(n1111) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1121) );
NAND2_X1 U804 ( .A1(KEYINPUT2), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U805 ( .A(KEYINPUT17), .B(n1118), .ZN(n1119) );
NAND2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1118) );
XNOR2_X1 U807 ( .A(G953), .B(KEYINPUT15), .ZN(n1126) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(G63) );
XNOR2_X1 U812 ( .A(n1128), .B(KEYINPUT13), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1136), .B(n1137), .Z(n1134) );
NOR2_X1 U814 ( .A1(KEYINPUT46), .A2(n1138), .ZN(n1137) );
NAND3_X1 U815 ( .A1(n1139), .A2(n1033), .A3(G478), .ZN(n1136) );
XNOR2_X1 U816 ( .A(KEYINPUT20), .B(n1140), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1128), .A2(n1141), .ZN(G60) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR3_X1 U819 ( .A1(n1133), .A2(KEYINPUT18), .A3(n1144), .ZN(n1142) );
XOR2_X1 U820 ( .A(G104), .B(n1145), .Z(G6) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(G57) );
XNOR2_X1 U822 ( .A(n1148), .B(n1149), .ZN(n1147) );
NAND2_X1 U823 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NAND2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1150) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1133), .ZN(n1155) );
OR2_X1 U827 ( .A1(n1153), .A2(n1152), .ZN(n1154) );
XNOR2_X1 U828 ( .A(n1157), .B(n1158), .ZN(n1152) );
XOR2_X1 U829 ( .A(KEYINPUT38), .B(KEYINPUT30), .Z(n1158) );
XOR2_X1 U830 ( .A(n1159), .B(n1160), .Z(n1157) );
INV_X1 U831 ( .A(KEYINPUT26), .ZN(n1153) );
NOR2_X1 U832 ( .A1(n1161), .A2(n1100), .ZN(n1146) );
XNOR2_X1 U833 ( .A(G952), .B(KEYINPUT9), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1128), .A2(n1162), .ZN(G54) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1133), .ZN(n1164) );
NAND2_X1 U837 ( .A1(KEYINPUT50), .A2(n1166), .ZN(n1163) );
XOR2_X1 U838 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U839 ( .A(n1169), .B(n1170), .ZN(n1168) );
XNOR2_X1 U840 ( .A(n1171), .B(G140), .ZN(n1167) );
NOR2_X1 U841 ( .A1(n1100), .A2(G952), .ZN(n1128) );
NOR2_X1 U842 ( .A1(n1172), .A2(n1173), .ZN(G51) );
XOR2_X1 U843 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U845 ( .A1(n1178), .A2(n1133), .ZN(n1176) );
NAND2_X1 U846 ( .A1(G902), .A2(n1033), .ZN(n1133) );
NAND4_X1 U847 ( .A1(n1179), .A2(n1180), .A3(n1101), .A4(n1104), .ZN(n1033) );
AND4_X1 U848 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1101) );
AND3_X1 U849 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
INV_X1 U850 ( .A(n1127), .ZN(n1180) );
NAND4_X1 U851 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1127) );
NOR4_X1 U852 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NOR2_X1 U853 ( .A1(n1079), .A2(n1196), .ZN(n1195) );
NOR3_X1 U854 ( .A1(n1197), .A2(n1054), .A3(n1198), .ZN(n1194) );
INV_X1 U855 ( .A(n1199), .ZN(n1054) );
INV_X1 U856 ( .A(n1200), .ZN(n1193) );
NOR2_X1 U857 ( .A1(n1145), .A2(n1025), .ZN(n1190) );
NOR3_X1 U858 ( .A1(n1069), .A2(n1065), .A3(n1198), .ZN(n1025) );
NOR3_X1 U859 ( .A1(n1198), .A2(n1065), .A3(n1068), .ZN(n1145) );
XOR2_X1 U860 ( .A(n1102), .B(KEYINPUT8), .Z(n1179) );
NAND3_X1 U861 ( .A1(n1046), .A2(n1201), .A3(n1202), .ZN(n1102) );
XOR2_X1 U862 ( .A(n1203), .B(KEYINPUT21), .Z(n1174) );
NAND3_X1 U863 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NAND2_X1 U864 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U865 ( .A(KEYINPUT0), .ZN(n1208) );
NAND2_X1 U866 ( .A1(KEYINPUT0), .A2(n1209), .ZN(n1204) );
NOR2_X1 U867 ( .A1(G952), .A2(n1210), .ZN(n1172) );
XNOR2_X1 U868 ( .A(KEYINPUT44), .B(n1100), .ZN(n1210) );
XNOR2_X1 U869 ( .A(G146), .B(n1183), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1063), .A2(n1211), .A3(n1212), .ZN(n1183) );
XOR2_X1 U871 ( .A(n1186), .B(n1213), .Z(G45) );
NAND2_X1 U872 ( .A1(KEYINPUT28), .A2(G143), .ZN(n1213) );
NAND4_X1 U873 ( .A1(n1214), .A2(n1046), .A3(n1063), .A4(n1215), .ZN(n1186) );
NOR3_X1 U874 ( .A1(n1079), .A2(n1216), .A3(n1217), .ZN(n1215) );
XNOR2_X1 U875 ( .A(G140), .B(n1181), .ZN(G42) );
NAND3_X1 U876 ( .A1(n1201), .A2(n1199), .A3(n1202), .ZN(n1181) );
XNOR2_X1 U877 ( .A(G137), .B(n1182), .ZN(G39) );
NAND4_X1 U878 ( .A1(n1202), .A2(n1045), .A3(n1218), .A4(n1219), .ZN(n1182) );
XNOR2_X1 U879 ( .A(G134), .B(n1185), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1046), .A2(n1220), .A3(n1202), .ZN(n1185) );
AND3_X1 U881 ( .A1(n1063), .A2(n1221), .A3(n1037), .ZN(n1202) );
XNOR2_X1 U882 ( .A(n1089), .B(n1222), .ZN(G33) );
AND4_X1 U883 ( .A1(n1223), .A2(n1046), .A3(n1212), .A4(n1037), .ZN(n1222) );
NOR2_X1 U884 ( .A1(n1224), .A2(n1082), .ZN(n1037) );
XNOR2_X1 U885 ( .A(n1063), .B(KEYINPUT43), .ZN(n1223) );
XNOR2_X1 U886 ( .A(n1225), .B(KEYINPUT22), .ZN(n1063) );
XNOR2_X1 U887 ( .A(G128), .B(n1104), .ZN(G30) );
NAND4_X1 U888 ( .A1(n1211), .A2(n1220), .A3(n1225), .A4(n1221), .ZN(n1104) );
XNOR2_X1 U889 ( .A(n1226), .B(n1188), .ZN(G3) );
OR3_X1 U890 ( .A1(n1227), .A2(n1198), .A3(n1197), .ZN(n1188) );
INV_X1 U891 ( .A(n1045), .ZN(n1197) );
NAND2_X1 U892 ( .A1(KEYINPUT16), .A2(n1228), .ZN(n1226) );
INV_X1 U893 ( .A(G101), .ZN(n1228) );
XNOR2_X1 U894 ( .A(G125), .B(n1187), .ZN(G27) );
NAND4_X1 U895 ( .A1(n1212), .A2(n1047), .A3(n1199), .A4(n1229), .ZN(n1187) );
NOR2_X1 U896 ( .A1(n1068), .A2(n1216), .ZN(n1212) );
INV_X1 U897 ( .A(n1221), .ZN(n1216) );
NAND2_X1 U898 ( .A1(n1230), .A2(n1078), .ZN(n1221) );
NAND3_X1 U899 ( .A1(G902), .A2(n1231), .A3(n1085), .ZN(n1230) );
NOR2_X1 U900 ( .A1(G900), .A2(n1100), .ZN(n1085) );
INV_X1 U901 ( .A(n1201), .ZN(n1068) );
XNOR2_X1 U902 ( .A(G122), .B(n1200), .ZN(G24) );
NAND3_X1 U903 ( .A1(n1214), .A2(n1232), .A3(n1233), .ZN(n1200) );
NOR3_X1 U904 ( .A1(n1079), .A2(n1065), .A3(n1217), .ZN(n1233) );
INV_X1 U905 ( .A(n1056), .ZN(n1065) );
NAND2_X1 U906 ( .A1(n1234), .A2(n1235), .ZN(n1056) );
OR3_X1 U907 ( .A1(n1074), .A2(n1219), .A3(KEYINPUT10), .ZN(n1235) );
NAND2_X1 U908 ( .A1(KEYINPUT10), .A2(n1199), .ZN(n1234) );
XOR2_X1 U909 ( .A(G119), .B(n1192), .Z(G21) );
AND3_X1 U910 ( .A1(n1232), .A2(n1211), .A3(n1045), .ZN(n1192) );
AND3_X1 U911 ( .A1(n1218), .A2(n1219), .A3(n1229), .ZN(n1211) );
XNOR2_X1 U912 ( .A(n1236), .B(n1237), .ZN(G18) );
NOR2_X1 U913 ( .A1(n1238), .A2(n1079), .ZN(n1237) );
XOR2_X1 U914 ( .A(n1196), .B(KEYINPUT27), .Z(n1238) );
NAND3_X1 U915 ( .A1(n1232), .A2(n1220), .A3(n1046), .ZN(n1196) );
INV_X1 U916 ( .A(n1069), .ZN(n1220) );
NAND2_X1 U917 ( .A1(n1239), .A2(n1214), .ZN(n1069) );
XNOR2_X1 U918 ( .A(n1075), .B(KEYINPUT40), .ZN(n1239) );
XNOR2_X1 U919 ( .A(G113), .B(n1189), .ZN(G15) );
NAND4_X1 U920 ( .A1(n1046), .A2(n1201), .A3(n1232), .A4(n1229), .ZN(n1189) );
AND2_X1 U921 ( .A1(n1047), .A2(n1240), .ZN(n1232) );
AND2_X1 U922 ( .A1(n1061), .A2(n1241), .ZN(n1047) );
NOR2_X1 U923 ( .A1(n1217), .A2(n1214), .ZN(n1201) );
INV_X1 U924 ( .A(n1075), .ZN(n1217) );
INV_X1 U925 ( .A(n1227), .ZN(n1046) );
NAND2_X1 U926 ( .A1(n1242), .A2(n1218), .ZN(n1227) );
XOR2_X1 U927 ( .A(n1074), .B(KEYINPUT57), .Z(n1218) );
XNOR2_X1 U928 ( .A(n1219), .B(KEYINPUT10), .ZN(n1242) );
XNOR2_X1 U929 ( .A(G110), .B(n1243), .ZN(G12) );
NAND4_X1 U930 ( .A1(n1045), .A2(n1199), .A3(n1244), .A4(n1245), .ZN(n1243) );
NAND2_X1 U931 ( .A1(n1198), .A2(n1246), .ZN(n1245) );
INV_X1 U932 ( .A(KEYINPUT42), .ZN(n1246) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1247), .ZN(n1198) );
NAND2_X1 U934 ( .A1(KEYINPUT42), .A2(n1248), .ZN(n1244) );
NAND2_X1 U935 ( .A1(n1247), .A2(n1079), .ZN(n1248) );
INV_X1 U936 ( .A(n1229), .ZN(n1079) );
NOR2_X1 U937 ( .A1(n1081), .A2(n1082), .ZN(n1229) );
AND2_X1 U938 ( .A1(G214), .A2(n1249), .ZN(n1082) );
INV_X1 U939 ( .A(n1224), .ZN(n1081) );
XOR2_X1 U940 ( .A(n1250), .B(n1178), .Z(n1224) );
NAND2_X1 U941 ( .A1(G210), .A2(n1249), .ZN(n1178) );
NAND2_X1 U942 ( .A1(n1251), .A2(n1140), .ZN(n1249) );
INV_X1 U943 ( .A(G237), .ZN(n1251) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1140), .ZN(n1250) );
XNOR2_X1 U945 ( .A(n1177), .B(n1253), .ZN(n1252) );
NOR2_X1 U946 ( .A1(n1207), .A2(n1254), .ZN(n1253) );
INV_X1 U947 ( .A(n1206), .ZN(n1254) );
NAND2_X1 U948 ( .A1(n1209), .A2(n1255), .ZN(n1206) );
NOR2_X1 U949 ( .A1(n1255), .A2(n1209), .ZN(n1207) );
NOR2_X1 U950 ( .A1(n1113), .A2(G953), .ZN(n1209) );
INV_X1 U951 ( .A(G224), .ZN(n1113) );
XOR2_X1 U952 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U953 ( .A(n1124), .B(n1125), .Z(n1177) );
XOR2_X1 U954 ( .A(n1236), .B(n1258), .Z(n1125) );
XOR2_X1 U955 ( .A(n1259), .B(n1260), .Z(n1124) );
XNOR2_X1 U956 ( .A(KEYINPUT45), .B(n1261), .ZN(n1260) );
XOR2_X1 U957 ( .A(n1262), .B(n1263), .Z(n1259) );
NOR2_X1 U958 ( .A1(G122), .A2(KEYINPUT54), .ZN(n1263) );
AND2_X1 U959 ( .A1(n1225), .A2(n1240), .ZN(n1247) );
NAND2_X1 U960 ( .A1(n1078), .A2(n1264), .ZN(n1240) );
NAND3_X1 U961 ( .A1(n1122), .A2(n1231), .A3(G902), .ZN(n1264) );
NOR2_X1 U962 ( .A1(G898), .A2(n1100), .ZN(n1122) );
NAND3_X1 U963 ( .A1(n1029), .A2(n1231), .A3(G952), .ZN(n1078) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1231) );
INV_X1 U965 ( .A(n1034), .ZN(n1029) );
XOR2_X1 U966 ( .A(G953), .B(KEYINPUT7), .Z(n1034) );
NOR2_X1 U967 ( .A1(n1061), .A2(n1062), .ZN(n1225) );
INV_X1 U968 ( .A(n1241), .ZN(n1062) );
NAND2_X1 U969 ( .A1(G221), .A2(n1265), .ZN(n1241) );
XOR2_X1 U970 ( .A(n1073), .B(KEYINPUT59), .Z(n1061) );
XOR2_X1 U971 ( .A(n1266), .B(n1165), .Z(n1073) );
INV_X1 U972 ( .A(G469), .ZN(n1165) );
NAND2_X1 U973 ( .A1(n1267), .A2(n1140), .ZN(n1266) );
XOR2_X1 U974 ( .A(n1268), .B(n1170), .Z(n1267) );
XNOR2_X1 U975 ( .A(n1261), .B(n1269), .ZN(n1170) );
NOR2_X1 U976 ( .A1(G953), .A2(n1098), .ZN(n1269) );
INV_X1 U977 ( .A(G227), .ZN(n1098) );
XOR2_X1 U978 ( .A(n1270), .B(n1271), .Z(n1268) );
NOR2_X1 U979 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U980 ( .A(n1274), .B(KEYINPUT29), .Z(n1273) );
NAND2_X1 U981 ( .A1(n1169), .A2(n1171), .ZN(n1274) );
NOR2_X1 U982 ( .A1(n1169), .A2(n1171), .ZN(n1272) );
XNOR2_X1 U983 ( .A(n1262), .B(n1275), .ZN(n1169) );
XOR2_X1 U984 ( .A(KEYINPUT55), .B(n1094), .Z(n1275) );
XNOR2_X1 U985 ( .A(n1276), .B(n1277), .ZN(n1094) );
XOR2_X1 U986 ( .A(KEYINPUT37), .B(G128), .Z(n1277) );
NAND2_X1 U987 ( .A1(KEYINPUT60), .A2(n1278), .ZN(n1276) );
XOR2_X1 U988 ( .A(G143), .B(n1279), .Z(n1278) );
XNOR2_X1 U989 ( .A(G101), .B(n1280), .ZN(n1262) );
XOR2_X1 U990 ( .A(G107), .B(G104), .Z(n1280) );
NAND2_X1 U991 ( .A1(KEYINPUT23), .A2(n1281), .ZN(n1270) );
XOR2_X1 U992 ( .A(KEYINPUT11), .B(G140), .Z(n1281) );
NOR2_X1 U993 ( .A1(n1074), .A2(n1070), .ZN(n1199) );
INV_X1 U994 ( .A(n1219), .ZN(n1070) );
XOR2_X1 U995 ( .A(n1282), .B(n1132), .Z(n1219) );
NAND2_X1 U996 ( .A1(G217), .A2(n1265), .ZN(n1132) );
NAND2_X1 U997 ( .A1(G234), .A2(n1140), .ZN(n1265) );
OR2_X1 U998 ( .A1(n1131), .A2(G902), .ZN(n1282) );
XNOR2_X1 U999 ( .A(n1283), .B(n1284), .ZN(n1131) );
XOR2_X1 U1000 ( .A(G137), .B(n1285), .Z(n1284) );
NOR2_X1 U1001 ( .A1(KEYINPUT62), .A2(n1286), .ZN(n1285) );
XOR2_X1 U1002 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1003 ( .A(G128), .B(G119), .Z(n1288) );
XNOR2_X1 U1004 ( .A(n1289), .B(n1290), .ZN(n1287) );
NAND2_X1 U1005 ( .A1(KEYINPUT14), .A2(n1261), .ZN(n1290) );
INV_X1 U1006 ( .A(G110), .ZN(n1261) );
NAND3_X1 U1007 ( .A1(n1291), .A2(n1292), .A3(KEYINPUT63), .ZN(n1289) );
NAND2_X1 U1008 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n1295), .Z(n1291) );
NOR2_X1 U1010 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
NAND2_X1 U1011 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
OR2_X1 U1012 ( .A1(n1093), .A2(KEYINPUT51), .ZN(n1297) );
NAND3_X1 U1013 ( .A1(G140), .A2(n1256), .A3(KEYINPUT51), .ZN(n1296) );
INV_X1 U1014 ( .A(G125), .ZN(n1256) );
NAND2_X1 U1015 ( .A1(n1298), .A2(G221), .ZN(n1283) );
XOR2_X1 U1016 ( .A(n1299), .B(n1156), .Z(n1074) );
INV_X1 U1017 ( .A(G472), .ZN(n1156) );
NAND2_X1 U1018 ( .A1(n1140), .A2(n1300), .ZN(n1299) );
NAND2_X1 U1019 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1020 ( .A1(n1149), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1021 ( .A(n1304), .B(KEYINPUT41), .Z(n1301) );
NAND2_X1 U1022 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XNOR2_X1 U1023 ( .A(KEYINPUT25), .B(n1149), .ZN(n1306) );
XOR2_X1 U1024 ( .A(n1307), .B(G101), .Z(n1149) );
NAND2_X1 U1025 ( .A1(n1308), .A2(G210), .ZN(n1307) );
INV_X1 U1026 ( .A(n1303), .ZN(n1305) );
XNOR2_X1 U1027 ( .A(n1309), .B(n1159), .ZN(n1303) );
XOR2_X1 U1028 ( .A(n1171), .B(n1257), .Z(n1159) );
XNOR2_X1 U1029 ( .A(n1310), .B(n1279), .ZN(n1257) );
XNOR2_X1 U1030 ( .A(n1294), .B(KEYINPUT12), .ZN(n1279) );
XOR2_X1 U1031 ( .A(G131), .B(n1311), .Z(n1171) );
XOR2_X1 U1032 ( .A(G137), .B(G134), .Z(n1311) );
NAND2_X1 U1033 ( .A1(KEYINPUT34), .A2(n1160), .ZN(n1309) );
XOR2_X1 U1034 ( .A(n1312), .B(n1258), .Z(n1160) );
XOR2_X1 U1035 ( .A(G113), .B(G119), .Z(n1258) );
NAND2_X1 U1036 ( .A1(KEYINPUT33), .A2(n1236), .ZN(n1312) );
INV_X1 U1037 ( .A(G902), .ZN(n1140) );
NOR2_X1 U1038 ( .A1(n1075), .A2(n1214), .ZN(n1045) );
XOR2_X1 U1039 ( .A(n1313), .B(G478), .Z(n1214) );
NAND2_X1 U1040 ( .A1(KEYINPUT61), .A2(n1076), .ZN(n1313) );
OR2_X1 U1041 ( .A1(n1138), .A2(G902), .ZN(n1076) );
XOR2_X1 U1042 ( .A(n1314), .B(n1315), .Z(n1138) );
XOR2_X1 U1043 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND3_X1 U1044 ( .A1(G217), .A2(n1298), .A3(KEYINPUT24), .ZN(n1317) );
AND2_X1 U1045 ( .A1(G234), .A2(n1100), .ZN(n1298) );
INV_X1 U1046 ( .A(G953), .ZN(n1100) );
NAND2_X1 U1047 ( .A1(KEYINPUT3), .A2(n1236), .ZN(n1316) );
INV_X1 U1048 ( .A(G116), .ZN(n1236) );
XOR2_X1 U1049 ( .A(n1318), .B(n1319), .Z(n1314) );
NOR2_X1 U1050 ( .A1(KEYINPUT36), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1051 ( .A(G134), .B(n1310), .ZN(n1320) );
XNOR2_X1 U1052 ( .A(G128), .B(G143), .ZN(n1310) );
XNOR2_X1 U1053 ( .A(G107), .B(G122), .ZN(n1318) );
XNOR2_X1 U1054 ( .A(n1321), .B(n1322), .ZN(n1075) );
XNOR2_X1 U1055 ( .A(KEYINPUT31), .B(n1144), .ZN(n1322) );
INV_X1 U1056 ( .A(G475), .ZN(n1144) );
OR2_X1 U1057 ( .A1(n1143), .A2(G902), .ZN(n1321) );
XNOR2_X1 U1058 ( .A(n1323), .B(n1324), .ZN(n1143) );
XOR2_X1 U1059 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1060 ( .A(G104), .B(n1327), .Z(n1326) );
NOR2_X1 U1061 ( .A1(KEYINPUT5), .A2(n1328), .ZN(n1327) );
XNOR2_X1 U1062 ( .A(n1294), .B(n1093), .ZN(n1328) );
XOR2_X1 U1063 ( .A(G125), .B(G140), .Z(n1093) );
INV_X1 U1064 ( .A(G146), .ZN(n1294) );
XOR2_X1 U1065 ( .A(G143), .B(G113), .Z(n1325) );
XOR2_X1 U1066 ( .A(n1329), .B(n1330), .Z(n1323) );
XOR2_X1 U1067 ( .A(n1331), .B(n1332), .Z(n1330) );
NAND2_X1 U1068 ( .A1(KEYINPUT56), .A2(n1333), .ZN(n1332) );
INV_X1 U1069 ( .A(G122), .ZN(n1333) );
NAND2_X1 U1070 ( .A1(KEYINPUT52), .A2(n1089), .ZN(n1331) );
INV_X1 U1071 ( .A(G131), .ZN(n1089) );
NAND3_X1 U1072 ( .A1(n1308), .A2(G214), .A3(KEYINPUT53), .ZN(n1329) );
NOR2_X1 U1073 ( .A1(G953), .A2(G237), .ZN(n1308) );
endmodule


