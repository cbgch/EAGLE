//Key = 1101000101101001101111010110101010011001110000111010111100110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;

XOR2_X1 U738 ( .A(G107), .B(n1023), .Z(G9) );
AND3_X1 U739 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NOR2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1030) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U744 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR3_X1 U745 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1041) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1038) );
NOR3_X1 U753 ( .A1(n1050), .A2(n1057), .A3(n1044), .ZN(n1056) );
NOR2_X1 U754 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR4_X1 U755 ( .A1(n1060), .A2(n1044), .A3(n1040), .A4(n1050), .ZN(n1035) );
INV_X1 U756 ( .A(n1061), .ZN(n1050) );
NOR2_X1 U757 ( .A1(n1024), .A2(n1062), .ZN(n1060) );
NOR3_X1 U758 ( .A1(n1032), .A2(G952), .A3(n1029), .ZN(n1027) );
AND4_X1 U759 ( .A1(n1054), .A2(n1055), .A3(n1063), .A4(n1064), .ZN(n1029) );
NOR4_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(n1067) );
XOR2_X1 U762 ( .A(KEYINPUT0), .B(G472), .Z(n1070) );
XOR2_X1 U763 ( .A(n1071), .B(n1072), .Z(n1066) );
NAND2_X1 U764 ( .A1(KEYINPUT47), .A2(n1073), .ZN(n1071) );
XOR2_X1 U765 ( .A(n1074), .B(n1075), .Z(n1063) );
NOR2_X1 U766 ( .A1(KEYINPUT61), .A2(n1076), .ZN(n1075) );
INV_X1 U767 ( .A(n1077), .ZN(n1032) );
XOR2_X1 U768 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U769 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND3_X1 U770 ( .A1(G953), .A2(n1082), .A3(KEYINPUT52), .ZN(n1081) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1082) );
NAND2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U774 ( .A(n1087), .B(KEYINPUT9), .Z(n1085) );
XOR2_X1 U775 ( .A(n1088), .B(n1089), .Z(n1083) );
XOR2_X1 U776 ( .A(n1090), .B(n1091), .Z(n1089) );
XNOR2_X1 U777 ( .A(G134), .B(KEYINPUT1), .ZN(n1091) );
XOR2_X1 U778 ( .A(n1092), .B(n1093), .Z(n1088) );
XNOR2_X1 U779 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U780 ( .A1(G131), .A2(KEYINPUT17), .ZN(n1094) );
NOR2_X1 U781 ( .A1(n1096), .A2(G953), .ZN(n1078) );
XOR2_X1 U782 ( .A(n1097), .B(n1098), .Z(G69) );
NOR2_X1 U783 ( .A1(n1099), .A2(n1087), .ZN(n1098) );
AND2_X1 U784 ( .A1(G224), .A2(G898), .ZN(n1099) );
NAND2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1087), .ZN(n1101) );
XOR2_X1 U787 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
OR3_X1 U789 ( .A1(n1107), .A2(n1104), .A3(n1087), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XNOR2_X1 U791 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1108), .A2(n1114), .ZN(G63) );
NOR3_X1 U794 ( .A1(n1072), .A2(n1115), .A3(n1116), .ZN(n1114) );
NOR3_X1 U795 ( .A1(n1117), .A2(n1073), .A3(n1113), .ZN(n1116) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
AND2_X1 U797 ( .A1(n1031), .A2(G478), .ZN(n1118) );
NOR2_X1 U798 ( .A1(n1108), .A2(n1120), .ZN(G60) );
XOR2_X1 U799 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U800 ( .A1(KEYINPUT6), .A2(n1123), .ZN(n1122) );
NAND2_X1 U801 ( .A1(n1124), .A2(G475), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1105), .B(n1125), .Z(G6) );
NOR2_X1 U803 ( .A1(KEYINPUT43), .A2(n1126), .ZN(n1125) );
XOR2_X1 U804 ( .A(KEYINPUT3), .B(G104), .Z(n1126) );
NOR2_X1 U805 ( .A1(n1108), .A2(n1127), .ZN(G57) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U808 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
OR2_X1 U809 ( .A1(n1134), .A2(KEYINPUT5), .ZN(n1133) );
NAND3_X1 U810 ( .A1(n1135), .A2(n1136), .A3(KEYINPUT5), .ZN(n1132) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1128) );
AND2_X1 U812 ( .A1(G472), .A2(n1124), .ZN(n1138) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
XOR2_X1 U814 ( .A(KEYINPUT36), .B(n1141), .Z(n1139) );
NOR2_X1 U815 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1108), .A2(n1144), .ZN(G54) );
XOR2_X1 U817 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U820 ( .A(n1151), .ZN(n1150) );
NOR3_X1 U821 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1149) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
AND3_X1 U823 ( .A1(n1156), .A2(n1155), .A3(KEYINPUT19), .ZN(n1153) );
NOR2_X1 U824 ( .A1(KEYINPUT19), .A2(n1157), .ZN(n1152) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1158), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
INV_X1 U827 ( .A(n1157), .ZN(n1160) );
NAND2_X1 U828 ( .A1(n1161), .A2(n1156), .ZN(n1157) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1156), .ZN(n1159) );
NAND2_X1 U830 ( .A1(n1163), .A2(n1164), .ZN(n1156) );
NAND2_X1 U831 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U832 ( .A(n1167), .B(KEYINPUT14), .Z(n1163) );
OR2_X1 U833 ( .A1(n1166), .A2(n1165), .ZN(n1167) );
INV_X1 U834 ( .A(n1090), .ZN(n1165) );
XNOR2_X1 U835 ( .A(n1161), .B(KEYINPUT19), .ZN(n1162) );
INV_X1 U836 ( .A(n1155), .ZN(n1161) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1169), .ZN(n1155) );
XOR2_X1 U838 ( .A(n1170), .B(KEYINPUT2), .Z(n1168) );
NOR2_X1 U839 ( .A1(KEYINPUT44), .A2(n1136), .ZN(n1151) );
AND2_X1 U840 ( .A1(G469), .A2(n1124), .ZN(n1145) );
INV_X1 U841 ( .A(n1113), .ZN(n1124) );
NOR2_X1 U842 ( .A1(n1108), .A2(n1171), .ZN(G51) );
XOR2_X1 U843 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U846 ( .A1(KEYINPUT22), .A2(n1178), .ZN(n1177) );
NOR2_X1 U847 ( .A1(G125), .A2(KEYINPUT49), .ZN(n1176) );
NOR2_X1 U848 ( .A1(n1074), .A2(n1113), .ZN(n1174) );
NAND2_X1 U849 ( .A1(G902), .A2(n1031), .ZN(n1113) );
NAND3_X1 U850 ( .A1(n1096), .A2(n1179), .A3(n1180), .ZN(n1031) );
INV_X1 U851 ( .A(n1106), .ZN(n1180) );
NAND4_X1 U852 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1106) );
NOR3_X1 U853 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
INV_X1 U854 ( .A(n1188), .ZN(n1185) );
NAND2_X1 U855 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
XOR2_X1 U856 ( .A(n1191), .B(KEYINPUT20), .Z(n1189) );
NAND4_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1059), .A4(n1194), .ZN(n1181) );
NAND2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
NAND3_X1 U859 ( .A1(n1024), .A2(n1025), .A3(n1197), .ZN(n1196) );
XOR2_X1 U860 ( .A(n1198), .B(KEYINPUT59), .Z(n1197) );
NAND3_X1 U861 ( .A1(n1199), .A2(n1200), .A3(n1052), .ZN(n1195) );
XOR2_X1 U862 ( .A(KEYINPUT38), .B(n1190), .Z(n1200) );
XOR2_X1 U863 ( .A(KEYINPUT23), .B(n1105), .Z(n1179) );
NOR3_X1 U864 ( .A1(n1201), .A2(n1044), .A3(n1202), .ZN(n1105) );
AND4_X1 U865 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1096) );
AND4_X1 U866 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND3_X1 U868 ( .A1(n1213), .A2(n1046), .A3(n1214), .ZN(n1204) );
NAND2_X1 U869 ( .A1(n1215), .A2(n1216), .ZN(n1203) );
XOR2_X1 U870 ( .A(KEYINPUT63), .B(n1062), .Z(n1216) );
INV_X1 U871 ( .A(n1217), .ZN(n1215) );
XOR2_X1 U872 ( .A(n1218), .B(n1135), .Z(n1172) );
NOR2_X1 U873 ( .A1(n1087), .A2(G952), .ZN(n1108) );
XOR2_X1 U874 ( .A(G146), .B(n1212), .Z(G48) );
AND3_X1 U875 ( .A1(n1053), .A2(n1046), .A3(n1219), .ZN(n1212) );
XNOR2_X1 U876 ( .A(G143), .B(n1220), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1221), .A2(KEYINPUT62), .A3(n1214), .A4(n1046), .ZN(n1220) );
XNOR2_X1 U878 ( .A(n1213), .B(KEYINPUT40), .ZN(n1221) );
XOR2_X1 U879 ( .A(n1211), .B(n1222), .Z(G42) );
NOR2_X1 U880 ( .A1(KEYINPUT27), .A2(n1223), .ZN(n1222) );
INV_X1 U881 ( .A(G140), .ZN(n1223) );
AND3_X1 U882 ( .A1(n1061), .A2(n1224), .A3(n1219), .ZN(n1211) );
AND3_X1 U883 ( .A1(n1062), .A2(n1225), .A3(n1226), .ZN(n1219) );
XOR2_X1 U884 ( .A(n1227), .B(n1209), .Z(G39) );
NAND3_X1 U885 ( .A1(n1228), .A2(n1199), .A3(n1061), .ZN(n1209) );
XNOR2_X1 U886 ( .A(G134), .B(n1210), .ZN(G36) );
NAND3_X1 U887 ( .A1(n1214), .A2(n1024), .A3(n1061), .ZN(n1210) );
XNOR2_X1 U888 ( .A(G131), .B(n1208), .ZN(G33) );
NAND3_X1 U889 ( .A1(n1214), .A2(n1062), .A3(n1061), .ZN(n1208) );
NOR2_X1 U890 ( .A1(n1047), .A2(n1065), .ZN(n1061) );
INV_X1 U891 ( .A(n1048), .ZN(n1065) );
AND2_X1 U892 ( .A1(n1226), .A2(n1052), .ZN(n1214) );
XNOR2_X1 U893 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U894 ( .A1(n1024), .A2(n1046), .A3(n1228), .ZN(n1207) );
AND3_X1 U895 ( .A1(n1053), .A2(n1225), .A3(n1226), .ZN(n1228) );
AND3_X1 U896 ( .A1(n1229), .A2(n1059), .A3(n1192), .ZN(n1226) );
XOR2_X1 U897 ( .A(G101), .B(n1230), .Z(G3) );
AND3_X1 U898 ( .A1(n1052), .A2(n1026), .A3(n1199), .ZN(n1230) );
INV_X1 U899 ( .A(n1201), .ZN(n1026) );
XOR2_X1 U900 ( .A(G125), .B(n1231), .Z(G27) );
NOR2_X1 U901 ( .A1(n1202), .A2(n1217), .ZN(n1231) );
NAND3_X1 U902 ( .A1(n1055), .A2(n1046), .A3(n1232), .ZN(n1217) );
AND3_X1 U903 ( .A1(n1225), .A2(n1229), .A3(n1224), .ZN(n1232) );
NAND2_X1 U904 ( .A1(n1034), .A2(n1233), .ZN(n1229) );
NAND4_X1 U905 ( .A1(n1234), .A2(G953), .A3(G902), .A4(n1235), .ZN(n1233) );
XOR2_X1 U906 ( .A(n1086), .B(KEYINPUT29), .Z(n1234) );
INV_X1 U907 ( .A(G900), .ZN(n1086) );
XOR2_X1 U908 ( .A(n1182), .B(n1236), .Z(G24) );
XOR2_X1 U909 ( .A(KEYINPUT32), .B(G122), .Z(n1236) );
NAND4_X1 U910 ( .A1(n1213), .A2(n1237), .A3(n1025), .A4(n1046), .ZN(n1182) );
INV_X1 U911 ( .A(n1044), .ZN(n1025) );
NAND2_X1 U912 ( .A1(n1238), .A2(n1224), .ZN(n1044) );
XOR2_X1 U913 ( .A(KEYINPUT55), .B(n1225), .Z(n1238) );
AND2_X1 U914 ( .A1(n1239), .A2(n1068), .ZN(n1213) );
XOR2_X1 U915 ( .A(KEYINPUT54), .B(n1240), .Z(n1239) );
NAND2_X1 U916 ( .A1(n1241), .A2(n1242), .ZN(G21) );
NAND2_X1 U917 ( .A1(G119), .A2(n1188), .ZN(n1242) );
XOR2_X1 U918 ( .A(n1243), .B(KEYINPUT56), .Z(n1241) );
OR2_X1 U919 ( .A1(n1188), .A2(G119), .ZN(n1243) );
NAND4_X1 U920 ( .A1(n1046), .A2(n1225), .A3(n1199), .A4(n1244), .ZN(n1188) );
NOR2_X1 U921 ( .A1(n1245), .A2(n1224), .ZN(n1244) );
XOR2_X1 U922 ( .A(G116), .B(n1187), .Z(G18) );
AND4_X1 U923 ( .A1(n1052), .A2(n1237), .A3(n1024), .A4(n1046), .ZN(n1187) );
XOR2_X1 U924 ( .A(n1190), .B(KEYINPUT37), .Z(n1046) );
NOR2_X1 U925 ( .A1(n1068), .A2(n1240), .ZN(n1024) );
XOR2_X1 U926 ( .A(n1246), .B(KEYINPUT35), .Z(n1240) );
XOR2_X1 U927 ( .A(G113), .B(n1247), .Z(G15) );
NOR2_X1 U928 ( .A1(n1198), .A2(n1191), .ZN(n1247) );
NAND3_X1 U929 ( .A1(n1052), .A2(n1237), .A3(n1062), .ZN(n1191) );
INV_X1 U930 ( .A(n1202), .ZN(n1062) );
NAND2_X1 U931 ( .A1(n1248), .A2(n1068), .ZN(n1202) );
INV_X1 U932 ( .A(n1245), .ZN(n1237) );
NAND2_X1 U933 ( .A1(n1055), .A2(n1194), .ZN(n1245) );
INV_X1 U934 ( .A(n1040), .ZN(n1055) );
NAND2_X1 U935 ( .A1(n1058), .A2(n1059), .ZN(n1040) );
NOR2_X1 U936 ( .A1(n1224), .A2(n1225), .ZN(n1052) );
INV_X1 U937 ( .A(n1054), .ZN(n1225) );
INV_X1 U938 ( .A(n1053), .ZN(n1224) );
XOR2_X1 U939 ( .A(n1249), .B(n1250), .Z(G12) );
NAND2_X1 U940 ( .A1(KEYINPUT21), .A2(n1186), .ZN(n1250) );
NOR4_X1 U941 ( .A1(n1037), .A2(n1201), .A3(n1054), .A4(n1053), .ZN(n1186) );
XOR2_X1 U942 ( .A(n1069), .B(n1251), .Z(n1053) );
NOR2_X1 U943 ( .A1(G472), .A2(KEYINPUT34), .ZN(n1251) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1253), .ZN(n1069) );
NAND2_X1 U945 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U946 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U947 ( .A(KEYINPUT50), .B(n1258), .Z(n1254) );
NOR2_X1 U948 ( .A1(n1256), .A2(n1257), .ZN(n1258) );
NAND2_X1 U949 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U950 ( .A1(KEYINPUT45), .A2(n1261), .ZN(n1260) );
NAND2_X1 U951 ( .A1(n1140), .A2(n1262), .ZN(n1261) );
OR2_X1 U952 ( .A1(n1143), .A2(n1142), .ZN(n1262) );
NAND2_X1 U953 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND2_X1 U954 ( .A1(n1263), .A2(n1264), .ZN(n1259) );
INV_X1 U955 ( .A(KEYINPUT45), .ZN(n1264) );
XOR2_X1 U956 ( .A(n1143), .B(n1142), .Z(n1263) );
NAND3_X1 U957 ( .A1(n1265), .A2(n1087), .A3(G210), .ZN(n1143) );
XOR2_X1 U958 ( .A(n1130), .B(n1134), .Z(n1256) );
XOR2_X1 U959 ( .A(n1135), .B(n1266), .Z(n1134) );
INV_X1 U960 ( .A(n1136), .ZN(n1266) );
XOR2_X1 U961 ( .A(n1267), .B(n1268), .Z(n1130) );
XOR2_X1 U962 ( .A(KEYINPUT18), .B(G113), .Z(n1268) );
NAND2_X1 U963 ( .A1(KEYINPUT48), .A2(n1269), .ZN(n1267) );
XOR2_X1 U964 ( .A(G119), .B(G116), .Z(n1269) );
XNOR2_X1 U965 ( .A(n1270), .B(n1112), .ZN(n1054) );
NAND2_X1 U966 ( .A1(G217), .A2(n1271), .ZN(n1112) );
NAND2_X1 U967 ( .A1(n1110), .A2(n1252), .ZN(n1270) );
XNOR2_X1 U968 ( .A(n1272), .B(n1273), .ZN(n1110) );
XOR2_X1 U969 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U970 ( .A(n1276), .B(n1277), .ZN(n1275) );
AND3_X1 U971 ( .A1(G221), .A2(n1087), .A3(G234), .ZN(n1276) );
INV_X1 U972 ( .A(n1092), .ZN(n1274) );
XOR2_X1 U973 ( .A(n1227), .B(G125), .Z(n1092) );
XOR2_X1 U974 ( .A(n1278), .B(n1279), .Z(n1272) );
XOR2_X1 U975 ( .A(G128), .B(G119), .Z(n1279) );
XNOR2_X1 U976 ( .A(n1280), .B(n1281), .ZN(n1278) );
NAND2_X1 U977 ( .A1(KEYINPUT30), .A2(n1095), .ZN(n1281) );
NAND2_X1 U978 ( .A1(n1282), .A2(KEYINPUT39), .ZN(n1280) );
XOR2_X1 U979 ( .A(n1249), .B(KEYINPUT60), .Z(n1282) );
NAND4_X1 U980 ( .A1(n1190), .A2(n1192), .A3(n1059), .A4(n1194), .ZN(n1201) );
NAND2_X1 U981 ( .A1(n1034), .A2(n1283), .ZN(n1194) );
NAND4_X1 U982 ( .A1(G953), .A2(G902), .A3(n1235), .A4(n1107), .ZN(n1283) );
INV_X1 U983 ( .A(G898), .ZN(n1107) );
NAND3_X1 U984 ( .A1(n1077), .A2(n1235), .A3(G952), .ZN(n1034) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1235) );
XOR2_X1 U986 ( .A(n1087), .B(KEYINPUT24), .Z(n1077) );
NAND2_X1 U987 ( .A1(G221), .A2(n1271), .ZN(n1059) );
NAND2_X1 U988 ( .A1(G234), .A2(n1284), .ZN(n1271) );
XOR2_X1 U989 ( .A(KEYINPUT4), .B(n1285), .Z(n1284) );
INV_X1 U990 ( .A(n1058), .ZN(n1192) );
XOR2_X1 U991 ( .A(n1286), .B(G469), .Z(n1058) );
NAND2_X1 U992 ( .A1(n1287), .A2(n1252), .ZN(n1286) );
XOR2_X1 U993 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U994 ( .A(n1166), .B(n1136), .Z(n1289) );
XNOR2_X1 U995 ( .A(G131), .B(n1290), .ZN(n1136) );
NOR2_X1 U996 ( .A1(KEYINPUT8), .A2(n1291), .ZN(n1290) );
XOR2_X1 U997 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U998 ( .A(G134), .B(KEYINPUT12), .ZN(n1293) );
NAND2_X1 U999 ( .A1(KEYINPUT46), .A2(n1227), .ZN(n1292) );
INV_X1 U1000 ( .A(G137), .ZN(n1227) );
XOR2_X1 U1001 ( .A(n1294), .B(n1142), .Z(n1166) );
XOR2_X1 U1002 ( .A(n1295), .B(G107), .Z(n1294) );
INV_X1 U1003 ( .A(G104), .ZN(n1295) );
XOR2_X1 U1004 ( .A(n1296), .B(n1297), .Z(n1288) );
NOR2_X1 U1005 ( .A1(KEYINPUT33), .A2(n1090), .ZN(n1297) );
NAND2_X1 U1006 ( .A1(n1298), .A2(n1299), .ZN(n1090) );
OR2_X1 U1007 ( .A1(n1300), .A2(G128), .ZN(n1299) );
XOR2_X1 U1008 ( .A(n1301), .B(KEYINPUT57), .Z(n1298) );
NAND2_X1 U1009 ( .A1(G128), .A2(n1300), .ZN(n1301) );
NAND2_X1 U1010 ( .A1(n1169), .A2(n1170), .ZN(n1296) );
NAND3_X1 U1011 ( .A1(n1302), .A2(n1087), .A3(G227), .ZN(n1170) );
INV_X1 U1012 ( .A(n1303), .ZN(n1302) );
NAND2_X1 U1013 ( .A1(n1303), .A2(n1304), .ZN(n1169) );
NAND2_X1 U1014 ( .A1(G227), .A2(n1087), .ZN(n1304) );
XOR2_X1 U1015 ( .A(n1249), .B(n1095), .Z(n1303) );
INV_X1 U1016 ( .A(n1198), .ZN(n1190) );
NAND2_X1 U1017 ( .A1(n1047), .A2(n1048), .ZN(n1198) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1305), .ZN(n1048) );
XNOR2_X1 U1019 ( .A(n1306), .B(n1074), .ZN(n1047) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1305), .ZN(n1074) );
NAND2_X1 U1021 ( .A1(n1285), .A2(n1265), .ZN(n1305) );
XOR2_X1 U1022 ( .A(G902), .B(KEYINPUT28), .Z(n1285) );
NAND2_X1 U1023 ( .A1(KEYINPUT41), .A2(n1076), .ZN(n1306) );
NAND2_X1 U1024 ( .A1(n1307), .A2(n1252), .ZN(n1076) );
INV_X1 U1025 ( .A(G902), .ZN(n1252) );
XOR2_X1 U1026 ( .A(n1218), .B(n1308), .Z(n1307) );
NOR2_X1 U1027 ( .A1(KEYINPUT11), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1028 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1029 ( .A(n1312), .B(n1135), .ZN(n1311) );
XNOR2_X1 U1030 ( .A(n1313), .B(n1314), .ZN(n1135) );
XOR2_X1 U1031 ( .A(n1315), .B(G128), .Z(n1313) );
NAND2_X1 U1032 ( .A1(KEYINPUT7), .A2(n1277), .ZN(n1315) );
NAND2_X1 U1033 ( .A1(KEYINPUT10), .A2(n1316), .ZN(n1312) );
INV_X1 U1034 ( .A(n1178), .ZN(n1316) );
NAND2_X1 U1035 ( .A1(G224), .A2(n1087), .ZN(n1178) );
XOR2_X1 U1036 ( .A(KEYINPUT25), .B(G125), .Z(n1310) );
XNOR2_X1 U1037 ( .A(n1104), .B(KEYINPUT16), .ZN(n1218) );
XNOR2_X1 U1038 ( .A(n1317), .B(n1318), .ZN(n1104) );
XOR2_X1 U1039 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1040 ( .A(G110), .B(G104), .Z(n1320) );
XOR2_X1 U1041 ( .A(G119), .B(G113), .Z(n1319) );
XOR2_X1 U1042 ( .A(n1321), .B(n1322), .Z(n1317) );
XNOR2_X1 U1043 ( .A(n1323), .B(n1142), .ZN(n1321) );
XNOR2_X1 U1044 ( .A(G101), .B(KEYINPUT42), .ZN(n1142) );
NAND2_X1 U1045 ( .A1(KEYINPUT15), .A2(G107), .ZN(n1323) );
INV_X1 U1046 ( .A(n1199), .ZN(n1037) );
NOR2_X1 U1047 ( .A1(n1068), .A2(n1246), .ZN(n1199) );
INV_X1 U1048 ( .A(n1248), .ZN(n1246) );
XOR2_X1 U1049 ( .A(n1072), .B(n1073), .Z(n1248) );
INV_X1 U1050 ( .A(G478), .ZN(n1073) );
NOR2_X1 U1051 ( .A1(n1119), .A2(G902), .ZN(n1072) );
INV_X1 U1052 ( .A(n1117), .ZN(n1119) );
NAND2_X1 U1053 ( .A1(n1324), .A2(n1325), .ZN(n1117) );
NAND2_X1 U1054 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND3_X1 U1055 ( .A1(G217), .A2(n1087), .A3(G234), .ZN(n1327) );
INV_X1 U1056 ( .A(n1328), .ZN(n1326) );
NAND4_X1 U1057 ( .A1(G217), .A2(n1087), .A3(G234), .A4(n1328), .ZN(n1324) );
XOR2_X1 U1058 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1059 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1060 ( .A(G134), .B(G128), .Z(n1332) );
XOR2_X1 U1061 ( .A(KEYINPUT58), .B(KEYINPUT13), .Z(n1331) );
XOR2_X1 U1062 ( .A(n1333), .B(n1322), .Z(n1329) );
XOR2_X1 U1063 ( .A(G116), .B(G122), .Z(n1322) );
XNOR2_X1 U1064 ( .A(G107), .B(n1314), .ZN(n1333) );
XNOR2_X1 U1065 ( .A(n1334), .B(G475), .ZN(n1068) );
OR2_X1 U1066 ( .A1(n1123), .A2(G902), .ZN(n1334) );
XNOR2_X1 U1067 ( .A(n1335), .B(n1336), .ZN(n1123) );
XOR2_X1 U1068 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1069 ( .A(G113), .B(G104), .Z(n1338) );
XOR2_X1 U1070 ( .A(G131), .B(G122), .Z(n1337) );
XNOR2_X1 U1071 ( .A(n1339), .B(n1300), .ZN(n1335) );
XOR2_X1 U1072 ( .A(n1277), .B(n1314), .Z(n1300) );
XOR2_X1 U1073 ( .A(G143), .B(KEYINPUT26), .Z(n1314) );
XNOR2_X1 U1074 ( .A(G146), .B(KEYINPUT51), .ZN(n1277) );
XOR2_X1 U1075 ( .A(n1340), .B(n1341), .Z(n1339) );
AND3_X1 U1076 ( .A1(G214), .A2(n1087), .A3(n1265), .ZN(n1341) );
INV_X1 U1077 ( .A(G237), .ZN(n1265) );
INV_X1 U1078 ( .A(G953), .ZN(n1087) );
NAND2_X1 U1079 ( .A1(KEYINPUT53), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1080 ( .A(G125), .B(n1095), .ZN(n1342) );
XNOR2_X1 U1081 ( .A(G140), .B(KEYINPUT31), .ZN(n1095) );
INV_X1 U1082 ( .A(G110), .ZN(n1249) );
endmodule


