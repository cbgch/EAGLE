//Key = 0111101101010111111111100010100111001100010011000001101011010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374;

XNOR2_X1 U751 ( .A(n1033), .B(n1034), .ZN(G9) );
NAND2_X1 U752 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND3_X1 U753 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
INV_X1 U754 ( .A(KEYINPUT52), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1040), .A2(KEYINPUT52), .ZN(n1035) );
NOR2_X1 U756 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR3_X1 U757 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NAND3_X1 U758 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1043) );
NAND2_X1 U759 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND4_X1 U761 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NAND2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
OR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U768 ( .A1(n1063), .A2(n1069), .A3(n1059), .ZN(n1051) );
NAND2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U770 ( .A1(n1072), .A2(n1073), .A3(n1054), .ZN(n1071) );
OR2_X1 U771 ( .A1(n1056), .A2(n1053), .ZN(n1073) );
NAND3_X1 U772 ( .A1(n1074), .A2(n1038), .A3(n1056), .ZN(n1072) );
INV_X1 U773 ( .A(n1075), .ZN(n1038) );
NAND2_X1 U774 ( .A1(n1053), .A2(n1076), .ZN(n1070) );
INV_X1 U775 ( .A(n1077), .ZN(n1049) );
NOR3_X1 U776 ( .A1(n1078), .A2(G953), .A3(G952), .ZN(n1041) );
INV_X1 U777 ( .A(n1046), .ZN(n1078) );
NAND4_X1 U778 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1046) );
NOR4_X1 U779 ( .A1(n1068), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1082) );
INV_X1 U780 ( .A(n1063), .ZN(n1085) );
INV_X1 U781 ( .A(n1086), .ZN(n1068) );
NOR3_X1 U782 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1081) );
NOR2_X1 U783 ( .A1(KEYINPUT26), .A2(n1090), .ZN(n1089) );
INV_X1 U784 ( .A(n1091), .ZN(n1090) );
AND2_X1 U785 ( .A1(n1092), .A2(KEYINPUT26), .ZN(n1088) );
XOR2_X1 U786 ( .A(KEYINPUT1), .B(n1093), .Z(n1087) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U789 ( .A(KEYINPUT41), .B(n1098), .ZN(n1097) );
XOR2_X1 U790 ( .A(n1099), .B(KEYINPUT34), .Z(n1079) );
NAND2_X1 U791 ( .A1(G469), .A2(n1100), .ZN(n1099) );
XOR2_X1 U792 ( .A(n1101), .B(n1102), .Z(G72) );
XOR2_X1 U793 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U795 ( .A1(G900), .A2(n1107), .ZN(n1106) );
XOR2_X1 U796 ( .A(KEYINPUT10), .B(G227), .Z(n1107) );
INV_X1 U797 ( .A(n1108), .ZN(n1105) );
NAND3_X1 U798 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1103) );
XOR2_X1 U799 ( .A(n1112), .B(KEYINPUT29), .Z(n1111) );
NAND2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
OR2_X1 U802 ( .A1(n1114), .A2(n1113), .ZN(n1109) );
XNOR2_X1 U803 ( .A(n1117), .B(n1118), .ZN(n1114) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1117) );
XNOR2_X1 U806 ( .A(G137), .B(n1123), .ZN(n1122) );
NAND2_X1 U807 ( .A1(KEYINPUT31), .A2(G134), .ZN(n1123) );
NAND2_X1 U808 ( .A1(KEYINPUT9), .A2(n1124), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1125), .A2(G953), .ZN(n1101) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U811 ( .A1(n1128), .A2(n1108), .ZN(n1127) );
XOR2_X1 U812 ( .A(G953), .B(KEYINPUT19), .Z(n1108) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U814 ( .A1(n1131), .A2(n1132), .A3(KEYINPUT14), .ZN(n1126) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XNOR2_X1 U816 ( .A(KEYINPUT38), .B(n1135), .ZN(n1134) );
XOR2_X1 U817 ( .A(KEYINPUT33), .B(n1136), .Z(n1133) );
NAND2_X1 U818 ( .A1(n1136), .A2(n1135), .ZN(n1131) );
NAND2_X1 U819 ( .A1(n1047), .A2(n1045), .ZN(n1135) );
AND2_X1 U820 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U821 ( .A1(n1116), .A2(n1130), .ZN(n1138) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U823 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR3_X1 U824 ( .A1(n1143), .A2(KEYINPUT48), .A3(n1144), .ZN(n1141) );
NOR2_X1 U825 ( .A1(n1145), .A2(n1146), .ZN(G63) );
XOR2_X1 U826 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1143), .ZN(n1147) );
NOR2_X1 U828 ( .A1(G952), .A2(n1150), .ZN(n1145) );
XNOR2_X1 U829 ( .A(KEYINPUT6), .B(n1047), .ZN(n1150) );
NOR2_X1 U830 ( .A1(n1139), .A2(n1151), .ZN(G60) );
XNOR2_X1 U831 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1143), .ZN(n1152) );
XNOR2_X1 U833 ( .A(n1155), .B(n1156), .ZN(G6) );
NOR3_X1 U834 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(G57) );
AND2_X1 U835 ( .A1(KEYINPUT57), .A2(n1139), .ZN(n1159) );
NOR3_X1 U836 ( .A1(KEYINPUT57), .A2(G953), .A3(G952), .ZN(n1158) );
XOR2_X1 U837 ( .A(n1160), .B(n1161), .Z(n1157) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U839 ( .A1(n1164), .A2(n1143), .ZN(n1163) );
NAND3_X1 U840 ( .A1(n1165), .A2(n1166), .A3(KEYINPUT11), .ZN(n1162) );
NAND2_X1 U841 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
INV_X1 U842 ( .A(n1169), .ZN(n1168) );
NAND2_X1 U843 ( .A1(KEYINPUT17), .A2(n1170), .ZN(n1167) );
OR2_X1 U844 ( .A1(n1171), .A2(KEYINPUT23), .ZN(n1170) );
NAND2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
NAND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U847 ( .A1(n1169), .A2(KEYINPUT17), .ZN(n1174) );
NOR2_X1 U848 ( .A1(n1175), .A2(n1176), .ZN(n1169) );
INV_X1 U849 ( .A(KEYINPUT23), .ZN(n1173) );
XNOR2_X1 U850 ( .A(G101), .B(n1177), .ZN(n1160) );
AND3_X1 U851 ( .A1(G210), .A2(n1178), .A3(n1179), .ZN(n1177) );
INV_X1 U852 ( .A(KEYINPUT30), .ZN(n1178) );
NOR2_X1 U853 ( .A1(n1139), .A2(n1180), .ZN(G54) );
XOR2_X1 U854 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U856 ( .A1(KEYINPUT3), .A2(n1185), .ZN(n1183) );
XOR2_X1 U857 ( .A(n1186), .B(n1187), .Z(n1181) );
XNOR2_X1 U858 ( .A(G140), .B(n1188), .ZN(n1187) );
NAND3_X1 U859 ( .A1(n1189), .A2(n1190), .A3(G469), .ZN(n1186) );
NAND2_X1 U860 ( .A1(n1143), .A2(n1191), .ZN(n1190) );
INV_X1 U861 ( .A(KEYINPUT27), .ZN(n1191) );
NAND2_X1 U862 ( .A1(KEYINPUT27), .A2(n1192), .ZN(n1189) );
OR2_X1 U863 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR3_X1 U864 ( .A1(n1139), .A2(n1195), .A3(n1196), .ZN(G51) );
NOR2_X1 U865 ( .A1(n1137), .A2(n1197), .ZN(n1196) );
XOR2_X1 U866 ( .A(KEYINPUT49), .B(n1198), .Z(n1197) );
NOR2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1195) );
XNOR2_X1 U868 ( .A(n1198), .B(KEYINPUT12), .ZN(n1200) );
XNOR2_X1 U869 ( .A(n1201), .B(n1202), .ZN(n1198) );
NOR3_X1 U870 ( .A1(n1143), .A2(KEYINPUT5), .A3(n1098), .ZN(n1202) );
NAND2_X1 U871 ( .A1(G902), .A2(n1193), .ZN(n1143) );
NAND2_X1 U872 ( .A1(n1203), .A2(n1125), .ZN(n1193) );
INV_X1 U873 ( .A(n1044), .ZN(n1125) );
NAND2_X1 U874 ( .A1(n1204), .A2(n1205), .ZN(n1044) );
AND4_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
NOR4_X1 U876 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1204) );
NOR2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U878 ( .A(n1076), .B(KEYINPUT53), .ZN(n1214) );
NOR3_X1 U879 ( .A1(n1216), .A2(n1065), .A3(n1217), .ZN(n1212) );
XOR2_X1 U880 ( .A(n1045), .B(KEYINPUT59), .Z(n1203) );
NAND2_X1 U881 ( .A1(n1218), .A2(n1219), .ZN(n1045) );
NOR4_X1 U882 ( .A1(n1220), .A2(n1156), .A3(n1040), .A4(n1221), .ZN(n1219) );
INV_X1 U883 ( .A(n1222), .ZN(n1221) );
AND2_X1 U884 ( .A1(n1075), .A2(n1037), .ZN(n1040) );
AND2_X1 U885 ( .A1(n1223), .A2(n1037), .ZN(n1156) );
AND2_X1 U886 ( .A1(n1063), .A2(n1224), .ZN(n1037) );
AND4_X1 U887 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1218) );
NAND3_X1 U888 ( .A1(n1229), .A2(n1063), .A3(n1230), .ZN(n1228) );
NAND2_X1 U889 ( .A1(n1231), .A2(n1232), .ZN(n1201) );
NAND2_X1 U890 ( .A1(G125), .A2(n1233), .ZN(n1232) );
NAND2_X1 U891 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U892 ( .A1(n1236), .A2(n1237), .ZN(n1231) );
XOR2_X1 U893 ( .A(n1238), .B(n1239), .Z(n1236) );
NOR2_X1 U894 ( .A1(n1047), .A2(G952), .ZN(n1139) );
XOR2_X1 U895 ( .A(n1240), .B(n1241), .Z(G48) );
NAND2_X1 U896 ( .A1(KEYINPUT62), .A2(G146), .ZN(n1241) );
NAND2_X1 U897 ( .A1(n1242), .A2(n1076), .ZN(n1240) );
INV_X1 U898 ( .A(n1215), .ZN(n1242) );
NAND4_X1 U899 ( .A1(n1223), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1215) );
XNOR2_X1 U900 ( .A(G143), .B(n1246), .ZN(G45) );
NAND3_X1 U901 ( .A1(n1247), .A2(n1229), .A3(n1248), .ZN(n1246) );
XNOR2_X1 U902 ( .A(n1243), .B(KEYINPUT22), .ZN(n1248) );
XNOR2_X1 U903 ( .A(n1211), .B(n1249), .ZN(G42) );
NAND2_X1 U904 ( .A1(KEYINPUT4), .A2(G140), .ZN(n1249) );
AND4_X1 U905 ( .A1(n1059), .A2(n1223), .A3(n1250), .A4(n1062), .ZN(n1211) );
AND2_X1 U906 ( .A1(n1245), .A2(n1076), .ZN(n1250) );
XOR2_X1 U907 ( .A(G137), .B(n1210), .Z(G39) );
AND3_X1 U908 ( .A1(n1251), .A2(n1053), .A3(n1059), .ZN(n1210) );
XNOR2_X1 U909 ( .A(G134), .B(n1209), .ZN(G36) );
NAND3_X1 U910 ( .A1(n1247), .A2(n1075), .A3(n1059), .ZN(n1209) );
XNOR2_X1 U911 ( .A(G131), .B(n1208), .ZN(G33) );
NAND3_X1 U912 ( .A1(n1247), .A2(n1223), .A3(n1059), .ZN(n1208) );
AND2_X1 U913 ( .A1(n1067), .A2(n1086), .ZN(n1059) );
INV_X1 U914 ( .A(n1216), .ZN(n1247) );
NAND3_X1 U915 ( .A1(n1061), .A2(n1245), .A3(n1076), .ZN(n1216) );
XNOR2_X1 U916 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U917 ( .A1(n1075), .A2(n1243), .A3(n1251), .ZN(n1207) );
AND3_X1 U918 ( .A1(n1244), .A2(n1245), .A3(n1076), .ZN(n1251) );
XNOR2_X1 U919 ( .A(G101), .B(n1227), .ZN(G3) );
NAND3_X1 U920 ( .A1(n1224), .A2(n1061), .A3(n1053), .ZN(n1227) );
XNOR2_X1 U921 ( .A(G125), .B(n1206), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1223), .A2(n1062), .A3(n1252), .A4(n1245), .ZN(n1206) );
NAND2_X1 U923 ( .A1(n1077), .A2(n1253), .ZN(n1245) );
NAND2_X1 U924 ( .A1(n1115), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U925 ( .A(G900), .B(KEYINPUT24), .ZN(n1115) );
XNOR2_X1 U926 ( .A(G122), .B(n1255), .ZN(G24) );
NAND4_X1 U927 ( .A1(n1256), .A2(n1229), .A3(n1252), .A4(n1063), .ZN(n1255) );
INV_X1 U928 ( .A(n1217), .ZN(n1229) );
NAND2_X1 U929 ( .A1(n1257), .A2(n1092), .ZN(n1217) );
XOR2_X1 U930 ( .A(n1258), .B(KEYINPUT40), .Z(n1256) );
XOR2_X1 U931 ( .A(n1220), .B(n1259), .Z(G21) );
NOR2_X1 U932 ( .A1(KEYINPUT58), .A2(n1260), .ZN(n1259) );
AND3_X1 U933 ( .A1(n1230), .A2(n1244), .A3(n1053), .ZN(n1220) );
NAND2_X1 U934 ( .A1(n1261), .A2(n1262), .ZN(n1244) );
NAND3_X1 U935 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
INV_X1 U936 ( .A(KEYINPUT42), .ZN(n1265) );
NAND2_X1 U937 ( .A1(KEYINPUT42), .A2(n1062), .ZN(n1261) );
XNOR2_X1 U938 ( .A(G116), .B(n1226), .ZN(G18) );
NAND3_X1 U939 ( .A1(n1075), .A2(n1061), .A3(n1230), .ZN(n1226) );
NOR2_X1 U940 ( .A1(n1092), .A2(n1080), .ZN(n1075) );
XOR2_X1 U941 ( .A(n1225), .B(n1266), .Z(G15) );
NAND2_X1 U942 ( .A1(n1267), .A2(G113), .ZN(n1266) );
XNOR2_X1 U943 ( .A(KEYINPUT56), .B(KEYINPUT16), .ZN(n1267) );
NAND3_X1 U944 ( .A1(n1230), .A2(n1061), .A3(n1223), .ZN(n1225) );
INV_X1 U945 ( .A(n1074), .ZN(n1223) );
NAND2_X1 U946 ( .A1(n1080), .A2(n1092), .ZN(n1074) );
INV_X1 U947 ( .A(n1257), .ZN(n1080) );
NAND2_X1 U948 ( .A1(n1268), .A2(n1269), .ZN(n1061) );
OR3_X1 U949 ( .A1(n1270), .A2(n1263), .A3(KEYINPUT42), .ZN(n1269) );
NAND2_X1 U950 ( .A1(KEYINPUT42), .A2(n1063), .ZN(n1268) );
NOR2_X1 U951 ( .A1(n1264), .A2(n1263), .ZN(n1063) );
AND2_X1 U952 ( .A1(n1252), .A2(n1258), .ZN(n1230) );
NOR3_X1 U953 ( .A1(n1065), .A2(n1083), .A3(n1271), .ZN(n1252) );
INV_X1 U954 ( .A(n1243), .ZN(n1065) );
XNOR2_X1 U955 ( .A(G110), .B(n1222), .ZN(G12) );
NAND3_X1 U956 ( .A1(n1062), .A2(n1224), .A3(n1053), .ZN(n1222) );
NOR2_X1 U957 ( .A1(n1257), .A2(n1092), .ZN(n1053) );
NAND2_X1 U958 ( .A1(n1091), .A2(n1272), .ZN(n1092) );
NAND3_X1 U959 ( .A1(n1154), .A2(n1194), .A3(n1153), .ZN(n1272) );
INV_X1 U960 ( .A(G475), .ZN(n1154) );
NAND2_X1 U961 ( .A1(G475), .A2(n1273), .ZN(n1091) );
NAND2_X1 U962 ( .A1(n1153), .A2(n1194), .ZN(n1273) );
XOR2_X1 U963 ( .A(n1274), .B(n1275), .Z(n1153) );
XNOR2_X1 U964 ( .A(n1276), .B(n1277), .ZN(n1275) );
NOR2_X1 U965 ( .A1(KEYINPUT47), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U966 ( .A(n1155), .B(n1279), .ZN(n1278) );
INV_X1 U967 ( .A(G104), .ZN(n1155) );
XNOR2_X1 U968 ( .A(n1280), .B(n1281), .ZN(n1274) );
NOR2_X1 U969 ( .A1(KEYINPUT60), .A2(n1282), .ZN(n1281) );
XOR2_X1 U970 ( .A(n1124), .B(n1283), .Z(n1282) );
XOR2_X1 U971 ( .A(n1284), .B(G143), .Z(n1283) );
NAND2_X1 U972 ( .A1(G214), .A2(n1179), .ZN(n1284) );
XOR2_X1 U973 ( .A(n1285), .B(n1149), .Z(n1257) );
INV_X1 U974 ( .A(G478), .ZN(n1149) );
OR2_X1 U975 ( .A1(n1148), .A2(G902), .ZN(n1285) );
XNOR2_X1 U976 ( .A(n1286), .B(n1287), .ZN(n1148) );
XOR2_X1 U977 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U978 ( .A(n1290), .B(G122), .ZN(n1289) );
XOR2_X1 U979 ( .A(G143), .B(G134), .Z(n1288) );
XOR2_X1 U980 ( .A(n1291), .B(n1292), .Z(n1286) );
AND2_X1 U981 ( .A1(n1293), .A2(G217), .ZN(n1292) );
XNOR2_X1 U982 ( .A(n1294), .B(n1034), .ZN(n1291) );
NAND2_X1 U983 ( .A1(KEYINPUT13), .A2(n1295), .ZN(n1294) );
INV_X1 U984 ( .A(G116), .ZN(n1295) );
AND3_X1 U985 ( .A1(n1076), .A2(n1258), .A3(n1243), .ZN(n1224) );
NOR2_X1 U986 ( .A1(n1296), .A2(n1067), .ZN(n1243) );
NOR2_X1 U987 ( .A1(n1297), .A2(n1094), .ZN(n1067) );
AND2_X1 U988 ( .A1(n1096), .A2(n1098), .ZN(n1094) );
NOR2_X1 U989 ( .A1(n1098), .A2(n1096), .ZN(n1297) );
AND2_X1 U990 ( .A1(n1298), .A2(n1194), .ZN(n1096) );
XNOR2_X1 U991 ( .A(n1299), .B(n1137), .ZN(n1298) );
INV_X1 U992 ( .A(n1199), .ZN(n1137) );
XNOR2_X1 U993 ( .A(n1300), .B(n1301), .ZN(n1199) );
XNOR2_X1 U994 ( .A(n1302), .B(n1279), .ZN(n1301) );
XOR2_X1 U995 ( .A(G113), .B(G122), .Z(n1279) );
NAND2_X1 U996 ( .A1(KEYINPUT63), .A2(n1303), .ZN(n1302) );
XOR2_X1 U997 ( .A(n1304), .B(n1305), .Z(n1300) );
NOR2_X1 U998 ( .A1(KEYINPUT0), .A2(n1306), .ZN(n1305) );
XOR2_X1 U999 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1000 ( .A(G104), .B(KEYINPUT25), .ZN(n1308) );
NAND2_X1 U1001 ( .A1(KEYINPUT44), .A2(n1034), .ZN(n1307) );
INV_X1 U1002 ( .A(G107), .ZN(n1034) );
XNOR2_X1 U1003 ( .A(G101), .B(G110), .ZN(n1304) );
NAND2_X1 U1004 ( .A1(n1309), .A2(n1310), .ZN(n1299) );
NAND3_X1 U1005 ( .A1(n1311), .A2(n1312), .A3(G125), .ZN(n1310) );
NAND3_X1 U1006 ( .A1(n1313), .A2(n1314), .A3(n1234), .ZN(n1311) );
NAND2_X1 U1007 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1008 ( .A1(KEYINPUT50), .A2(n1239), .ZN(n1313) );
NAND4_X1 U1009 ( .A1(n1317), .A2(n1235), .A3(n1318), .A4(n1319), .ZN(n1309) );
OR2_X1 U1010 ( .A1(n1316), .A2(n1239), .ZN(n1319) );
INV_X1 U1011 ( .A(KEYINPUT50), .ZN(n1316) );
OR2_X1 U1012 ( .A1(n1234), .A2(KEYINPUT50), .ZN(n1318) );
NAND2_X1 U1013 ( .A1(n1239), .A2(n1238), .ZN(n1234) );
INV_X1 U1014 ( .A(n1315), .ZN(n1235) );
NOR2_X1 U1015 ( .A1(n1238), .A2(n1239), .ZN(n1315) );
NOR2_X1 U1016 ( .A1(n1129), .A2(G953), .ZN(n1239) );
INV_X1 U1017 ( .A(G224), .ZN(n1129) );
NAND2_X1 U1018 ( .A1(G125), .A2(n1312), .ZN(n1317) );
INV_X1 U1019 ( .A(KEYINPUT61), .ZN(n1312) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1320), .ZN(n1098) );
XNOR2_X1 U1021 ( .A(n1086), .B(KEYINPUT35), .ZN(n1296) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1320), .ZN(n1086) );
NAND2_X1 U1023 ( .A1(n1321), .A2(n1194), .ZN(n1320) );
INV_X1 U1024 ( .A(G237), .ZN(n1321) );
NAND2_X1 U1025 ( .A1(n1322), .A2(n1077), .ZN(n1258) );
NAND3_X1 U1026 ( .A1(n1323), .A2(n1047), .A3(G952), .ZN(n1077) );
NAND2_X1 U1027 ( .A1(n1254), .A2(n1130), .ZN(n1322) );
INV_X1 U1028 ( .A(G898), .ZN(n1130) );
AND3_X1 U1029 ( .A1(n1116), .A2(n1323), .A3(G902), .ZN(n1254) );
NAND2_X1 U1030 ( .A1(G237), .A2(G234), .ZN(n1323) );
XNOR2_X1 U1031 ( .A(G953), .B(KEYINPUT7), .ZN(n1116) );
NOR2_X1 U1032 ( .A1(n1083), .A2(n1054), .ZN(n1076) );
INV_X1 U1033 ( .A(n1271), .ZN(n1054) );
NAND2_X1 U1034 ( .A1(n1324), .A2(n1325), .ZN(n1271) );
NAND2_X1 U1035 ( .A1(G469), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1036 ( .A1(KEYINPUT54), .A2(n1327), .ZN(n1326) );
INV_X1 U1037 ( .A(n1100), .ZN(n1327) );
NAND2_X1 U1038 ( .A1(n1084), .A2(KEYINPUT54), .ZN(n1324) );
NOR2_X1 U1039 ( .A1(n1100), .A2(G469), .ZN(n1084) );
NAND2_X1 U1040 ( .A1(n1328), .A2(n1194), .ZN(n1100) );
XOR2_X1 U1041 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1042 ( .A(KEYINPUT21), .B(n1188), .Z(n1330) );
AND2_X1 U1043 ( .A1(G227), .A2(n1047), .ZN(n1188) );
XOR2_X1 U1044 ( .A(n1331), .B(n1332), .Z(n1329) );
NOR2_X1 U1045 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NOR2_X1 U1046 ( .A1(G110), .A2(n1335), .ZN(n1334) );
XNOR2_X1 U1047 ( .A(KEYINPUT45), .B(n1336), .ZN(n1335) );
INV_X1 U1048 ( .A(G140), .ZN(n1336) );
NOR2_X1 U1049 ( .A1(G140), .A2(n1185), .ZN(n1333) );
NAND2_X1 U1050 ( .A1(KEYINPUT20), .A2(n1184), .ZN(n1331) );
XOR2_X1 U1051 ( .A(n1337), .B(n1338), .Z(n1184) );
XOR2_X1 U1052 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1053 ( .A(KEYINPUT18), .B(G101), .Z(n1340) );
NOR2_X1 U1054 ( .A1(KEYINPUT55), .A2(n1341), .ZN(n1339) );
XNOR2_X1 U1055 ( .A(G104), .B(G107), .ZN(n1341) );
XOR2_X1 U1056 ( .A(n1342), .B(n1120), .Z(n1337) );
XOR2_X1 U1057 ( .A(G143), .B(KEYINPUT46), .Z(n1120) );
XNOR2_X1 U1058 ( .A(n1343), .B(n1344), .ZN(n1342) );
INV_X1 U1059 ( .A(n1056), .ZN(n1083) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1345), .ZN(n1056) );
AND2_X1 U1061 ( .A1(n1270), .A2(n1263), .ZN(n1062) );
XOR2_X1 U1062 ( .A(n1346), .B(n1144), .Z(n1263) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1345), .ZN(n1144) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1194), .ZN(n1345) );
OR2_X1 U1065 ( .A1(n1142), .A2(G902), .ZN(n1346) );
XNOR2_X1 U1066 ( .A(n1347), .B(n1348), .ZN(n1142) );
XNOR2_X1 U1067 ( .A(n1349), .B(n1113), .ZN(n1348) );
INV_X1 U1068 ( .A(n1280), .ZN(n1113) );
XNOR2_X1 U1069 ( .A(G140), .B(n1237), .ZN(n1280) );
INV_X1 U1070 ( .A(G125), .ZN(n1237) );
XNOR2_X1 U1071 ( .A(n1350), .B(n1351), .ZN(n1347) );
INV_X1 U1072 ( .A(n1343), .ZN(n1351) );
XOR2_X1 U1073 ( .A(G137), .B(n1119), .Z(n1343) );
XNOR2_X1 U1074 ( .A(n1290), .B(G146), .ZN(n1119) );
XNOR2_X1 U1075 ( .A(n1352), .B(n1185), .ZN(n1350) );
INV_X1 U1076 ( .A(G110), .ZN(n1185) );
NAND2_X1 U1077 ( .A1(G221), .A2(n1293), .ZN(n1352) );
AND2_X1 U1078 ( .A1(G234), .A2(n1047), .ZN(n1293) );
INV_X1 U1079 ( .A(G953), .ZN(n1047) );
INV_X1 U1080 ( .A(n1264), .ZN(n1270) );
XOR2_X1 U1081 ( .A(n1353), .B(n1164), .Z(n1264) );
INV_X1 U1082 ( .A(G472), .ZN(n1164) );
NAND2_X1 U1083 ( .A1(n1354), .A2(n1194), .ZN(n1353) );
INV_X1 U1084 ( .A(G902), .ZN(n1194) );
XOR2_X1 U1085 ( .A(n1355), .B(n1356), .Z(n1354) );
XNOR2_X1 U1086 ( .A(n1171), .B(n1357), .ZN(n1356) );
NOR3_X1 U1087 ( .A1(n1175), .A2(n1358), .A3(n1359), .ZN(n1357) );
AND2_X1 U1088 ( .A1(KEYINPUT28), .A2(n1176), .ZN(n1359) );
AND2_X1 U1089 ( .A1(n1360), .A2(n1238), .ZN(n1176) );
NOR2_X1 U1090 ( .A1(KEYINPUT28), .A2(n1238), .ZN(n1358) );
NOR2_X1 U1091 ( .A1(n1238), .A2(n1360), .ZN(n1175) );
XNOR2_X1 U1092 ( .A(n1344), .B(G137), .ZN(n1360) );
XNOR2_X1 U1093 ( .A(G134), .B(n1124), .ZN(n1344) );
XNOR2_X1 U1094 ( .A(G131), .B(KEYINPUT36), .ZN(n1124) );
NAND2_X1 U1095 ( .A1(n1361), .A2(n1362), .ZN(n1238) );
NAND2_X1 U1096 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1097 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1098 ( .A1(KEYINPUT15), .A2(n1290), .ZN(n1366) );
INV_X1 U1099 ( .A(G128), .ZN(n1290) );
INV_X1 U1100 ( .A(KEYINPUT39), .ZN(n1365) );
NAND2_X1 U1101 ( .A1(G128), .A2(n1367), .ZN(n1361) );
NAND2_X1 U1102 ( .A1(KEYINPUT15), .A2(n1368), .ZN(n1367) );
OR2_X1 U1103 ( .A1(n1363), .A2(KEYINPUT39), .ZN(n1368) );
XNOR2_X1 U1104 ( .A(n1369), .B(n1370), .ZN(n1363) );
XOR2_X1 U1105 ( .A(KEYINPUT32), .B(G143), .Z(n1370) );
NAND2_X1 U1106 ( .A1(KEYINPUT2), .A2(n1276), .ZN(n1369) );
INV_X1 U1107 ( .A(G146), .ZN(n1276) );
XNOR2_X1 U1108 ( .A(n1371), .B(n1372), .ZN(n1171) );
XOR2_X1 U1109 ( .A(KEYINPUT8), .B(KEYINPUT43), .Z(n1372) );
XOR2_X1 U1110 ( .A(n1303), .B(G113), .Z(n1371) );
XNOR2_X1 U1111 ( .A(G116), .B(n1349), .ZN(n1303) );
XNOR2_X1 U1112 ( .A(n1260), .B(KEYINPUT37), .ZN(n1349) );
INV_X1 U1113 ( .A(G119), .ZN(n1260) );
XOR2_X1 U1114 ( .A(n1373), .B(G101), .Z(n1355) );
NAND2_X1 U1115 ( .A1(KEYINPUT51), .A2(n1374), .ZN(n1373) );
NAND2_X1 U1116 ( .A1(G210), .A2(n1179), .ZN(n1374) );
NOR2_X1 U1117 ( .A1(G953), .A2(G237), .ZN(n1179) );
endmodule


