//Key = 1011100100011000000110000110100111110011011100001100100111000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
n1472, n1473, n1474;

XOR2_X1 U794 ( .A(n1122), .B(n1123), .Z(G9) );
NAND2_X1 U795 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U796 ( .A1(KEYINPUT32), .A2(G107), .ZN(n1122) );
NAND3_X1 U797 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(G75) );
NAND2_X1 U798 ( .A1(G952), .A2(n1129), .ZN(n1128) );
NAND2_X1 U799 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U800 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U801 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NAND3_X1 U802 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
NAND2_X1 U803 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U804 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U805 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U806 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NAND2_X1 U807 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U808 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND3_X1 U809 ( .A1(n1145), .A2(n1151), .A3(n1141), .ZN(n1134) );
NAND2_X1 U810 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U811 ( .A1(n1138), .A2(n1154), .ZN(n1153) );
NAND2_X1 U812 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U813 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U814 ( .A(n1159), .ZN(n1155) );
NAND2_X1 U815 ( .A1(n1136), .A2(n1160), .ZN(n1152) );
NAND2_X1 U816 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U817 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U818 ( .A(n1165), .ZN(n1130) );
NAND4_X1 U819 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1126) );
NOR4_X1 U820 ( .A1(n1158), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1169) );
XOR2_X1 U821 ( .A(G469), .B(n1173), .Z(n1172) );
XOR2_X1 U822 ( .A(n1174), .B(n1175), .Z(n1171) );
XOR2_X1 U823 ( .A(G478), .B(n1176), .Z(n1170) );
NOR2_X1 U824 ( .A1(KEYINPUT30), .A2(n1177), .ZN(n1176) );
NOR3_X1 U825 ( .A1(n1163), .A2(n1178), .A3(n1149), .ZN(n1168) );
NAND2_X1 U826 ( .A1(n1179), .A2(n1180), .ZN(n1167) );
XNOR2_X1 U827 ( .A(KEYINPUT3), .B(n1181), .ZN(n1180) );
XNOR2_X1 U828 ( .A(G475), .B(KEYINPUT19), .ZN(n1179) );
XNOR2_X1 U829 ( .A(n1164), .B(KEYINPUT62), .ZN(n1166) );
XOR2_X1 U830 ( .A(n1182), .B(n1183), .Z(G72) );
NOR2_X1 U831 ( .A1(n1184), .A2(n1127), .ZN(n1183) );
AND2_X1 U832 ( .A1(G227), .A2(G900), .ZN(n1184) );
NAND2_X1 U833 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
NAND2_X1 U834 ( .A1(n1187), .A2(n1127), .ZN(n1186) );
XNOR2_X1 U835 ( .A(n1188), .B(n1189), .ZN(n1187) );
NAND3_X1 U836 ( .A1(G900), .A2(n1189), .A3(G953), .ZN(n1185) );
NAND3_X1 U837 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
NAND2_X1 U838 ( .A1(KEYINPUT22), .A2(n1193), .ZN(n1192) );
NAND3_X1 U839 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1191) );
INV_X1 U840 ( .A(KEYINPUT22), .ZN(n1195) );
OR2_X1 U841 ( .A1(n1196), .A2(n1194), .ZN(n1190) );
NOR2_X1 U842 ( .A1(n1197), .A2(n1193), .ZN(n1194) );
XNOR2_X1 U843 ( .A(n1198), .B(n1199), .ZN(n1193) );
INV_X1 U844 ( .A(n1200), .ZN(n1199) );
XNOR2_X1 U845 ( .A(KEYINPUT46), .B(n1201), .ZN(n1198) );
NOR2_X1 U846 ( .A1(KEYINPUT21), .A2(n1202), .ZN(n1201) );
INV_X1 U847 ( .A(KEYINPUT63), .ZN(n1197) );
AND2_X1 U848 ( .A1(n1203), .A2(n1204), .ZN(n1196) );
NAND2_X1 U849 ( .A1(KEYINPUT33), .A2(n1205), .ZN(n1204) );
NAND2_X1 U850 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U851 ( .A1(n1208), .A2(n1209), .ZN(n1203) );
INV_X1 U852 ( .A(KEYINPUT33), .ZN(n1209) );
XOR2_X1 U853 ( .A(n1210), .B(G125), .Z(n1208) );
NAND2_X1 U854 ( .A1(n1211), .A2(n1212), .ZN(G69) );
NAND2_X1 U855 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR2_X1 U856 ( .A1(n1127), .A2(G224), .ZN(n1214) );
INV_X1 U857 ( .A(n1215), .ZN(n1213) );
NAND3_X1 U858 ( .A1(G953), .A2(n1216), .A3(n1215), .ZN(n1211) );
XOR2_X1 U859 ( .A(n1217), .B(n1218), .Z(n1215) );
NOR2_X1 U860 ( .A1(n1219), .A2(G953), .ZN(n1218) );
NOR2_X1 U861 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U862 ( .A1(n1222), .A2(n1223), .ZN(n1217) );
NAND2_X1 U863 ( .A1(G953), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U864 ( .A(n1225), .B(n1226), .ZN(n1222) );
XNOR2_X1 U865 ( .A(n1227), .B(n1228), .ZN(n1225) );
NAND2_X1 U866 ( .A1(KEYINPUT48), .A2(n1229), .ZN(n1228) );
NAND2_X1 U867 ( .A1(KEYINPUT34), .A2(n1230), .ZN(n1227) );
NAND2_X1 U868 ( .A1(G898), .A2(G224), .ZN(n1216) );
NOR2_X1 U869 ( .A1(n1231), .A2(n1232), .ZN(G66) );
XOR2_X1 U870 ( .A(n1233), .B(n1234), .Z(n1232) );
NAND4_X1 U871 ( .A1(G217), .A2(n1235), .A3(n1236), .A4(n1165), .ZN(n1233) );
XOR2_X1 U872 ( .A(KEYINPUT38), .B(n1237), .Z(n1235) );
INV_X1 U873 ( .A(n1238), .ZN(n1237) );
NOR2_X1 U874 ( .A1(n1231), .A2(n1239), .ZN(G63) );
NOR2_X1 U875 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U876 ( .A(n1242), .B(KEYINPUT39), .Z(n1241) );
NAND2_X1 U877 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NOR2_X1 U878 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
AND2_X1 U879 ( .A1(n1245), .A2(G478), .ZN(n1243) );
NOR2_X1 U880 ( .A1(n1231), .A2(n1246), .ZN(G60) );
XNOR2_X1 U881 ( .A(n1247), .B(n1248), .ZN(n1246) );
AND2_X1 U882 ( .A1(G475), .A2(n1245), .ZN(n1248) );
NAND3_X1 U883 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(G6) );
NAND2_X1 U884 ( .A1(G104), .A2(n1252), .ZN(n1251) );
NAND2_X1 U885 ( .A1(KEYINPUT17), .A2(n1253), .ZN(n1250) );
NAND2_X1 U886 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U887 ( .A(n1252), .ZN(n1255) );
XNOR2_X1 U888 ( .A(KEYINPUT16), .B(G104), .ZN(n1254) );
NAND2_X1 U889 ( .A1(n1256), .A2(n1257), .ZN(n1249) );
INV_X1 U890 ( .A(KEYINPUT17), .ZN(n1257) );
NAND2_X1 U891 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
OR3_X1 U892 ( .A1(n1252), .A2(G104), .A3(KEYINPUT16), .ZN(n1259) );
NAND2_X1 U893 ( .A1(KEYINPUT16), .A2(G104), .ZN(n1258) );
NOR2_X1 U894 ( .A1(n1231), .A2(n1260), .ZN(G57) );
XOR2_X1 U895 ( .A(n1261), .B(n1262), .Z(n1260) );
NAND2_X1 U896 ( .A1(n1263), .A2(KEYINPUT43), .ZN(n1261) );
XOR2_X1 U897 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U898 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U899 ( .A1(n1174), .A2(n1268), .ZN(n1267) );
NOR2_X1 U900 ( .A1(KEYINPUT18), .A2(n1269), .ZN(n1266) );
XNOR2_X1 U901 ( .A(n1270), .B(n1271), .ZN(n1269) );
NOR2_X1 U902 ( .A1(n1231), .A2(n1272), .ZN(G54) );
XOR2_X1 U903 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U904 ( .A(n1200), .B(n1275), .Z(n1274) );
XOR2_X1 U905 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U906 ( .A(n1278), .B(n1279), .ZN(n1200) );
XOR2_X1 U907 ( .A(n1280), .B(n1281), .Z(n1273) );
XOR2_X1 U908 ( .A(n1282), .B(n1283), .Z(n1281) );
AND2_X1 U909 ( .A1(G469), .A2(n1245), .ZN(n1283) );
INV_X1 U910 ( .A(n1268), .ZN(n1245) );
NOR2_X1 U911 ( .A1(KEYINPUT6), .A2(n1284), .ZN(n1282) );
XOR2_X1 U912 ( .A(n1285), .B(KEYINPUT51), .Z(n1284) );
XOR2_X1 U913 ( .A(n1210), .B(KEYINPUT4), .Z(n1280) );
NOR2_X1 U914 ( .A1(n1231), .A2(n1286), .ZN(G51) );
XOR2_X1 U915 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U916 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR2_X1 U917 ( .A1(n1291), .A2(n1268), .ZN(n1290) );
NAND2_X1 U918 ( .A1(n1238), .A2(n1165), .ZN(n1268) );
NAND3_X1 U919 ( .A1(n1188), .A2(n1292), .A3(n1293), .ZN(n1165) );
XOR2_X1 U920 ( .A(n1220), .B(KEYINPUT25), .Z(n1293) );
NAND4_X1 U921 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1220) );
INV_X1 U922 ( .A(n1298), .ZN(n1297) );
NAND4_X1 U923 ( .A1(n1299), .A2(n1300), .A3(n1136), .A4(n1301), .ZN(n1295) );
NOR2_X1 U924 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U925 ( .A1(KEYINPUT31), .A2(n1304), .ZN(n1300) );
NAND2_X1 U926 ( .A1(n1305), .A2(n1306), .ZN(n1299) );
INV_X1 U927 ( .A(KEYINPUT31), .ZN(n1306) );
NAND2_X1 U928 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND3_X1 U929 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1294) );
XOR2_X1 U930 ( .A(KEYINPUT45), .B(n1159), .Z(n1310) );
INV_X1 U931 ( .A(n1221), .ZN(n1292) );
NAND4_X1 U932 ( .A1(n1312), .A2(n1252), .A3(n1313), .A4(n1314), .ZN(n1221) );
NAND2_X1 U933 ( .A1(n1309), .A2(n1125), .ZN(n1252) );
AND2_X1 U934 ( .A1(n1315), .A2(n1136), .ZN(n1125) );
NAND3_X1 U935 ( .A1(n1315), .A2(n1316), .A3(n1124), .ZN(n1312) );
XOR2_X1 U936 ( .A(KEYINPUT37), .B(n1136), .Z(n1316) );
AND4_X1 U937 ( .A1(n1317), .A2(n1318), .A3(n1319), .A4(n1320), .ZN(n1188) );
NOR4_X1 U938 ( .A1(n1321), .A2(n1322), .A3(n1323), .A4(n1324), .ZN(n1320) );
AND2_X1 U939 ( .A1(n1325), .A2(n1326), .ZN(n1319) );
XOR2_X1 U940 ( .A(n1327), .B(KEYINPUT20), .Z(n1238) );
XOR2_X1 U941 ( .A(n1328), .B(KEYINPUT44), .Z(n1291) );
NOR3_X1 U942 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1289) );
AND3_X1 U943 ( .A1(n1270), .A2(n1332), .A3(G125), .ZN(n1331) );
NOR3_X1 U944 ( .A1(n1270), .A2(n1333), .A3(n1332), .ZN(n1330) );
NOR2_X1 U945 ( .A1(G125), .A2(n1334), .ZN(n1329) );
NOR2_X1 U946 ( .A1(KEYINPUT5), .A2(n1335), .ZN(n1287) );
NOR2_X1 U947 ( .A1(n1127), .A2(G952), .ZN(n1231) );
XOR2_X1 U948 ( .A(G146), .B(n1324), .Z(G48) );
AND3_X1 U949 ( .A1(n1336), .A2(n1337), .A3(n1309), .ZN(n1324) );
XNOR2_X1 U950 ( .A(G143), .B(n1318), .ZN(G45) );
NAND4_X1 U951 ( .A1(n1338), .A2(n1337), .A3(n1339), .A4(n1340), .ZN(n1318) );
XOR2_X1 U952 ( .A(n1210), .B(n1326), .Z(G42) );
NAND3_X1 U953 ( .A1(n1138), .A2(n1341), .A3(n1342), .ZN(n1326) );
XOR2_X1 U954 ( .A(G137), .B(n1323), .Z(G39) );
AND3_X1 U955 ( .A1(n1336), .A2(n1145), .A3(n1138), .ZN(n1323) );
NAND2_X1 U956 ( .A1(n1343), .A2(n1344), .ZN(G36) );
OR2_X1 U957 ( .A1(n1325), .A2(G134), .ZN(n1344) );
XOR2_X1 U958 ( .A(n1345), .B(KEYINPUT23), .Z(n1343) );
NAND2_X1 U959 ( .A1(G134), .A2(n1325), .ZN(n1345) );
NAND3_X1 U960 ( .A1(n1338), .A2(n1124), .A3(n1138), .ZN(n1325) );
XOR2_X1 U961 ( .A(G131), .B(n1322), .Z(G33) );
AND3_X1 U962 ( .A1(n1309), .A2(n1338), .A3(n1138), .ZN(n1322) );
AND2_X1 U963 ( .A1(n1164), .A2(n1346), .ZN(n1138) );
AND3_X1 U964 ( .A1(n1341), .A2(n1347), .A3(n1159), .ZN(n1338) );
XOR2_X1 U965 ( .A(G128), .B(n1321), .Z(G30) );
AND3_X1 U966 ( .A1(n1124), .A2(n1337), .A3(n1336), .ZN(n1321) );
AND4_X1 U967 ( .A1(n1341), .A2(n1347), .A3(n1158), .A4(n1348), .ZN(n1336) );
INV_X1 U968 ( .A(n1143), .ZN(n1124) );
XNOR2_X1 U969 ( .A(G101), .B(n1313), .ZN(G3) );
NAND3_X1 U970 ( .A1(n1315), .A2(n1145), .A3(n1159), .ZN(n1313) );
XOR2_X1 U971 ( .A(n1333), .B(n1349), .Z(G27) );
NOR2_X1 U972 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NOR2_X1 U973 ( .A1(n1352), .A2(n1317), .ZN(n1351) );
NAND2_X1 U974 ( .A1(n1353), .A2(n1337), .ZN(n1317) );
INV_X1 U975 ( .A(KEYINPUT42), .ZN(n1352) );
NOR3_X1 U976 ( .A1(KEYINPUT42), .A2(n1353), .A3(n1161), .ZN(n1350) );
INV_X1 U977 ( .A(n1337), .ZN(n1161) );
AND2_X1 U978 ( .A1(n1141), .A2(n1342), .ZN(n1353) );
AND4_X1 U979 ( .A1(n1309), .A2(n1157), .A3(n1347), .A4(n1158), .ZN(n1342) );
NAND2_X1 U980 ( .A1(n1354), .A2(n1355), .ZN(n1347) );
NAND4_X1 U981 ( .A1(G953), .A2(G902), .A3(n1133), .A4(n1356), .ZN(n1355) );
INV_X1 U982 ( .A(G900), .ZN(n1356) );
INV_X1 U983 ( .A(n1144), .ZN(n1309) );
XNOR2_X1 U984 ( .A(G122), .B(n1357), .ZN(G24) );
NAND4_X1 U985 ( .A1(n1311), .A2(n1136), .A3(n1339), .A4(n1340), .ZN(n1357) );
NOR2_X1 U986 ( .A1(n1348), .A2(n1158), .ZN(n1136) );
XOR2_X1 U987 ( .A(n1358), .B(n1296), .Z(G21) );
NAND4_X1 U988 ( .A1(n1311), .A2(n1145), .A3(n1158), .A4(n1348), .ZN(n1296) );
XOR2_X1 U989 ( .A(G116), .B(n1298), .Z(G18) );
NOR2_X1 U990 ( .A1(n1359), .A2(n1143), .ZN(n1298) );
XOR2_X1 U991 ( .A(G113), .B(n1360), .Z(G15) );
NOR2_X1 U992 ( .A1(n1144), .A2(n1359), .ZN(n1360) );
NAND2_X1 U993 ( .A1(n1311), .A2(n1159), .ZN(n1359) );
NOR2_X1 U994 ( .A1(n1158), .A2(n1157), .ZN(n1159) );
INV_X1 U995 ( .A(n1304), .ZN(n1311) );
NAND2_X1 U996 ( .A1(n1141), .A2(n1307), .ZN(n1304) );
INV_X1 U997 ( .A(n1308), .ZN(n1141) );
NAND2_X1 U998 ( .A1(n1361), .A2(n1150), .ZN(n1308) );
INV_X1 U999 ( .A(n1362), .ZN(n1150) );
NAND2_X1 U1000 ( .A1(n1363), .A2(n1340), .ZN(n1144) );
INV_X1 U1001 ( .A(n1302), .ZN(n1340) );
XOR2_X1 U1002 ( .A(KEYINPUT12), .B(n1339), .Z(n1363) );
XOR2_X1 U1003 ( .A(n1364), .B(n1314), .Z(G12) );
NAND4_X1 U1004 ( .A1(n1315), .A2(n1157), .A3(n1145), .A4(n1158), .ZN(n1314) );
NAND3_X1 U1005 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1158) );
NAND2_X1 U1006 ( .A1(G902), .A2(G217), .ZN(n1367) );
NAND3_X1 U1007 ( .A1(n1234), .A2(n1327), .A3(n1368), .ZN(n1366) );
OR2_X1 U1008 ( .A1(n1368), .A2(n1234), .ZN(n1365) );
XNOR2_X1 U1009 ( .A(n1369), .B(n1370), .ZN(n1234) );
XNOR2_X1 U1010 ( .A(n1277), .B(n1371), .ZN(n1370) );
XOR2_X1 U1011 ( .A(n1372), .B(n1373), .Z(n1371) );
AND3_X1 U1012 ( .A1(G221), .A2(n1127), .A3(G234), .ZN(n1373) );
NAND2_X1 U1013 ( .A1(n1374), .A2(n1206), .ZN(n1372) );
XOR2_X1 U1014 ( .A(n1207), .B(KEYINPUT47), .Z(n1374) );
XOR2_X1 U1015 ( .A(n1364), .B(n1202), .Z(n1277) );
XOR2_X1 U1016 ( .A(n1375), .B(n1376), .Z(n1369) );
XOR2_X1 U1017 ( .A(G128), .B(n1377), .Z(n1376) );
NOR2_X1 U1018 ( .A1(G119), .A2(KEYINPUT61), .ZN(n1377) );
XNOR2_X1 U1019 ( .A(G146), .B(KEYINPUT58), .ZN(n1375) );
NAND2_X1 U1020 ( .A1(G217), .A2(n1378), .ZN(n1368) );
INV_X1 U1021 ( .A(G234), .ZN(n1378) );
NAND2_X1 U1022 ( .A1(n1379), .A2(n1380), .ZN(n1145) );
OR2_X1 U1023 ( .A1(n1143), .A2(KEYINPUT12), .ZN(n1380) );
NAND2_X1 U1024 ( .A1(n1302), .A2(n1339), .ZN(n1143) );
INV_X1 U1025 ( .A(n1303), .ZN(n1339) );
NAND3_X1 U1026 ( .A1(n1302), .A2(n1303), .A3(KEYINPUT12), .ZN(n1379) );
XOR2_X1 U1027 ( .A(n1177), .B(G478), .Z(n1303) );
OR2_X1 U1028 ( .A1(n1244), .A2(G902), .ZN(n1177) );
XNOR2_X1 U1029 ( .A(n1381), .B(n1382), .ZN(n1244) );
XOR2_X1 U1030 ( .A(n1383), .B(n1384), .Z(n1382) );
XOR2_X1 U1031 ( .A(G128), .B(G122), .Z(n1384) );
XOR2_X1 U1032 ( .A(G143), .B(G134), .Z(n1383) );
XOR2_X1 U1033 ( .A(n1385), .B(n1386), .Z(n1381) );
XOR2_X1 U1034 ( .A(G107), .B(n1387), .Z(n1386) );
AND3_X1 U1035 ( .A1(G234), .A2(n1127), .A3(G217), .ZN(n1387) );
NAND2_X1 U1036 ( .A1(KEYINPUT41), .A2(n1388), .ZN(n1385) );
NOR2_X1 U1037 ( .A1(n1178), .A2(n1389), .ZN(n1302) );
AND2_X1 U1038 ( .A1(G475), .A2(n1181), .ZN(n1389) );
NOR2_X1 U1039 ( .A1(n1181), .A2(G475), .ZN(n1178) );
NAND2_X1 U1040 ( .A1(n1247), .A2(n1327), .ZN(n1181) );
XNOR2_X1 U1041 ( .A(n1390), .B(n1391), .ZN(n1247) );
XOR2_X1 U1042 ( .A(n1392), .B(n1393), .Z(n1391) );
XOR2_X1 U1043 ( .A(n1394), .B(n1395), .Z(n1393) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1396), .ZN(n1394) );
XOR2_X1 U1045 ( .A(n1397), .B(n1398), .Z(n1392) );
NOR2_X1 U1046 ( .A1(G122), .A2(KEYINPUT40), .ZN(n1398) );
NAND3_X1 U1047 ( .A1(n1399), .A2(n1400), .A3(n1207), .ZN(n1397) );
NAND2_X1 U1048 ( .A1(G125), .A2(n1210), .ZN(n1207) );
OR2_X1 U1049 ( .A1(n1333), .A2(KEYINPUT11), .ZN(n1400) );
NAND2_X1 U1050 ( .A1(n1401), .A2(KEYINPUT11), .ZN(n1399) );
INV_X1 U1051 ( .A(n1206), .ZN(n1401) );
NAND2_X1 U1052 ( .A1(G140), .A2(n1333), .ZN(n1206) );
XOR2_X1 U1053 ( .A(n1402), .B(n1403), .Z(n1390) );
XOR2_X1 U1054 ( .A(G113), .B(G104), .Z(n1403) );
XNOR2_X1 U1055 ( .A(G131), .B(KEYINPUT58), .ZN(n1402) );
INV_X1 U1056 ( .A(n1348), .ZN(n1157) );
NAND3_X1 U1057 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n1348) );
NAND2_X1 U1058 ( .A1(n1407), .A2(n1174), .ZN(n1406) );
OR3_X1 U1059 ( .A1(n1174), .A2(n1407), .A3(n1408), .ZN(n1405) );
NOR2_X1 U1060 ( .A1(n1409), .A2(n1175), .ZN(n1407) );
INV_X1 U1061 ( .A(KEYINPUT7), .ZN(n1409) );
INV_X1 U1062 ( .A(G472), .ZN(n1174) );
NAND2_X1 U1063 ( .A1(n1410), .A2(n1408), .ZN(n1404) );
INV_X1 U1064 ( .A(KEYINPUT49), .ZN(n1408) );
NAND2_X1 U1065 ( .A1(G472), .A2(n1175), .ZN(n1410) );
NAND2_X1 U1066 ( .A1(n1411), .A2(n1327), .ZN(n1175) );
XOR2_X1 U1067 ( .A(n1412), .B(n1413), .Z(n1411) );
XOR2_X1 U1068 ( .A(n1262), .B(n1270), .Z(n1413) );
XOR2_X1 U1069 ( .A(n1414), .B(n1415), .Z(n1262) );
NAND2_X1 U1070 ( .A1(G210), .A2(n1396), .ZN(n1414) );
NOR2_X1 U1071 ( .A1(G953), .A2(G237), .ZN(n1396) );
XOR2_X1 U1072 ( .A(n1264), .B(n1416), .Z(n1412) );
XNOR2_X1 U1073 ( .A(KEYINPUT8), .B(n1417), .ZN(n1416) );
NOR2_X1 U1074 ( .A1(KEYINPUT1), .A2(n1271), .ZN(n1417) );
XOR2_X1 U1075 ( .A(n1418), .B(n1419), .Z(n1264) );
XOR2_X1 U1076 ( .A(G119), .B(G113), .Z(n1419) );
NAND2_X1 U1077 ( .A1(KEYINPUT52), .A2(G116), .ZN(n1418) );
AND2_X1 U1078 ( .A1(n1341), .A2(n1307), .ZN(n1315) );
AND2_X1 U1079 ( .A1(n1337), .A2(n1420), .ZN(n1307) );
NAND2_X1 U1080 ( .A1(n1421), .A2(n1354), .ZN(n1420) );
NAND3_X1 U1081 ( .A1(G952), .A2(n1127), .A3(n1422), .ZN(n1354) );
XOR2_X1 U1082 ( .A(n1133), .B(KEYINPUT14), .Z(n1422) );
NAND4_X1 U1083 ( .A1(G953), .A2(G902), .A3(n1133), .A4(n1224), .ZN(n1421) );
INV_X1 U1084 ( .A(G898), .ZN(n1224) );
NAND2_X1 U1085 ( .A1(G237), .A2(G234), .ZN(n1133) );
NOR2_X1 U1086 ( .A1(n1164), .A2(n1163), .ZN(n1337) );
INV_X1 U1087 ( .A(n1346), .ZN(n1163) );
NAND2_X1 U1088 ( .A1(G214), .A2(n1423), .ZN(n1346) );
XNOR2_X1 U1089 ( .A(n1424), .B(n1425), .ZN(n1164) );
NOR2_X1 U1090 ( .A1(n1426), .A2(n1427), .ZN(n1425) );
NOR2_X1 U1091 ( .A1(n1428), .A2(n1328), .ZN(n1427) );
NAND2_X1 U1092 ( .A1(G210), .A2(n1423), .ZN(n1328) );
INV_X1 U1093 ( .A(KEYINPUT0), .ZN(n1428) );
NOR3_X1 U1094 ( .A1(KEYINPUT0), .A2(n1429), .A3(n1423), .ZN(n1426) );
NAND2_X1 U1095 ( .A1(n1430), .A2(n1327), .ZN(n1423) );
XNOR2_X1 U1096 ( .A(G237), .B(KEYINPUT27), .ZN(n1430) );
INV_X1 U1097 ( .A(G210), .ZN(n1429) );
NAND2_X1 U1098 ( .A1(n1431), .A2(n1327), .ZN(n1424) );
XOR2_X1 U1099 ( .A(n1432), .B(n1433), .Z(n1431) );
XNOR2_X1 U1100 ( .A(n1335), .B(n1334), .ZN(n1433) );
XNOR2_X1 U1101 ( .A(n1270), .B(n1332), .ZN(n1334) );
NAND2_X1 U1102 ( .A1(G224), .A2(n1127), .ZN(n1332) );
NAND2_X1 U1103 ( .A1(n1434), .A2(n1435), .ZN(n1270) );
NAND2_X1 U1104 ( .A1(n1436), .A2(n1437), .ZN(n1435) );
INV_X1 U1105 ( .A(G128), .ZN(n1437) );
NAND2_X1 U1106 ( .A1(n1395), .A2(n1438), .ZN(n1436) );
OR2_X1 U1107 ( .A1(KEYINPUT35), .A2(KEYINPUT29), .ZN(n1438) );
NAND3_X1 U1108 ( .A1(KEYINPUT35), .A2(n1439), .A3(G128), .ZN(n1434) );
XOR2_X1 U1109 ( .A(KEYINPUT29), .B(n1395), .Z(n1439) );
XNOR2_X1 U1110 ( .A(n1229), .B(n1440), .ZN(n1335) );
XOR2_X1 U1111 ( .A(n1230), .B(n1441), .Z(n1440) );
NOR2_X1 U1112 ( .A1(KEYINPUT59), .A2(n1226), .ZN(n1441) );
XOR2_X1 U1113 ( .A(n1442), .B(G104), .Z(n1226) );
AND2_X1 U1114 ( .A1(n1443), .A2(n1444), .ZN(n1230) );
NAND2_X1 U1115 ( .A1(G122), .A2(n1364), .ZN(n1444) );
XOR2_X1 U1116 ( .A(n1445), .B(KEYINPUT36), .Z(n1443) );
OR2_X1 U1117 ( .A1(n1364), .A2(G122), .ZN(n1445) );
XOR2_X1 U1118 ( .A(n1446), .B(G113), .Z(n1229) );
NAND4_X1 U1119 ( .A1(n1447), .A2(n1448), .A3(n1449), .A4(n1450), .ZN(n1446) );
NAND3_X1 U1120 ( .A1(n1451), .A2(n1358), .A3(n1452), .ZN(n1450) );
INV_X1 U1121 ( .A(KEYINPUT15), .ZN(n1452) );
XNOR2_X1 U1122 ( .A(KEYINPUT24), .B(n1453), .ZN(n1451) );
NAND2_X1 U1123 ( .A1(G119), .A2(KEYINPUT15), .ZN(n1449) );
OR3_X1 U1124 ( .A1(n1453), .A2(n1454), .A3(KEYINPUT56), .ZN(n1448) );
AND2_X1 U1125 ( .A1(KEYINPUT24), .A2(n1358), .ZN(n1454) );
INV_X1 U1126 ( .A(G119), .ZN(n1358) );
NAND3_X1 U1127 ( .A1(n1453), .A2(n1455), .A3(KEYINPUT56), .ZN(n1447) );
OR2_X1 U1128 ( .A1(KEYINPUT24), .A2(G119), .ZN(n1455) );
XNOR2_X1 U1129 ( .A(n1388), .B(KEYINPUT10), .ZN(n1453) );
INV_X1 U1130 ( .A(G116), .ZN(n1388) );
XNOR2_X1 U1131 ( .A(n1456), .B(KEYINPUT54), .ZN(n1432) );
NAND2_X1 U1132 ( .A1(KEYINPUT26), .A2(n1333), .ZN(n1456) );
INV_X1 U1133 ( .A(G125), .ZN(n1333) );
INV_X1 U1134 ( .A(n1147), .ZN(n1341) );
NAND2_X1 U1135 ( .A1(n1361), .A2(n1362), .ZN(n1147) );
XNOR2_X1 U1136 ( .A(G469), .B(n1457), .ZN(n1362) );
NOR2_X1 U1137 ( .A1(n1173), .A2(KEYINPUT50), .ZN(n1457) );
AND3_X1 U1138 ( .A1(n1458), .A2(n1459), .A3(n1327), .ZN(n1173) );
NAND2_X1 U1139 ( .A1(n1460), .A2(n1210), .ZN(n1459) );
INV_X1 U1140 ( .A(G140), .ZN(n1210) );
NAND2_X1 U1141 ( .A1(n1461), .A2(G140), .ZN(n1458) );
XNOR2_X1 U1142 ( .A(KEYINPUT60), .B(n1460), .ZN(n1461) );
XNOR2_X1 U1143 ( .A(n1462), .B(n1285), .ZN(n1460) );
NAND2_X1 U1144 ( .A1(G227), .A2(n1127), .ZN(n1285) );
INV_X1 U1145 ( .A(G953), .ZN(n1127) );
XOR2_X1 U1146 ( .A(n1463), .B(G110), .Z(n1462) );
NAND3_X1 U1147 ( .A1(n1464), .A2(n1465), .A3(n1466), .ZN(n1463) );
NAND2_X1 U1148 ( .A1(n1271), .A2(n1467), .ZN(n1466) );
OR3_X1 U1149 ( .A1(n1467), .A2(n1271), .A3(n1468), .ZN(n1465) );
INV_X1 U1150 ( .A(KEYINPUT55), .ZN(n1467) );
NAND2_X1 U1151 ( .A1(n1468), .A2(n1469), .ZN(n1464) );
NAND2_X1 U1152 ( .A1(n1470), .A2(KEYINPUT55), .ZN(n1469) );
XOR2_X1 U1153 ( .A(n1271), .B(KEYINPUT28), .Z(n1470) );
XOR2_X1 U1154 ( .A(n1202), .B(n1278), .Z(n1271) );
XOR2_X1 U1155 ( .A(G131), .B(G134), .Z(n1278) );
INV_X1 U1156 ( .A(G137), .ZN(n1202) );
XNOR2_X1 U1157 ( .A(n1471), .B(n1472), .ZN(n1468) );
INV_X1 U1158 ( .A(n1276), .ZN(n1472) );
XOR2_X1 U1159 ( .A(n1442), .B(n1473), .Z(n1276) );
NOR2_X1 U1160 ( .A1(G104), .A2(KEYINPUT53), .ZN(n1473) );
XNOR2_X1 U1161 ( .A(G107), .B(n1415), .ZN(n1442) );
XOR2_X1 U1162 ( .A(G101), .B(KEYINPUT9), .Z(n1415) );
NAND2_X1 U1163 ( .A1(KEYINPUT57), .A2(n1279), .ZN(n1471) );
XOR2_X1 U1164 ( .A(G128), .B(n1395), .Z(n1279) );
XOR2_X1 U1165 ( .A(G143), .B(G146), .Z(n1395) );
XNOR2_X1 U1166 ( .A(n1149), .B(KEYINPUT13), .ZN(n1361) );
AND2_X1 U1167 ( .A1(n1474), .A2(n1236), .ZN(n1149) );
NAND2_X1 U1168 ( .A1(G234), .A2(n1327), .ZN(n1236) );
INV_X1 U1169 ( .A(G902), .ZN(n1327) );
XNOR2_X1 U1170 ( .A(G221), .B(KEYINPUT2), .ZN(n1474) );
INV_X1 U1171 ( .A(G110), .ZN(n1364) );
endmodule


