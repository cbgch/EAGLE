//Key = 1010110000100000100111010110000110101001100101001110111010010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307;

XNOR2_X1 U723 ( .A(G107), .B(n994), .ZN(G9) );
NOR2_X1 U724 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U725 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n996) );
INV_X1 U726 ( .A(G952), .ZN(n1000) );
XOR2_X1 U727 ( .A(n1001), .B(KEYINPUT57), .Z(n999) );
NAND2_X1 U728 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND3_X1 U729 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NAND2_X1 U730 ( .A1(KEYINPUT13), .A2(n1007), .ZN(n1005) );
NAND2_X1 U731 ( .A1(n1008), .A2(n1009), .ZN(n1004) );
INV_X1 U732 ( .A(KEYINPUT13), .ZN(n1009) );
OR2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NAND2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(n1002) );
NAND2_X1 U735 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND4_X1 U736 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1015) );
AND2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
XNOR2_X1 U738 ( .A(n1022), .B(KEYINPUT43), .ZN(n1016) );
NAND3_X1 U739 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND3_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1019), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1029), .A2(n1020), .ZN(n1025) );
INV_X1 U743 ( .A(n1030), .ZN(n998) );
NAND4_X1 U744 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n997) );
NAND3_X1 U745 ( .A1(n1022), .A2(n1035), .A3(n1012), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U747 ( .A1(n1019), .A2(n1038), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1020), .A2(n1041), .ZN(n1040) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1024), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1031) );
XNOR2_X1 U753 ( .A(n1006), .B(KEYINPUT54), .ZN(n1045) );
AND3_X1 U754 ( .A1(n1019), .A2(n1044), .A3(n1012), .ZN(n1006) );
INV_X1 U755 ( .A(n1047), .ZN(n1012) );
NOR3_X1 U756 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n995) );
NOR2_X1 U757 ( .A1(KEYINPUT9), .A2(n1051), .ZN(n1050) );
NOR2_X1 U758 ( .A1(G953), .A2(G952), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
INV_X1 U760 ( .A(KEYINPUT9), .ZN(n1053) );
INV_X1 U761 ( .A(n1033), .ZN(n1048) );
NAND4_X1 U762 ( .A1(n1044), .A2(n1022), .A3(n1054), .A4(n1055), .ZN(n1033) );
XNOR2_X1 U763 ( .A(n1056), .B(n1057), .ZN(n1055) );
NAND2_X1 U764 ( .A1(KEYINPUT10), .A2(n1058), .ZN(n1057) );
XNOR2_X1 U765 ( .A(n1059), .B(n1060), .ZN(n1054) );
XNOR2_X1 U766 ( .A(G478), .B(KEYINPUT20), .ZN(n1060) );
XOR2_X1 U767 ( .A(n1061), .B(n1062), .Z(G72) );
XOR2_X1 U768 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U769 ( .A1(n1065), .A2(G953), .ZN(n1064) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
NAND2_X1 U772 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U773 ( .A(n1072), .B(n1073), .Z(n1068) );
XNOR2_X1 U774 ( .A(KEYINPUT26), .B(n1074), .ZN(n1073) );
XOR2_X1 U775 ( .A(n1075), .B(n1076), .Z(n1072) );
NOR2_X1 U776 ( .A1(KEYINPUT15), .A2(n1077), .ZN(n1076) );
NAND2_X1 U777 ( .A1(G953), .A2(n1078), .ZN(n1061) );
NAND2_X1 U778 ( .A1(G900), .A2(G227), .ZN(n1078) );
XOR2_X1 U779 ( .A(n1079), .B(n1080), .Z(G69) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U782 ( .A(n1085), .B(KEYINPUT34), .Z(n1084) );
NAND3_X1 U783 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NAND2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
OR3_X1 U785 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1087) );
INV_X1 U786 ( .A(KEYINPUT0), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1091), .ZN(n1086) );
NAND2_X1 U788 ( .A1(KEYINPUT16), .A2(n1093), .ZN(n1091) );
AND2_X1 U789 ( .A1(n1094), .A2(n1070), .ZN(n1083) );
NAND2_X1 U790 ( .A1(G953), .A2(n1095), .ZN(n1081) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1095) );
NAND2_X1 U792 ( .A1(n1034), .A2(n1096), .ZN(n1079) );
NOR3_X1 U793 ( .A1(n1052), .A2(n1097), .A3(n1098), .ZN(G66) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U795 ( .A(KEYINPUT19), .B(n1101), .Z(n1100) );
INV_X1 U796 ( .A(n1102), .ZN(n1099) );
NOR2_X1 U797 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
NAND2_X1 U798 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1052), .A2(n1105), .ZN(G63) );
NOR3_X1 U800 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NOR2_X1 U801 ( .A1(KEYINPUT28), .A2(n1109), .ZN(n1108) );
NOR2_X1 U802 ( .A1(n1110), .A2(n1059), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1030), .A2(n1113), .ZN(n1112) );
AND2_X1 U805 ( .A1(KEYINPUT28), .A2(n1111), .ZN(n1107) );
NOR3_X1 U806 ( .A1(n1114), .A2(n1115), .A3(n1113), .ZN(n1106) );
XNOR2_X1 U807 ( .A(G478), .B(KEYINPUT18), .ZN(n1113) );
NOR2_X1 U808 ( .A1(n1111), .A2(KEYINPUT28), .ZN(n1115) );
INV_X1 U809 ( .A(n1103), .ZN(n1114) );
NOR2_X1 U810 ( .A1(n1052), .A2(n1116), .ZN(G60) );
NOR3_X1 U811 ( .A1(n1056), .A2(n1117), .A3(n1118), .ZN(n1116) );
AND3_X1 U812 ( .A1(n1119), .A2(n1103), .A3(G475), .ZN(n1118) );
NOR2_X1 U813 ( .A1(n1120), .A2(n1119), .ZN(n1117) );
NOR2_X1 U814 ( .A1(n1030), .A2(n1058), .ZN(n1120) );
INV_X1 U815 ( .A(G475), .ZN(n1058) );
XOR2_X1 U816 ( .A(G104), .B(n1121), .Z(G6) );
NOR2_X1 U817 ( .A1(n1052), .A2(n1122), .ZN(G57) );
XOR2_X1 U818 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U819 ( .A(KEYINPUT39), .B(n1125), .Z(n1124) );
NOR2_X1 U820 ( .A1(KEYINPUT7), .A2(n1126), .ZN(n1125) );
XOR2_X1 U821 ( .A(n1127), .B(n1128), .Z(n1123) );
AND2_X1 U822 ( .A1(G472), .A2(n1103), .ZN(n1128) );
NOR2_X1 U823 ( .A1(n1052), .A2(n1129), .ZN(G54) );
XOR2_X1 U824 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U825 ( .A(n1132), .B(n1133), .Z(n1131) );
AND2_X1 U826 ( .A1(G469), .A2(n1103), .ZN(n1133) );
NOR2_X1 U827 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XOR2_X1 U828 ( .A(n1136), .B(KEYINPUT5), .Z(n1135) );
NAND2_X1 U829 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U830 ( .A(n1139), .B(KEYINPUT24), .Z(n1137) );
NOR2_X1 U831 ( .A1(n1140), .A2(n1138), .ZN(n1134) );
XNOR2_X1 U832 ( .A(n1141), .B(G110), .ZN(n1138) );
XOR2_X1 U833 ( .A(n1139), .B(KEYINPUT3), .Z(n1140) );
NAND3_X1 U834 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1130) );
OR2_X1 U835 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND3_X1 U836 ( .A1(n1147), .A2(n1145), .A3(n1077), .ZN(n1143) );
INV_X1 U837 ( .A(KEYINPUT60), .ZN(n1145) );
OR2_X1 U838 ( .A1(n1077), .A2(n1147), .ZN(n1142) );
AND2_X1 U839 ( .A1(KEYINPUT36), .A2(n1146), .ZN(n1147) );
XNOR2_X1 U840 ( .A(n1148), .B(n1149), .ZN(n1146) );
XNOR2_X1 U841 ( .A(G101), .B(n1150), .ZN(n1148) );
NOR2_X1 U842 ( .A1(n1052), .A2(n1151), .ZN(G51) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U844 ( .A(n1154), .B(KEYINPUT63), .Z(n1153) );
NAND2_X1 U845 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U846 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
XNOR2_X1 U847 ( .A(n1157), .B(n1158), .ZN(n1156) );
XNOR2_X1 U848 ( .A(G125), .B(n1159), .ZN(n1158) );
XNOR2_X1 U849 ( .A(n1160), .B(n1126), .ZN(n1157) );
AND2_X1 U850 ( .A1(n1103), .A2(G210), .ZN(n1155) );
NOR2_X1 U851 ( .A1(n1161), .A2(n1030), .ZN(n1103) );
NOR3_X1 U852 ( .A1(n1096), .A2(n1067), .A3(n1162), .ZN(n1030) );
XNOR2_X1 U853 ( .A(n1066), .B(KEYINPUT40), .ZN(n1162) );
NAND4_X1 U854 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1066) );
NAND3_X1 U855 ( .A1(n1019), .A2(n1022), .A3(n1167), .ZN(n1163) );
NAND4_X1 U856 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1067) );
NAND2_X1 U857 ( .A1(n1172), .A2(n1173), .ZN(n1096) );
NOR4_X1 U858 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1121), .ZN(n1173) );
AND3_X1 U859 ( .A1(n1020), .A2(n1177), .A3(n1043), .ZN(n1121) );
AND4_X1 U860 ( .A1(n994), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1172) );
NAND3_X1 U861 ( .A1(n1020), .A2(n1177), .A3(n1029), .ZN(n994) );
NOR2_X1 U862 ( .A1(n1034), .A2(G952), .ZN(n1052) );
XNOR2_X1 U863 ( .A(G146), .B(n1164), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1043), .A2(n1046), .A3(n1167), .ZN(n1164) );
XNOR2_X1 U865 ( .A(G143), .B(n1165), .ZN(G45) );
NAND4_X1 U866 ( .A1(n1181), .A2(n1042), .A3(n1182), .A4(n1183), .ZN(n1165) );
AND2_X1 U867 ( .A1(n1046), .A2(n1184), .ZN(n1182) );
NAND2_X1 U868 ( .A1(n1185), .A2(n1186), .ZN(G42) );
OR2_X1 U869 ( .A1(n1166), .A2(G140), .ZN(n1186) );
XOR2_X1 U870 ( .A(n1187), .B(KEYINPUT51), .Z(n1185) );
NAND2_X1 U871 ( .A1(G140), .A2(n1166), .ZN(n1187) );
NAND2_X1 U872 ( .A1(n1188), .A2(n1189), .ZN(n1166) );
XOR2_X1 U873 ( .A(G137), .B(n1190), .Z(G39) );
NOR3_X1 U874 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
INV_X1 U875 ( .A(n1019), .ZN(n1193) );
XNOR2_X1 U876 ( .A(n1022), .B(KEYINPUT8), .ZN(n1192) );
XNOR2_X1 U877 ( .A(G134), .B(n1168), .ZN(G36) );
NAND3_X1 U878 ( .A1(n1042), .A2(n1029), .A3(n1188), .ZN(n1168) );
XNOR2_X1 U879 ( .A(G131), .B(n1169), .ZN(G33) );
NAND3_X1 U880 ( .A1(n1043), .A2(n1042), .A3(n1188), .ZN(n1169) );
AND2_X1 U881 ( .A1(n1181), .A2(n1022), .ZN(n1188) );
XNOR2_X1 U882 ( .A(G128), .B(n1170), .ZN(G30) );
NAND3_X1 U883 ( .A1(n1029), .A2(n1046), .A3(n1167), .ZN(n1170) );
INV_X1 U884 ( .A(n1191), .ZN(n1167) );
NAND3_X1 U885 ( .A1(n1194), .A2(n1028), .A3(n1181), .ZN(n1191) );
AND2_X1 U886 ( .A1(n1041), .A2(n1195), .ZN(n1181) );
XOR2_X1 U887 ( .A(n1196), .B(n1176), .Z(G3) );
AND3_X1 U888 ( .A1(n1042), .A2(n1177), .A3(n1019), .ZN(n1176) );
AND2_X1 U889 ( .A1(n1197), .A2(n1041), .ZN(n1177) );
NAND2_X1 U890 ( .A1(KEYINPUT23), .A2(n1198), .ZN(n1196) );
XOR2_X1 U891 ( .A(n1171), .B(n1199), .Z(G27) );
NOR2_X1 U892 ( .A1(G125), .A2(KEYINPUT58), .ZN(n1199) );
NAND4_X1 U893 ( .A1(n1189), .A2(n1024), .A3(n1046), .A4(n1195), .ZN(n1171) );
NAND2_X1 U894 ( .A1(n1047), .A2(n1200), .ZN(n1195) );
NAND4_X1 U895 ( .A1(G902), .A2(n1070), .A3(n1201), .A4(n1071), .ZN(n1200) );
INV_X1 U896 ( .A(G900), .ZN(n1071) );
AND3_X1 U897 ( .A1(n1027), .A2(n1028), .A3(n1043), .ZN(n1189) );
XNOR2_X1 U898 ( .A(G122), .B(n1180), .ZN(G24) );
NAND4_X1 U899 ( .A1(n1183), .A2(n1044), .A3(n1184), .A4(n1197), .ZN(n1180) );
AND2_X1 U900 ( .A1(n1024), .A2(n1020), .ZN(n1044) );
NOR2_X1 U901 ( .A1(n1028), .A2(n1194), .ZN(n1020) );
XNOR2_X1 U902 ( .A(G119), .B(n1179), .ZN(G21) );
NAND3_X1 U903 ( .A1(n1024), .A2(n1194), .A3(n1202), .ZN(n1179) );
XOR2_X1 U904 ( .A(G116), .B(n1175), .Z(G18) );
AND2_X1 U905 ( .A1(n1203), .A2(n1029), .ZN(n1175) );
AND2_X1 U906 ( .A1(n1184), .A2(n1204), .ZN(n1029) );
XNOR2_X1 U907 ( .A(n1205), .B(n1174), .ZN(G15) );
AND2_X1 U908 ( .A1(n1043), .A2(n1203), .ZN(n1174) );
AND3_X1 U909 ( .A1(n1024), .A2(n1197), .A3(n1042), .ZN(n1203) );
NOR2_X1 U910 ( .A1(n1028), .A2(n1027), .ZN(n1042) );
NOR2_X1 U911 ( .A1(n1206), .A2(n1017), .ZN(n1024) );
NOR2_X1 U912 ( .A1(n1204), .A2(n1184), .ZN(n1043) );
XNOR2_X1 U913 ( .A(G110), .B(n1178), .ZN(G12) );
NAND3_X1 U914 ( .A1(n1027), .A2(n1041), .A3(n1202), .ZN(n1178) );
AND3_X1 U915 ( .A1(n1197), .A2(n1028), .A3(n1019), .ZN(n1202) );
NOR2_X1 U916 ( .A1(n1184), .A2(n1183), .ZN(n1019) );
INV_X1 U917 ( .A(n1204), .ZN(n1183) );
XOR2_X1 U918 ( .A(n1056), .B(n1207), .Z(n1204) );
NOR2_X1 U919 ( .A1(G475), .A2(KEYINPUT46), .ZN(n1207) );
NOR2_X1 U920 ( .A1(n1119), .A2(G902), .ZN(n1056) );
XOR2_X1 U921 ( .A(n1208), .B(n1209), .Z(n1119) );
NOR2_X1 U922 ( .A1(KEYINPUT38), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U923 ( .A(G113), .B(G122), .ZN(n1210) );
XNOR2_X1 U924 ( .A(G104), .B(n1211), .ZN(n1208) );
NOR3_X1 U925 ( .A1(n1212), .A2(KEYINPUT6), .A3(n1213), .ZN(n1211) );
NOR2_X1 U926 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U927 ( .A(KEYINPUT42), .B(n1216), .Z(n1212) );
NOR2_X1 U928 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XNOR2_X1 U929 ( .A(n1214), .B(KEYINPUT37), .ZN(n1218) );
XOR2_X1 U930 ( .A(n1219), .B(n1220), .Z(n1214) );
INV_X1 U931 ( .A(G131), .ZN(n1220) );
NAND2_X1 U932 ( .A1(n1221), .A2(KEYINPUT32), .ZN(n1219) );
XNOR2_X1 U933 ( .A(n1222), .B(n1074), .ZN(n1221) );
NAND2_X1 U934 ( .A1(G214), .A2(n1223), .ZN(n1222) );
INV_X1 U935 ( .A(n1215), .ZN(n1217) );
XNOR2_X1 U936 ( .A(n1224), .B(n1225), .ZN(n1215) );
XNOR2_X1 U937 ( .A(KEYINPUT49), .B(n1226), .ZN(n1225) );
NAND3_X1 U938 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1224) );
NAND2_X1 U939 ( .A1(KEYINPUT35), .A2(G125), .ZN(n1229) );
NAND3_X1 U940 ( .A1(n1230), .A2(n1231), .A3(n1141), .ZN(n1228) );
INV_X1 U941 ( .A(KEYINPUT35), .ZN(n1231) );
OR2_X1 U942 ( .A1(n1141), .A2(n1230), .ZN(n1227) );
NOR2_X1 U943 ( .A1(G125), .A2(KEYINPUT29), .ZN(n1230) );
INV_X1 U944 ( .A(G140), .ZN(n1141) );
XOR2_X1 U945 ( .A(n1232), .B(G478), .Z(n1184) );
NAND2_X1 U946 ( .A1(KEYINPUT21), .A2(n1233), .ZN(n1232) );
XOR2_X1 U947 ( .A(KEYINPUT52), .B(n1059), .Z(n1233) );
NOR2_X1 U948 ( .A1(n1111), .A2(G902), .ZN(n1059) );
AND2_X1 U949 ( .A1(n1234), .A2(n1235), .ZN(n1111) );
NAND3_X1 U950 ( .A1(n1236), .A2(n1237), .A3(G217), .ZN(n1235) );
XNOR2_X1 U951 ( .A(n1238), .B(n1239), .ZN(n1237) );
NAND2_X1 U952 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
NAND2_X1 U953 ( .A1(G217), .A2(n1236), .ZN(n1241) );
XNOR2_X1 U954 ( .A(n1238), .B(n1242), .ZN(n1240) );
INV_X1 U955 ( .A(n1239), .ZN(n1242) );
XNOR2_X1 U956 ( .A(n1243), .B(n1244), .ZN(n1239) );
NAND2_X1 U957 ( .A1(KEYINPUT2), .A2(n1245), .ZN(n1243) );
XOR2_X1 U958 ( .A(n1246), .B(n1247), .Z(n1238) );
NOR2_X1 U959 ( .A1(KEYINPUT11), .A2(n1248), .ZN(n1247) );
XOR2_X1 U960 ( .A(G122), .B(G116), .Z(n1248) );
XNOR2_X1 U961 ( .A(G128), .B(G143), .ZN(n1246) );
XNOR2_X1 U962 ( .A(n1249), .B(n1104), .ZN(n1028) );
AND2_X1 U963 ( .A1(G217), .A2(n1250), .ZN(n1104) );
OR2_X1 U964 ( .A1(n1101), .A2(G902), .ZN(n1249) );
XNOR2_X1 U965 ( .A(n1251), .B(n1252), .ZN(n1101) );
XNOR2_X1 U966 ( .A(n1253), .B(n1254), .ZN(n1252) );
XOR2_X1 U967 ( .A(KEYINPUT49), .B(G137), .Z(n1254) );
XOR2_X1 U968 ( .A(n1075), .B(n1255), .Z(n1251) );
XNOR2_X1 U969 ( .A(G110), .B(n1256), .ZN(n1255) );
NAND2_X1 U970 ( .A1(G221), .A2(n1236), .ZN(n1256) );
AND2_X1 U971 ( .A1(G234), .A2(n1034), .ZN(n1236) );
XOR2_X1 U972 ( .A(n1257), .B(G125), .Z(n1075) );
AND2_X1 U973 ( .A1(n1046), .A2(n1258), .ZN(n1197) );
NAND2_X1 U974 ( .A1(n1047), .A2(n1259), .ZN(n1258) );
NAND4_X1 U975 ( .A1(G902), .A2(n1070), .A3(n1201), .A4(n1094), .ZN(n1259) );
INV_X1 U976 ( .A(G898), .ZN(n1094) );
XOR2_X1 U977 ( .A(G953), .B(KEYINPUT33), .Z(n1070) );
NAND3_X1 U978 ( .A1(n1201), .A2(n1034), .A3(G952), .ZN(n1047) );
NAND2_X1 U979 ( .A1(G237), .A2(n1260), .ZN(n1201) );
NAND2_X1 U980 ( .A1(n1261), .A2(n1262), .ZN(n1046) );
OR2_X1 U981 ( .A1(n1007), .A2(KEYINPUT53), .ZN(n1262) );
INV_X1 U982 ( .A(n1022), .ZN(n1007) );
NOR2_X1 U983 ( .A1(n1011), .A2(n1263), .ZN(n1022) );
NAND3_X1 U984 ( .A1(n1011), .A2(n1010), .A3(KEYINPUT53), .ZN(n1261) );
INV_X1 U985 ( .A(n1263), .ZN(n1010) );
NOR2_X1 U986 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
INV_X1 U987 ( .A(G214), .ZN(n1264) );
XNOR2_X1 U988 ( .A(n1266), .B(n1267), .ZN(n1011) );
NOR2_X1 U989 ( .A1(n1265), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U990 ( .A(G210), .B(KEYINPUT62), .ZN(n1268) );
NOR2_X1 U991 ( .A1(G902), .A2(G237), .ZN(n1265) );
NAND2_X1 U992 ( .A1(n1269), .A2(n1161), .ZN(n1266) );
XOR2_X1 U993 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U994 ( .A(n1159), .B(n1272), .Z(n1271) );
NAND2_X1 U995 ( .A1(n1273), .A2(KEYINPUT48), .ZN(n1272) );
XNOR2_X1 U996 ( .A(n1126), .B(n1274), .ZN(n1273) );
NOR2_X1 U997 ( .A1(G125), .A2(KEYINPUT22), .ZN(n1274) );
NAND2_X1 U998 ( .A1(n1275), .A2(n1034), .ZN(n1159) );
XNOR2_X1 U999 ( .A(G224), .B(KEYINPUT31), .ZN(n1275) );
NOR2_X1 U1000 ( .A1(KEYINPUT55), .A2(n1160), .ZN(n1270) );
XNOR2_X1 U1001 ( .A(n1092), .B(n1089), .ZN(n1160) );
INV_X1 U1002 ( .A(n1093), .ZN(n1089) );
XOR2_X1 U1003 ( .A(G110), .B(n1276), .Z(n1093) );
XOR2_X1 U1004 ( .A(KEYINPUT45), .B(G122), .Z(n1276) );
XNOR2_X1 U1005 ( .A(n1277), .B(n1278), .ZN(n1092) );
XOR2_X1 U1006 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U1007 ( .A(n1281), .B(n1205), .ZN(n1280) );
NAND2_X1 U1008 ( .A1(n1282), .A2(n1253), .ZN(n1281) );
XNOR2_X1 U1009 ( .A(KEYINPUT17), .B(KEYINPUT1), .ZN(n1282) );
NAND2_X1 U1010 ( .A1(KEYINPUT61), .A2(n1198), .ZN(n1279) );
INV_X1 U1011 ( .A(G101), .ZN(n1198) );
XOR2_X1 U1012 ( .A(n1283), .B(n1284), .Z(n1277) );
NOR2_X1 U1013 ( .A1(n1021), .A2(n1017), .ZN(n1041) );
AND2_X1 U1014 ( .A1(G221), .A2(n1250), .ZN(n1017) );
NAND2_X1 U1015 ( .A1(n1260), .A2(n1161), .ZN(n1250) );
XOR2_X1 U1016 ( .A(G234), .B(KEYINPUT30), .Z(n1260) );
INV_X1 U1017 ( .A(n1206), .ZN(n1021) );
XNOR2_X1 U1018 ( .A(n1285), .B(G469), .ZN(n1206) );
NAND2_X1 U1019 ( .A1(n1286), .A2(n1161), .ZN(n1285) );
XOR2_X1 U1020 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1021 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1022 ( .A(n1291), .B(n1292), .ZN(n1290) );
NOR2_X1 U1023 ( .A1(G110), .A2(KEYINPUT41), .ZN(n1292) );
NOR2_X1 U1024 ( .A1(KEYINPUT27), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U1025 ( .A(KEYINPUT14), .B(n1139), .ZN(n1293) );
NAND2_X1 U1026 ( .A1(G227), .A2(n1034), .ZN(n1139) );
INV_X1 U1027 ( .A(G953), .ZN(n1034) );
XNOR2_X1 U1028 ( .A(KEYINPUT47), .B(KEYINPUT44), .ZN(n1289) );
XNOR2_X1 U1029 ( .A(n1149), .B(n1294), .ZN(n1287) );
XOR2_X1 U1030 ( .A(n1295), .B(n1257), .Z(n1294) );
XNOR2_X1 U1031 ( .A(G140), .B(n1150), .ZN(n1257) );
XNOR2_X1 U1032 ( .A(G128), .B(n1226), .ZN(n1150) );
INV_X1 U1033 ( .A(G146), .ZN(n1226) );
XOR2_X1 U1034 ( .A(n1296), .B(n1074), .Z(n1149) );
INV_X1 U1035 ( .A(G143), .ZN(n1074) );
NAND2_X1 U1036 ( .A1(n1297), .A2(KEYINPUT56), .ZN(n1296) );
XOR2_X1 U1037 ( .A(n1283), .B(KEYINPUT50), .Z(n1297) );
XNOR2_X1 U1038 ( .A(G104), .B(n1244), .ZN(n1283) );
XOR2_X1 U1039 ( .A(G107), .B(KEYINPUT4), .Z(n1244) );
INV_X1 U1040 ( .A(n1194), .ZN(n1027) );
XNOR2_X1 U1041 ( .A(n1298), .B(G472), .ZN(n1194) );
NAND2_X1 U1042 ( .A1(n1299), .A2(n1161), .ZN(n1298) );
INV_X1 U1043 ( .A(G902), .ZN(n1161) );
XNOR2_X1 U1044 ( .A(n1126), .B(n1127), .ZN(n1299) );
XOR2_X1 U1045 ( .A(n1300), .B(n1301), .Z(n1127) );
XNOR2_X1 U1046 ( .A(n1205), .B(n1302), .ZN(n1301) );
XNOR2_X1 U1047 ( .A(KEYINPUT59), .B(n1253), .ZN(n1302) );
INV_X1 U1048 ( .A(G119), .ZN(n1253) );
INV_X1 U1049 ( .A(G113), .ZN(n1205) );
XOR2_X1 U1050 ( .A(n1303), .B(n1284), .Z(n1300) );
XOR2_X1 U1051 ( .A(G116), .B(KEYINPUT25), .Z(n1284) );
XOR2_X1 U1052 ( .A(n1295), .B(n1304), .Z(n1303) );
AND2_X1 U1053 ( .A1(n1223), .A2(G210), .ZN(n1304) );
NOR2_X1 U1054 ( .A1(G953), .A2(G237), .ZN(n1223) );
XNOR2_X1 U1055 ( .A(n1077), .B(G101), .ZN(n1295) );
XOR2_X1 U1056 ( .A(G131), .B(n1305), .Z(n1077) );
XNOR2_X1 U1057 ( .A(G137), .B(n1245), .ZN(n1305) );
INV_X1 U1058 ( .A(G134), .ZN(n1245) );
XOR2_X1 U1059 ( .A(G128), .B(n1306), .Z(n1126) );
NOR2_X1 U1060 ( .A1(KEYINPUT12), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1061 ( .A(G146), .B(G143), .ZN(n1307) );
endmodule


