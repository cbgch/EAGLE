//Key = 0010001011011011100111011101010101010110001111100101010111110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320;

XNOR2_X1 U714 ( .A(G107), .B(n1000), .ZN(G9) );
NOR2_X1 U715 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR3_X1 U716 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NAND3_X1 U717 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1003) );
NAND2_X1 U718 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U719 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND3_X1 U720 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NAND2_X1 U721 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U722 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U723 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U724 ( .A1(n1022), .A2(n1023), .ZN(n1016) );
NAND2_X1 U725 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XOR2_X1 U726 ( .A(KEYINPUT9), .B(n1026), .Z(n1024) );
NOR2_X1 U727 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U728 ( .A(KEYINPUT1), .B(n1029), .Z(n1028) );
NAND3_X1 U729 ( .A1(n1018), .A2(n1030), .A3(n1022), .ZN(n1011) );
NAND2_X1 U730 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U731 ( .A1(n1013), .A2(n1033), .ZN(n1032) );
NAND2_X1 U732 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U733 ( .A1(n1036), .A2(n1037), .A3(KEYINPUT56), .ZN(n1035) );
INV_X1 U734 ( .A(n1038), .ZN(n1034) );
NAND2_X1 U735 ( .A1(n1015), .A2(n1039), .ZN(n1031) );
NAND3_X1 U736 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
XNOR2_X1 U737 ( .A(KEYINPUT3), .B(n1043), .ZN(n1042) );
NAND2_X1 U738 ( .A1(n1013), .A2(n1044), .ZN(n1040) );
INV_X1 U739 ( .A(KEYINPUT56), .ZN(n1044) );
INV_X1 U740 ( .A(n1045), .ZN(n1009) );
NOR3_X1 U741 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1001) );
INV_X1 U742 ( .A(n1006), .ZN(n1046) );
NAND2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1006) );
NOR4_X1 U744 ( .A1(n1037), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1048) );
XOR2_X1 U745 ( .A(n1052), .B(n1053), .Z(n1051) );
XOR2_X1 U746 ( .A(KEYINPUT4), .B(n1054), .Z(n1053) );
NOR2_X1 U747 ( .A1(KEYINPUT22), .A2(G469), .ZN(n1054) );
XOR2_X1 U748 ( .A(n1055), .B(n1056), .Z(n1050) );
XOR2_X1 U749 ( .A(KEYINPUT14), .B(G472), .Z(n1056) );
NOR4_X1 U750 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1047) );
XOR2_X1 U751 ( .A(KEYINPUT48), .B(n1061), .Z(n1060) );
NOR3_X1 U752 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NOR2_X1 U753 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
AND3_X1 U754 ( .A1(n1066), .A2(n1065), .A3(KEYINPUT15), .ZN(n1063) );
NOR2_X1 U755 ( .A1(n1067), .A2(KEYINPUT28), .ZN(n1065) );
NOR2_X1 U756 ( .A1(KEYINPUT15), .A2(n1068), .ZN(n1062) );
XNOR2_X1 U757 ( .A(n1069), .B(KEYINPUT11), .ZN(n1057) );
XOR2_X1 U758 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U759 ( .A1(n1072), .A2(n1007), .ZN(n1071) );
NOR2_X1 U760 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U761 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
NAND2_X1 U762 ( .A1(n1077), .A2(n1007), .ZN(n1076) );
XNOR2_X1 U763 ( .A(n1004), .B(n1078), .ZN(n1077) );
OR3_X1 U764 ( .A1(n1074), .A2(n1078), .A3(n1007), .ZN(n1075) );
XNOR2_X1 U765 ( .A(n1079), .B(n1080), .ZN(n1078) );
XNOR2_X1 U766 ( .A(n1081), .B(n1082), .ZN(n1080) );
XNOR2_X1 U767 ( .A(G125), .B(n1083), .ZN(n1079) );
XNOR2_X1 U768 ( .A(KEYINPUT30), .B(n1084), .ZN(n1083) );
XOR2_X1 U769 ( .A(n1085), .B(n1086), .Z(G69) );
XOR2_X1 U770 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U771 ( .A1(G953), .A2(n1089), .ZN(n1088) );
NAND2_X1 U772 ( .A1(G898), .A2(G224), .ZN(n1089) );
NAND2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U774 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(n1090) );
XOR2_X1 U776 ( .A(n1095), .B(KEYINPUT55), .Z(n1094) );
NAND3_X1 U777 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
OR2_X1 U778 ( .A1(n1099), .A2(KEYINPUT43), .ZN(n1098) );
NAND3_X1 U779 ( .A1(KEYINPUT43), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U780 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NAND2_X1 U781 ( .A1(n1103), .A2(KEYINPUT43), .ZN(n1102) );
XNOR2_X1 U782 ( .A(n1099), .B(KEYINPUT42), .ZN(n1103) );
INV_X1 U783 ( .A(n1100), .ZN(n1101) );
AND2_X1 U784 ( .A1(n1005), .A2(n1007), .ZN(n1085) );
NOR2_X1 U785 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U786 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1110), .ZN(G63) );
XOR2_X1 U789 ( .A(KEYINPUT31), .B(n1111), .Z(n1110) );
NOR3_X1 U790 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR4_X1 U791 ( .A1(n1115), .A2(n1109), .A3(n1066), .A4(n1116), .ZN(n1114) );
INV_X1 U792 ( .A(KEYINPUT29), .ZN(n1115) );
NOR2_X1 U793 ( .A1(KEYINPUT29), .A2(n1117), .ZN(n1113) );
NOR2_X1 U794 ( .A1(n1066), .A2(n1109), .ZN(n1117) );
NOR2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
AND3_X1 U796 ( .A1(n1120), .A2(n1116), .A3(G478), .ZN(n1118) );
XOR2_X1 U797 ( .A(n1119), .B(KEYINPUT46), .Z(n1116) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1121), .ZN(G60) );
XNOR2_X1 U799 ( .A(n1122), .B(n1123), .ZN(n1121) );
AND2_X1 U800 ( .A1(G475), .A2(n1120), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(G6) );
NAND2_X1 U802 ( .A1(KEYINPUT63), .A2(n1126), .ZN(n1124) );
NOR2_X1 U803 ( .A1(n1104), .A2(n1127), .ZN(G57) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1129) );
AND2_X1 U806 ( .A1(G472), .A2(n1120), .ZN(n1130) );
XOR2_X1 U807 ( .A(n1132), .B(KEYINPUT58), .Z(n1128) );
NAND2_X1 U808 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1132) );
NAND2_X1 U809 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
XOR2_X1 U811 ( .A(KEYINPUT51), .B(n1139), .Z(n1134) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1138), .ZN(n1139) );
AND2_X1 U813 ( .A1(n1137), .A2(n1136), .ZN(n1140) );
NAND2_X1 U814 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
XNOR2_X1 U815 ( .A(n1143), .B(KEYINPUT57), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1104), .A2(n1144), .ZN(G54) );
XOR2_X1 U817 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U818 ( .A(n1147), .B(n1081), .ZN(n1146) );
NAND3_X1 U819 ( .A1(n1120), .A2(G469), .A3(KEYINPUT6), .ZN(n1147) );
INV_X1 U820 ( .A(n1109), .ZN(n1120) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1145) );
XNOR2_X1 U822 ( .A(n1150), .B(KEYINPUT24), .ZN(n1149) );
NAND2_X1 U823 ( .A1(KEYINPUT59), .A2(n1151), .ZN(n1150) );
XOR2_X1 U824 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U825 ( .A1(KEYINPUT38), .A2(n1154), .ZN(n1152) );
NAND2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
INV_X1 U827 ( .A(n1157), .ZN(n1156) );
XOR2_X1 U828 ( .A(n1158), .B(KEYINPUT50), .Z(n1155) );
NAND2_X1 U829 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U830 ( .A1(n1104), .A2(n1161), .ZN(G51) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U832 ( .A1(n1164), .A2(n1109), .ZN(n1163) );
NAND2_X1 U833 ( .A1(G902), .A2(n1165), .ZN(n1109) );
OR2_X1 U834 ( .A1(n1005), .A2(n1004), .ZN(n1165) );
NAND4_X1 U835 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1004) );
NOR4_X1 U836 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
AND2_X1 U837 ( .A1(n1174), .A2(n1175), .ZN(n1168) );
NAND3_X1 U838 ( .A1(n1015), .A2(n1176), .A3(n1177), .ZN(n1167) );
NAND2_X1 U839 ( .A1(n1038), .A2(n1178), .ZN(n1166) );
XOR2_X1 U840 ( .A(KEYINPUT26), .B(n1179), .Z(n1178) );
NAND2_X1 U841 ( .A1(n1180), .A2(n1181), .ZN(n1005) );
NOR4_X1 U842 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1125), .ZN(n1181) );
AND3_X1 U843 ( .A1(n1013), .A2(n1185), .A3(n1186), .ZN(n1125) );
INV_X1 U844 ( .A(n1187), .ZN(n1184) );
AND4_X1 U845 ( .A1(n1000), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1180) );
NAND3_X1 U846 ( .A1(n1186), .A2(n1191), .A3(n1192), .ZN(n1190) );
NAND3_X1 U847 ( .A1(n1176), .A2(n1185), .A3(n1013), .ZN(n1000) );
NOR2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1162) );
XOR2_X1 U849 ( .A(KEYINPUT13), .B(n1195), .Z(n1194) );
NOR2_X1 U850 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
AND2_X1 U851 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
XNOR2_X1 U852 ( .A(n1198), .B(n1199), .ZN(n1197) );
NAND2_X1 U853 ( .A1(KEYINPUT25), .A2(n1200), .ZN(n1198) );
XOR2_X1 U854 ( .A(KEYINPUT10), .B(n1201), .Z(n1200) );
NOR2_X1 U855 ( .A1(n1007), .A2(G952), .ZN(n1104) );
XNOR2_X1 U856 ( .A(G146), .B(n1202), .ZN(G48) );
NAND2_X1 U857 ( .A1(n1179), .A2(n1038), .ZN(n1202) );
AND2_X1 U858 ( .A1(n1203), .A2(n1186), .ZN(n1179) );
XNOR2_X1 U859 ( .A(G143), .B(n1175), .ZN(G45) );
NAND4_X1 U860 ( .A1(n1177), .A2(n1038), .A3(n1204), .A4(n1059), .ZN(n1175) );
NAND2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(G42) );
NAND2_X1 U862 ( .A1(n1207), .A2(n1084), .ZN(n1206) );
NAND2_X1 U863 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U864 ( .A1(n1174), .A2(n1210), .ZN(n1209) );
OR2_X1 U865 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
INV_X1 U866 ( .A(KEYINPUT61), .ZN(n1210) );
NAND2_X1 U867 ( .A1(G140), .A2(n1211), .ZN(n1205) );
NOR2_X1 U868 ( .A1(n1212), .A2(KEYINPUT60), .ZN(n1211) );
INV_X1 U869 ( .A(n1174), .ZN(n1212) );
NAND4_X1 U870 ( .A1(n1043), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1174) );
AND2_X1 U871 ( .A1(n1186), .A2(n1015), .ZN(n1215) );
XOR2_X1 U872 ( .A(G137), .B(n1173), .Z(G39) );
AND3_X1 U873 ( .A1(n1203), .A2(n1022), .A3(n1015), .ZN(n1173) );
XNOR2_X1 U874 ( .A(n1216), .B(n1217), .ZN(G36) );
NOR3_X1 U875 ( .A1(n1218), .A2(n1021), .A3(n1219), .ZN(n1217) );
XOR2_X1 U876 ( .A(KEYINPUT8), .B(n1015), .Z(n1218) );
XOR2_X1 U877 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U878 ( .A1(n1015), .A2(n1186), .A3(n1177), .ZN(n1172) );
INV_X1 U879 ( .A(n1219), .ZN(n1177) );
NAND3_X1 U880 ( .A1(n1214), .A2(n1213), .A3(n1191), .ZN(n1219) );
NOR2_X1 U881 ( .A1(n1069), .A2(n1037), .ZN(n1015) );
XOR2_X1 U882 ( .A(G128), .B(n1171), .Z(G30) );
AND3_X1 U883 ( .A1(n1176), .A2(n1038), .A3(n1203), .ZN(n1171) );
AND4_X1 U884 ( .A1(n1220), .A2(n1214), .A3(n1058), .A4(n1213), .ZN(n1203) );
XNOR2_X1 U885 ( .A(G101), .B(n1187), .ZN(G3) );
NAND3_X1 U886 ( .A1(n1022), .A2(n1185), .A3(n1191), .ZN(n1187) );
XNOR2_X1 U887 ( .A(G125), .B(n1221), .ZN(G27) );
NAND2_X1 U888 ( .A1(KEYINPUT16), .A2(n1170), .ZN(n1221) );
AND4_X1 U889 ( .A1(n1186), .A2(n1038), .A3(n1222), .A4(n1018), .ZN(n1170) );
AND2_X1 U890 ( .A1(n1213), .A2(n1043), .ZN(n1222) );
NAND2_X1 U891 ( .A1(n1045), .A2(n1223), .ZN(n1213) );
NAND4_X1 U892 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1074), .ZN(n1223) );
INV_X1 U893 ( .A(G900), .ZN(n1074) );
XOR2_X1 U894 ( .A(G122), .B(n1225), .Z(G24) );
NOR2_X1 U895 ( .A1(KEYINPUT62), .A2(n1189), .ZN(n1225) );
NAND4_X1 U896 ( .A1(n1192), .A2(n1013), .A3(n1204), .A4(n1059), .ZN(n1189) );
XNOR2_X1 U897 ( .A(G119), .B(n1188), .ZN(G21) );
NAND4_X1 U898 ( .A1(n1220), .A2(n1192), .A3(n1022), .A4(n1058), .ZN(n1188) );
XOR2_X1 U899 ( .A(G116), .B(n1183), .Z(G18) );
NOR3_X1 U900 ( .A1(n1041), .A2(n1021), .A3(n1226), .ZN(n1183) );
INV_X1 U901 ( .A(n1176), .ZN(n1021) );
NOR2_X1 U902 ( .A1(n1059), .A2(n1227), .ZN(n1176) );
INV_X1 U903 ( .A(n1191), .ZN(n1041) );
XNOR2_X1 U904 ( .A(G113), .B(n1228), .ZN(G15) );
NAND3_X1 U905 ( .A1(n1186), .A2(n1192), .A3(n1229), .ZN(n1228) );
XNOR2_X1 U906 ( .A(n1191), .B(KEYINPUT21), .ZN(n1229) );
NOR2_X1 U907 ( .A1(n1230), .A2(n1058), .ZN(n1191) );
INV_X1 U908 ( .A(n1226), .ZN(n1192) );
NAND2_X1 U909 ( .A1(n1231), .A2(n1018), .ZN(n1226) );
NAND2_X1 U910 ( .A1(n1232), .A2(n1233), .ZN(n1018) );
OR3_X1 U911 ( .A1(n1029), .A2(n1049), .A3(KEYINPUT1), .ZN(n1233) );
INV_X1 U912 ( .A(n1027), .ZN(n1049) );
NAND2_X1 U913 ( .A1(KEYINPUT1), .A2(n1214), .ZN(n1232) );
INV_X1 U914 ( .A(n1020), .ZN(n1186) );
NAND2_X1 U915 ( .A1(n1227), .A2(n1059), .ZN(n1020) );
INV_X1 U916 ( .A(n1204), .ZN(n1227) );
XNOR2_X1 U917 ( .A(G110), .B(n1234), .ZN(G12) );
NAND2_X1 U918 ( .A1(KEYINPUT49), .A2(n1182), .ZN(n1234) );
AND3_X1 U919 ( .A1(n1185), .A2(n1043), .A3(n1022), .ZN(n1182) );
NOR2_X1 U920 ( .A1(n1204), .A2(n1059), .ZN(n1022) );
XNOR2_X1 U921 ( .A(n1235), .B(G475), .ZN(n1059) );
NAND2_X1 U922 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XNOR2_X1 U923 ( .A(KEYINPUT7), .B(n1238), .ZN(n1236) );
INV_X1 U924 ( .A(n1122), .ZN(n1238) );
XNOR2_X1 U925 ( .A(n1239), .B(G113), .ZN(n1122) );
XOR2_X1 U926 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U927 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U928 ( .A(G122), .B(n1126), .ZN(n1243) );
XNOR2_X1 U929 ( .A(G143), .B(n1084), .ZN(n1242) );
XOR2_X1 U930 ( .A(n1244), .B(n1245), .Z(n1240) );
XOR2_X1 U931 ( .A(n1246), .B(n1247), .Z(n1245) );
NAND2_X1 U932 ( .A1(KEYINPUT44), .A2(n1248), .ZN(n1247) );
NAND2_X1 U933 ( .A1(KEYINPUT12), .A2(n1249), .ZN(n1246) );
XOR2_X1 U934 ( .A(n1250), .B(n1251), .Z(n1244) );
NAND2_X1 U935 ( .A1(G214), .A2(n1252), .ZN(n1250) );
XOR2_X1 U936 ( .A(n1253), .B(n1066), .Z(n1204) );
INV_X1 U937 ( .A(G478), .ZN(n1066) );
NAND2_X1 U938 ( .A1(KEYINPUT27), .A2(n1067), .ZN(n1253) );
INV_X1 U939 ( .A(n1068), .ZN(n1067) );
NAND2_X1 U940 ( .A1(n1119), .A2(n1237), .ZN(n1068) );
XNOR2_X1 U941 ( .A(n1254), .B(n1255), .ZN(n1119) );
XNOR2_X1 U942 ( .A(n1216), .B(n1256), .ZN(n1255) );
NOR2_X1 U943 ( .A1(KEYINPUT17), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U944 ( .A(G128), .B(n1258), .ZN(n1257) );
XOR2_X1 U945 ( .A(KEYINPUT54), .B(G143), .Z(n1258) );
INV_X1 U946 ( .A(G134), .ZN(n1216) );
XOR2_X1 U947 ( .A(n1259), .B(n1260), .Z(n1254) );
NOR2_X1 U948 ( .A1(KEYINPUT18), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U949 ( .A(G107), .B(n1262), .ZN(n1261) );
XOR2_X1 U950 ( .A(G122), .B(G116), .Z(n1262) );
NAND3_X1 U951 ( .A1(G234), .A2(n1007), .A3(G217), .ZN(n1259) );
NAND2_X1 U952 ( .A1(n1263), .A2(n1264), .ZN(n1043) );
NAND3_X1 U953 ( .A1(n1230), .A2(n1058), .A3(n1265), .ZN(n1264) );
INV_X1 U954 ( .A(KEYINPUT40), .ZN(n1265) );
NAND2_X1 U955 ( .A1(KEYINPUT40), .A2(n1013), .ZN(n1263) );
NOR2_X1 U956 ( .A1(n1058), .A2(n1220), .ZN(n1013) );
INV_X1 U957 ( .A(n1230), .ZN(n1220) );
XNOR2_X1 U958 ( .A(n1055), .B(n1266), .ZN(n1230) );
NOR2_X1 U959 ( .A1(G472), .A2(KEYINPUT32), .ZN(n1266) );
NAND2_X1 U960 ( .A1(n1267), .A2(n1237), .ZN(n1055) );
XOR2_X1 U961 ( .A(n1138), .B(n1268), .Z(n1267) );
XNOR2_X1 U962 ( .A(n1269), .B(n1131), .ZN(n1268) );
XOR2_X1 U963 ( .A(n1270), .B(n1271), .Z(n1131) );
INV_X1 U964 ( .A(G101), .ZN(n1271) );
NAND2_X1 U965 ( .A1(G210), .A2(n1252), .ZN(n1270) );
NOR2_X1 U966 ( .A1(G953), .A2(G237), .ZN(n1252) );
NAND3_X1 U967 ( .A1(n1272), .A2(n1273), .A3(n1137), .ZN(n1269) );
NAND2_X1 U968 ( .A1(n1081), .A2(n1274), .ZN(n1137) );
NAND2_X1 U969 ( .A1(KEYINPUT36), .A2(n1081), .ZN(n1273) );
OR3_X1 U970 ( .A1(n1274), .A2(KEYINPUT36), .A3(n1081), .ZN(n1272) );
XOR2_X1 U971 ( .A(n1275), .B(n1276), .Z(n1138) );
NOR2_X1 U972 ( .A1(G113), .A2(KEYINPUT34), .ZN(n1276) );
XNOR2_X1 U973 ( .A(G119), .B(n1277), .ZN(n1275) );
NOR2_X1 U974 ( .A1(G116), .A2(KEYINPUT5), .ZN(n1277) );
XOR2_X1 U975 ( .A(n1278), .B(n1108), .Z(n1058) );
NAND2_X1 U976 ( .A1(G217), .A2(n1279), .ZN(n1108) );
OR2_X1 U977 ( .A1(n1107), .A2(G902), .ZN(n1278) );
XNOR2_X1 U978 ( .A(n1280), .B(n1281), .ZN(n1107) );
XOR2_X1 U979 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U980 ( .A(n1284), .B(n1285), .ZN(n1283) );
AND3_X1 U981 ( .A1(G221), .A2(n1007), .A3(G234), .ZN(n1285) );
INV_X1 U982 ( .A(G110), .ZN(n1284) );
XNOR2_X1 U983 ( .A(n1248), .B(G119), .ZN(n1282) );
INV_X1 U984 ( .A(G125), .ZN(n1248) );
XOR2_X1 U985 ( .A(n1286), .B(n1287), .Z(n1280) );
XNOR2_X1 U986 ( .A(n1288), .B(n1289), .ZN(n1286) );
NAND2_X1 U987 ( .A1(KEYINPUT19), .A2(G137), .ZN(n1289) );
NAND2_X1 U988 ( .A1(KEYINPUT2), .A2(n1084), .ZN(n1288) );
INV_X1 U989 ( .A(G140), .ZN(n1084) );
AND2_X1 U990 ( .A1(n1231), .A2(n1214), .ZN(n1185) );
INV_X1 U991 ( .A(n1025), .ZN(n1214) );
NAND2_X1 U992 ( .A1(n1029), .A2(n1027), .ZN(n1025) );
NAND2_X1 U993 ( .A1(G221), .A2(n1279), .ZN(n1027) );
NAND2_X1 U994 ( .A1(G234), .A2(n1237), .ZN(n1279) );
XNOR2_X1 U995 ( .A(n1052), .B(G469), .ZN(n1029) );
NAND2_X1 U996 ( .A1(n1290), .A2(n1237), .ZN(n1052) );
XOR2_X1 U997 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U998 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U999 ( .A1(KEYINPUT39), .A2(n1153), .ZN(n1294) );
XNOR2_X1 U1000 ( .A(G110), .B(G140), .ZN(n1153) );
NAND3_X1 U1001 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1293) );
NAND2_X1 U1002 ( .A1(n1157), .A2(n1081), .ZN(n1297) );
NOR2_X1 U1003 ( .A1(n1160), .A2(n1159), .ZN(n1157) );
NAND2_X1 U1004 ( .A1(n1298), .A2(n1159), .ZN(n1296) );
XNOR2_X1 U1005 ( .A(n1160), .B(n1081), .ZN(n1298) );
INV_X1 U1006 ( .A(n1143), .ZN(n1081) );
NAND3_X1 U1007 ( .A1(n1143), .A2(n1160), .A3(n1299), .ZN(n1295) );
INV_X1 U1008 ( .A(n1159), .ZN(n1299) );
XOR2_X1 U1009 ( .A(G101), .B(n1300), .Z(n1159) );
NOR2_X1 U1010 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
AND3_X1 U1011 ( .A1(KEYINPUT52), .A2(n1303), .A3(G104), .ZN(n1302) );
INV_X1 U1012 ( .A(G107), .ZN(n1303) );
NOR2_X1 U1013 ( .A1(KEYINPUT52), .A2(n1304), .ZN(n1301) );
XNOR2_X1 U1014 ( .A(n1082), .B(KEYINPUT33), .ZN(n1160) );
XOR2_X1 U1015 ( .A(G143), .B(n1287), .Z(n1082) );
XNOR2_X1 U1016 ( .A(G128), .B(n1249), .ZN(n1287) );
INV_X1 U1017 ( .A(G146), .ZN(n1249) );
XNOR2_X1 U1018 ( .A(n1305), .B(n1251), .ZN(n1143) );
XOR2_X1 U1019 ( .A(G131), .B(KEYINPUT41), .Z(n1251) );
XNOR2_X1 U1020 ( .A(G134), .B(G137), .ZN(n1305) );
XNOR2_X1 U1021 ( .A(n1154), .B(KEYINPUT0), .ZN(n1291) );
NOR2_X1 U1022 ( .A1(n1073), .A2(G953), .ZN(n1154) );
INV_X1 U1023 ( .A(G227), .ZN(n1073) );
AND2_X1 U1024 ( .A1(n1038), .A2(n1306), .ZN(n1231) );
NAND2_X1 U1025 ( .A1(n1045), .A2(n1307), .ZN(n1306) );
NAND4_X1 U1026 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1092), .ZN(n1307) );
INV_X1 U1027 ( .A(G898), .ZN(n1092) );
NAND3_X1 U1028 ( .A1(n1224), .A2(n1007), .A3(G952), .ZN(n1045) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1224) );
NOR2_X1 U1030 ( .A1(n1036), .A2(n1037), .ZN(n1038) );
AND2_X1 U1031 ( .A1(n1308), .A2(G214), .ZN(n1037) );
XOR2_X1 U1032 ( .A(n1309), .B(KEYINPUT47), .Z(n1308) );
INV_X1 U1033 ( .A(n1069), .ZN(n1036) );
XOR2_X1 U1034 ( .A(n1310), .B(n1164), .Z(n1069) );
NAND2_X1 U1035 ( .A1(G210), .A2(n1309), .ZN(n1164) );
OR2_X1 U1036 ( .A1(G902), .A2(G237), .ZN(n1309) );
NAND2_X1 U1037 ( .A1(n1311), .A2(n1237), .ZN(n1310) );
INV_X1 U1038 ( .A(G902), .ZN(n1237) );
XOR2_X1 U1039 ( .A(n1312), .B(n1313), .Z(n1311) );
XNOR2_X1 U1040 ( .A(n1314), .B(n1196), .ZN(n1313) );
XNOR2_X1 U1041 ( .A(n1093), .B(n1315), .ZN(n1196) );
XNOR2_X1 U1042 ( .A(n1316), .B(n1099), .ZN(n1315) );
XNOR2_X1 U1043 ( .A(n1317), .B(n1304), .ZN(n1099) );
XNOR2_X1 U1044 ( .A(n1126), .B(G107), .ZN(n1304) );
INV_X1 U1045 ( .A(G104), .ZN(n1126) );
NAND2_X1 U1046 ( .A1(KEYINPUT20), .A2(G101), .ZN(n1317) );
NAND2_X1 U1047 ( .A1(KEYINPUT37), .A2(n1100), .ZN(n1316) );
XOR2_X1 U1048 ( .A(G113), .B(n1318), .Z(n1100) );
XOR2_X1 U1049 ( .A(G119), .B(G116), .Z(n1318) );
XNOR2_X1 U1050 ( .A(G110), .B(G122), .ZN(n1093) );
NAND2_X1 U1051 ( .A1(KEYINPUT53), .A2(n1199), .ZN(n1314) );
XNOR2_X1 U1052 ( .A(n1274), .B(G125), .ZN(n1199) );
INV_X1 U1053 ( .A(n1142), .ZN(n1274) );
XNOR2_X1 U1054 ( .A(n1319), .B(G128), .ZN(n1142) );
NAND2_X1 U1055 ( .A1(n1320), .A2(KEYINPUT23), .ZN(n1319) );
XNOR2_X1 U1056 ( .A(G143), .B(G146), .ZN(n1320) );
XOR2_X1 U1057 ( .A(KEYINPUT35), .B(n1201), .Z(n1312) );
AND2_X1 U1058 ( .A1(G224), .A2(n1007), .ZN(n1201) );
INV_X1 U1059 ( .A(G953), .ZN(n1007) );
endmodule


